// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_outs_enb,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_spare_0,
    i_spare_1,
    i_test_uc2,
    i_test_wci,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_outs_enb;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_spare_0;
 input i_spare_1;
 input i_test_uc2;
 input i_test_wci;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire net90;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net91;
 wire net106;
 wire net107;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net124;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net108;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire _00000_;
 wire _00001_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire clknet_0__03773_;
 wire clknet_0__03774_;
 wire clknet_0__03775_;
 wire clknet_0__03776_;
 wire clknet_0__03777_;
 wire clknet_0__03778_;
 wire clknet_0__03779_;
 wire clknet_0__03780_;
 wire clknet_0__03781_;
 wire clknet_0__03980_;
 wire clknet_0__03981_;
 wire clknet_0__03982_;
 wire clknet_0__03983_;
 wire clknet_0__03984_;
 wire clknet_0__03985_;
 wire clknet_0__03986_;
 wire clknet_0__03987_;
 wire clknet_0__03988_;
 wire clknet_0__03989_;
 wire clknet_0__03990_;
 wire clknet_0__03991_;
 wire clknet_0__03992_;
 wire clknet_0__03993_;
 wire clknet_0__03994_;
 wire clknet_0__03995_;
 wire clknet_0__03996_;
 wire clknet_0__03997_;
 wire clknet_0__03998_;
 wire clknet_0__03999_;
 wire clknet_0__04000_;
 wire clknet_0__04001_;
 wire clknet_0__04002_;
 wire clknet_0__04003_;
 wire clknet_0__04004_;
 wire clknet_0__04005_;
 wire clknet_0__04006_;
 wire clknet_0__04007_;
 wire clknet_0__04008_;
 wire clknet_0__04009_;
 wire clknet_0__04010_;
 wire clknet_0__04011_;
 wire clknet_0__04012_;
 wire clknet_0__04800_;
 wire clknet_0__05840_;
 wire clknet_0__05891_;
 wire clknet_0__05942_;
 wire clknet_0__05994_;
 wire clknet_0__06044_;
 wire clknet_0__06092_;
 wire clknet_0_i_clk;
 wire clknet_1_0__leaf__03773_;
 wire clknet_1_0__leaf__03774_;
 wire clknet_1_0__leaf__03775_;
 wire clknet_1_0__leaf__03776_;
 wire clknet_1_0__leaf__03777_;
 wire clknet_1_0__leaf__03778_;
 wire clknet_1_0__leaf__03779_;
 wire clknet_1_0__leaf__03780_;
 wire clknet_1_0__leaf__03781_;
 wire clknet_1_0__leaf__03980_;
 wire clknet_1_0__leaf__03981_;
 wire clknet_1_0__leaf__03982_;
 wire clknet_1_0__leaf__03983_;
 wire clknet_1_0__leaf__03984_;
 wire clknet_1_0__leaf__03985_;
 wire clknet_1_0__leaf__03986_;
 wire clknet_1_0__leaf__03987_;
 wire clknet_1_0__leaf__03988_;
 wire clknet_1_0__leaf__03989_;
 wire clknet_1_0__leaf__03990_;
 wire clknet_1_0__leaf__03991_;
 wire clknet_1_0__leaf__03992_;
 wire clknet_1_0__leaf__03993_;
 wire clknet_1_0__leaf__03994_;
 wire clknet_1_0__leaf__03995_;
 wire clknet_1_0__leaf__03996_;
 wire clknet_1_0__leaf__03997_;
 wire clknet_1_0__leaf__03998_;
 wire clknet_1_0__leaf__03999_;
 wire clknet_1_0__leaf__04000_;
 wire clknet_1_0__leaf__04001_;
 wire clknet_1_0__leaf__04002_;
 wire clknet_1_0__leaf__04003_;
 wire clknet_1_0__leaf__04004_;
 wire clknet_1_0__leaf__04005_;
 wire clknet_1_0__leaf__04006_;
 wire clknet_1_0__leaf__04007_;
 wire clknet_1_0__leaf__04008_;
 wire clknet_1_0__leaf__04009_;
 wire clknet_1_0__leaf__04010_;
 wire clknet_1_0__leaf__04011_;
 wire clknet_1_0__leaf__04012_;
 wire clknet_1_0__leaf__04800_;
 wire clknet_1_0__leaf__05840_;
 wire clknet_1_0__leaf__05891_;
 wire clknet_1_0__leaf__05942_;
 wire clknet_1_0__leaf__05994_;
 wire clknet_1_0__leaf__06044_;
 wire clknet_1_0__leaf__06092_;
 wire clknet_1_1__leaf__03773_;
 wire clknet_1_1__leaf__03774_;
 wire clknet_1_1__leaf__03775_;
 wire clknet_1_1__leaf__03776_;
 wire clknet_1_1__leaf__03777_;
 wire clknet_1_1__leaf__03778_;
 wire clknet_1_1__leaf__03779_;
 wire clknet_1_1__leaf__03780_;
 wire clknet_1_1__leaf__03781_;
 wire clknet_1_1__leaf__03980_;
 wire clknet_1_1__leaf__03981_;
 wire clknet_1_1__leaf__03982_;
 wire clknet_1_1__leaf__03983_;
 wire clknet_1_1__leaf__03984_;
 wire clknet_1_1__leaf__03985_;
 wire clknet_1_1__leaf__03986_;
 wire clknet_1_1__leaf__03987_;
 wire clknet_1_1__leaf__03988_;
 wire clknet_1_1__leaf__03989_;
 wire clknet_1_1__leaf__03990_;
 wire clknet_1_1__leaf__03991_;
 wire clknet_1_1__leaf__03992_;
 wire clknet_1_1__leaf__03993_;
 wire clknet_1_1__leaf__03994_;
 wire clknet_1_1__leaf__03995_;
 wire clknet_1_1__leaf__03996_;
 wire clknet_1_1__leaf__03997_;
 wire clknet_1_1__leaf__03998_;
 wire clknet_1_1__leaf__03999_;
 wire clknet_1_1__leaf__04000_;
 wire clknet_1_1__leaf__04001_;
 wire clknet_1_1__leaf__04002_;
 wire clknet_1_1__leaf__04003_;
 wire clknet_1_1__leaf__04004_;
 wire clknet_1_1__leaf__04005_;
 wire clknet_1_1__leaf__04006_;
 wire clknet_1_1__leaf__04007_;
 wire clknet_1_1__leaf__04008_;
 wire clknet_1_1__leaf__04009_;
 wire clknet_1_1__leaf__04010_;
 wire clknet_1_1__leaf__04011_;
 wire clknet_1_1__leaf__04012_;
 wire clknet_1_1__leaf__04800_;
 wire clknet_1_1__leaf__05840_;
 wire clknet_1_1__leaf__05891_;
 wire clknet_1_1__leaf__05942_;
 wire clknet_1_1__leaf__05994_;
 wire clknet_1_1__leaf__06044_;
 wire clknet_1_1__leaf__06092_;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_leaf_0_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_9_i_clk;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net1;
 wire net10;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net303;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net356;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net358;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net363;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net368;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net371;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net372;
 wire net3720;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net373;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net374;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net375;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net376;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3769;
 wire net377;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net378;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net379;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net38;
 wire net380;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net381;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net382;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net383;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net384;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3848;
 wire net3849;
 wire net385;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net386;
 wire net3860;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net387;
 wire net3870;
 wire net3871;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net388;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net389;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net39;
 wire net390;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net391;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net392;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net393;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net394;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net395;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net396;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net397;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net398;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net399;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4;
 wire net40;
 wire net400;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net401;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net402;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net403;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net404;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net405;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net406;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net407;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net408;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net409;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net41;
 wire net410;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net411;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net412;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net413;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net414;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net415;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net416;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net417;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net418;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net419;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net42;
 wire net420;
 wire net4200;
 wire net4201;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net421;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net422;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net423;
 wire net4230;
 wire net4231;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net424;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net425;
 wire net4250;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net426;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net427;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net428;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net429;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4298;
 wire net4299;
 wire net43;
 wire net430;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net431;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net432;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net433;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net434;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net435;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net436;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net437;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net438;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net439;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net44;
 wire net440;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net441;
 wire net4410;
 wire net4411;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4419;
 wire net442;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net443;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net444;
 wire net4440;
 wire net4441;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net445;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net446;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net447;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net448;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net449;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net45;
 wire net450;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net451;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net452;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net453;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net454;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net455;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net456;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net457;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net458;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net459;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net46;
 wire net460;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net461;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net462;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net463;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net464;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net465;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net466;
 wire net4660;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net467;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net468;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net469;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net47;
 wire net470;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net471;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net472;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net473;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net474;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net475;
 wire net4750;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4758;
 wire net4759;
 wire net476;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net477;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net478;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net479;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net48;
 wire net480;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net481;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net482;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net483;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net484;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net485;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net486;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net487;
 wire net4870;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net488;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net489;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net49;
 wire net490;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net491;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net492;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net493;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net494;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net495;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net496;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net497;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net498;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net499;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5;
 wire net50;
 wire net500;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net501;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net502;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net503;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net504;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net505;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net506;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net507;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net508;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net509;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net51;
 wire net510;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net511;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net512;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net513;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net514;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net515;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net516;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net517;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net518;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net519;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net52;
 wire net520;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net521;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net522;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net523;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net524;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net525;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net526;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net527;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net528;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net529;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net53;
 wire net530;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net531;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net532;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net533;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net534;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net535;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net536;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net537;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net538;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net539;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net54;
 wire net540;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net541;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net542;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net543;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net544;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net545;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net546;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net547;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net548;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net549;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net55;
 wire net550;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net551;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net552;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net553;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net554;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net555;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net556;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net557;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net558;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net559;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net56;
 wire net560;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net561;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net562;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net563;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net564;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net565;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net566;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net567;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net568;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net569;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net57;
 wire net570;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net571;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net572;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net573;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net574;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net575;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net576;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net577;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net578;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net579;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net58;
 wire net580;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net581;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net582;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net583;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net584;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net585;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net586;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net587;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net588;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net589;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net59;
 wire net590;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net591;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net592;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net593;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net594;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net595;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net596;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net597;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net598;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net599;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6;
 wire net60;
 wire net600;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net601;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net602;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net603;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net604;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net605;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net606;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6068;
 wire net6069;
 wire net607;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6079;
 wire net608;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6085;
 wire net6086;
 wire net6088;
 wire net6089;
 wire net609;
 wire net6091;
 wire net6092;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net61;
 wire net610;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6108;
 wire net6109;
 wire net611;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6116;
 wire net6117;
 wire net6119;
 wire net612;
 wire net6120;
 wire net6122;
 wire net6123;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net613;
 wire net6130;
 wire net6131;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6138;
 wire net6139;
 wire net614;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net615;
 wire net6150;
 wire net6151;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net616;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net617;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net618;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net619;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net62;
 wire net620;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net621;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net622;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net623;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net624;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net625;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net626;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net627;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net628;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net629;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net63;
 wire net630;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net631;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net632;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net633;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net634;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net635;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net636;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net637;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net638;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net639;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net64;
 wire net640;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net641;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net642;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net643;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net644;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net645;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net646;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net647;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net648;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net649;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net65;
 wire net650;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net651;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net652;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net653;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net654;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net655;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net656;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net657;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net658;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net659;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net66;
 wire net660;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net661;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net662;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net663;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net664;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net665;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net666;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net667;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net668;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net669;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net67;
 wire net670;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net671;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net672;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net673;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net674;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net675;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net676;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net677;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net678;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net679;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net68;
 wire net680;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net681;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net682;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net683;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net684;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net685;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net686;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net687;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net688;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net689;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net69;
 wire net690;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net691;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net692;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net693;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net694;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net695;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net696;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net697;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net698;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net699;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7;
 wire net70;
 wire net700;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net701;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net702;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net703;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net704;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net705;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net706;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net707;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net708;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net709;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net71;
 wire net710;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net711;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net712;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net713;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net714;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net715;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net716;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net717;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net718;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net719;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net72;
 wire net720;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net721;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net722;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net723;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net724;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net725;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net726;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net727;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net728;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net729;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net73;
 wire net730;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net731;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net732;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net733;
 wire net7330;
 wire net7331;
 wire net7333;
 wire net7335;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net734;
 wire net7341;
 wire net7343;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7349;
 wire net735;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net736;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net737;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net738;
 wire net7380;
 wire net7381;
 wire net739;
 wire net74;
 wire net740;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net741;
 wire net742;
 wire net7427;
 wire net7428;
 wire net743;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net744;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net745;
 wire net7450;
 wire net7451;
 wire net7453;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net746;
 wire net7460;
 wire net7464;
 wire net7467;
 wire net7468;
 wire net747;
 wire net7471;
 wire net7472;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net748;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net749;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net75;
 wire net750;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7506;
 wire net7507;
 wire net751;
 wire net7510;
 wire net7511;
 wire net7513;
 wire net7514;
 wire net7516;
 wire net7517;
 wire net7519;
 wire net752;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net753;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net754;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net755;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7557;
 wire net7558;
 wire net756;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7566;
 wire net7568;
 wire net7569;
 wire net757;
 wire net7571;
 wire net7572;
 wire net7573;
 wire net7575;
 wire net7576;
 wire net7577;
 wire net758;
 wire net7580;
 wire net7581;
 wire net7582;
 wire net7583;
 wire net7585;
 wire net7586;
 wire net7589;
 wire net759;
 wire net7590;
 wire net7594;
 wire net7595;
 wire net7596;
 wire net7598;
 wire net7599;
 wire net76;
 wire net760;
 wire net7601;
 wire net7602;
 wire net7606;
 wire net7608;
 wire net7609;
 wire net761;
 wire net7611;
 wire net7612;
 wire net7613;
 wire net7614;
 wire net7615;
 wire net7616;
 wire net7617;
 wire net7619;
 wire net762;
 wire net7620;
 wire net7621;
 wire net7622;
 wire net7623;
 wire net7624;
 wire net7625;
 wire net7627;
 wire net7628;
 wire net7629;
 wire net763;
 wire net7631;
 wire net7632;
 wire net7633;
 wire net7634;
 wire net7635;
 wire net7636;
 wire net7637;
 wire net7638;
 wire net7639;
 wire net764;
 wire net7640;
 wire net7641;
 wire net7642;
 wire net7643;
 wire net7644;
 wire net7645;
 wire net7646;
 wire net7647;
 wire net7648;
 wire net7649;
 wire net765;
 wire net7650;
 wire net7651;
 wire net7652;
 wire net7653;
 wire net7654;
 wire net7655;
 wire net7656;
 wire net7657;
 wire net7658;
 wire net7659;
 wire net766;
 wire net7660;
 wire net7661;
 wire net7662;
 wire net7663;
 wire net7664;
 wire net7665;
 wire net7666;
 wire net7667;
 wire net7668;
 wire net7669;
 wire net767;
 wire net7670;
 wire net7671;
 wire net7672;
 wire net7673;
 wire net7674;
 wire net7675;
 wire net7676;
 wire net7677;
 wire net7678;
 wire net7679;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net7711;
 wire net7712;
 wire net7717;
 wire net7718;
 wire net772;
 wire net7721;
 wire net7722;
 wire net7723;
 wire net7724;
 wire net7725;
 wire net7726;
 wire net773;
 wire net7731;
 wire net7732;
 wire net7733;
 wire net7735;
 wire net7736;
 wire net7737;
 wire net7738;
 wire net7739;
 wire net774;
 wire net7740;
 wire net7741;
 wire net7742;
 wire net7743;
 wire net7744;
 wire net7747;
 wire net7748;
 wire net775;
 wire net7750;
 wire net7751;
 wire net7752;
 wire net7753;
 wire net7754;
 wire net7757;
 wire net7759;
 wire net776;
 wire net7761;
 wire net7762;
 wire net7764;
 wire net7766;
 wire net7767;
 wire net7769;
 wire net777;
 wire net7770;
 wire net7771;
 wire net7773;
 wire net7775;
 wire net7777;
 wire net7779;
 wire net778;
 wire net7780;
 wire net7781;
 wire net7782;
 wire net7787;
 wire net7788;
 wire net7789;
 wire net779;
 wire net7790;
 wire net7791;
 wire net7792;
 wire net7793;
 wire net7794;
 wire net7795;
 wire net7796;
 wire net7797;
 wire net7798;
 wire net7799;
 wire net78;
 wire net780;
 wire net7800;
 wire net7801;
 wire net7804;
 wire net7805;
 wire net7806;
 wire net7807;
 wire net7809;
 wire net781;
 wire net7810;
 wire net7811;
 wire net7812;
 wire net7813;
 wire net7814;
 wire net7815;
 wire net7816;
 wire net7817;
 wire net7818;
 wire net7819;
 wire net782;
 wire net7820;
 wire net7822;
 wire net7823;
 wire net7824;
 wire net7825;
 wire net7826;
 wire net7827;
 wire net7828;
 wire net783;
 wire net7833;
 wire net7834;
 wire net7836;
 wire net7838;
 wire net7839;
 wire net784;
 wire net7840;
 wire net7843;
 wire net7844;
 wire net7845;
 wire net7846;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net7880;
 wire net7881;
 wire net7886;
 wire net7887;
 wire net7888;
 wire net789;
 wire net7891;
 wire net7892;
 wire net7899;
 wire net79;
 wire net790;
 wire net7900;
 wire net7901;
 wire net7902;
 wire net7904;
 wire net7906;
 wire net7907;
 wire net7908;
 wire net791;
 wire net7912;
 wire net7914;
 wire net7915;
 wire net7916;
 wire net7918;
 wire net792;
 wire net7923;
 wire net7924;
 wire net793;
 wire net7939;
 wire net794;
 wire net7942;
 wire net7945;
 wire net795;
 wire net7951;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net7999;
 wire net8;
 wire net80;
 wire net800;
 wire net8009;
 wire net801;
 wire net8010;
 wire net8016;
 wire net8017;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net8126;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.buf_floor[0] ;
 wire \rbzero.spi_registers.buf_floor[1] ;
 wire \rbzero.spi_registers.buf_floor[2] ;
 wire \rbzero.spi_registers.buf_floor[3] ;
 wire \rbzero.spi_registers.buf_floor[4] ;
 wire \rbzero.spi_registers.buf_floor[5] ;
 wire \rbzero.spi_registers.buf_leak[0] ;
 wire \rbzero.spi_registers.buf_leak[1] ;
 wire \rbzero.spi_registers.buf_leak[2] ;
 wire \rbzero.spi_registers.buf_leak[3] ;
 wire \rbzero.spi_registers.buf_leak[4] ;
 wire \rbzero.spi_registers.buf_leak[5] ;
 wire \rbzero.spi_registers.buf_mapdx[0] ;
 wire \rbzero.spi_registers.buf_mapdx[1] ;
 wire \rbzero.spi_registers.buf_mapdx[2] ;
 wire \rbzero.spi_registers.buf_mapdx[3] ;
 wire \rbzero.spi_registers.buf_mapdx[4] ;
 wire \rbzero.spi_registers.buf_mapdx[5] ;
 wire \rbzero.spi_registers.buf_mapdxw[0] ;
 wire \rbzero.spi_registers.buf_mapdxw[1] ;
 wire \rbzero.spi_registers.buf_mapdy[0] ;
 wire \rbzero.spi_registers.buf_mapdy[1] ;
 wire \rbzero.spi_registers.buf_mapdy[2] ;
 wire \rbzero.spi_registers.buf_mapdy[3] ;
 wire \rbzero.spi_registers.buf_mapdy[4] ;
 wire \rbzero.spi_registers.buf_mapdy[5] ;
 wire \rbzero.spi_registers.buf_mapdyw[0] ;
 wire \rbzero.spi_registers.buf_mapdyw[1] ;
 wire \rbzero.spi_registers.buf_otherx[0] ;
 wire \rbzero.spi_registers.buf_otherx[1] ;
 wire \rbzero.spi_registers.buf_otherx[2] ;
 wire \rbzero.spi_registers.buf_otherx[3] ;
 wire \rbzero.spi_registers.buf_otherx[4] ;
 wire \rbzero.spi_registers.buf_othery[0] ;
 wire \rbzero.spi_registers.buf_othery[1] ;
 wire \rbzero.spi_registers.buf_othery[2] ;
 wire \rbzero.spi_registers.buf_othery[3] ;
 wire \rbzero.spi_registers.buf_othery[4] ;
 wire \rbzero.spi_registers.buf_sky[0] ;
 wire \rbzero.spi_registers.buf_sky[1] ;
 wire \rbzero.spi_registers.buf_sky[2] ;
 wire \rbzero.spi_registers.buf_sky[3] ;
 wire \rbzero.spi_registers.buf_sky[4] ;
 wire \rbzero.spi_registers.buf_sky[5] ;
 wire \rbzero.spi_registers.buf_texadd0[0] ;
 wire \rbzero.spi_registers.buf_texadd0[10] ;
 wire \rbzero.spi_registers.buf_texadd0[11] ;
 wire \rbzero.spi_registers.buf_texadd0[12] ;
 wire \rbzero.spi_registers.buf_texadd0[13] ;
 wire \rbzero.spi_registers.buf_texadd0[14] ;
 wire \rbzero.spi_registers.buf_texadd0[15] ;
 wire \rbzero.spi_registers.buf_texadd0[16] ;
 wire \rbzero.spi_registers.buf_texadd0[17] ;
 wire \rbzero.spi_registers.buf_texadd0[18] ;
 wire \rbzero.spi_registers.buf_texadd0[19] ;
 wire \rbzero.spi_registers.buf_texadd0[1] ;
 wire \rbzero.spi_registers.buf_texadd0[20] ;
 wire \rbzero.spi_registers.buf_texadd0[21] ;
 wire \rbzero.spi_registers.buf_texadd0[22] ;
 wire \rbzero.spi_registers.buf_texadd0[23] ;
 wire \rbzero.spi_registers.buf_texadd0[2] ;
 wire \rbzero.spi_registers.buf_texadd0[3] ;
 wire \rbzero.spi_registers.buf_texadd0[4] ;
 wire \rbzero.spi_registers.buf_texadd0[5] ;
 wire \rbzero.spi_registers.buf_texadd0[6] ;
 wire \rbzero.spi_registers.buf_texadd0[7] ;
 wire \rbzero.spi_registers.buf_texadd0[8] ;
 wire \rbzero.spi_registers.buf_texadd0[9] ;
 wire \rbzero.spi_registers.buf_texadd1[0] ;
 wire \rbzero.spi_registers.buf_texadd1[10] ;
 wire \rbzero.spi_registers.buf_texadd1[11] ;
 wire \rbzero.spi_registers.buf_texadd1[12] ;
 wire \rbzero.spi_registers.buf_texadd1[13] ;
 wire \rbzero.spi_registers.buf_texadd1[14] ;
 wire \rbzero.spi_registers.buf_texadd1[15] ;
 wire \rbzero.spi_registers.buf_texadd1[16] ;
 wire \rbzero.spi_registers.buf_texadd1[17] ;
 wire \rbzero.spi_registers.buf_texadd1[18] ;
 wire \rbzero.spi_registers.buf_texadd1[19] ;
 wire \rbzero.spi_registers.buf_texadd1[1] ;
 wire \rbzero.spi_registers.buf_texadd1[20] ;
 wire \rbzero.spi_registers.buf_texadd1[21] ;
 wire \rbzero.spi_registers.buf_texadd1[22] ;
 wire \rbzero.spi_registers.buf_texadd1[23] ;
 wire \rbzero.spi_registers.buf_texadd1[2] ;
 wire \rbzero.spi_registers.buf_texadd1[3] ;
 wire \rbzero.spi_registers.buf_texadd1[4] ;
 wire \rbzero.spi_registers.buf_texadd1[5] ;
 wire \rbzero.spi_registers.buf_texadd1[6] ;
 wire \rbzero.spi_registers.buf_texadd1[7] ;
 wire \rbzero.spi_registers.buf_texadd1[8] ;
 wire \rbzero.spi_registers.buf_texadd1[9] ;
 wire \rbzero.spi_registers.buf_texadd2[0] ;
 wire \rbzero.spi_registers.buf_texadd2[10] ;
 wire \rbzero.spi_registers.buf_texadd2[11] ;
 wire \rbzero.spi_registers.buf_texadd2[12] ;
 wire \rbzero.spi_registers.buf_texadd2[13] ;
 wire \rbzero.spi_registers.buf_texadd2[14] ;
 wire \rbzero.spi_registers.buf_texadd2[15] ;
 wire \rbzero.spi_registers.buf_texadd2[16] ;
 wire \rbzero.spi_registers.buf_texadd2[17] ;
 wire \rbzero.spi_registers.buf_texadd2[18] ;
 wire \rbzero.spi_registers.buf_texadd2[19] ;
 wire \rbzero.spi_registers.buf_texadd2[1] ;
 wire \rbzero.spi_registers.buf_texadd2[20] ;
 wire \rbzero.spi_registers.buf_texadd2[21] ;
 wire \rbzero.spi_registers.buf_texadd2[22] ;
 wire \rbzero.spi_registers.buf_texadd2[23] ;
 wire \rbzero.spi_registers.buf_texadd2[2] ;
 wire \rbzero.spi_registers.buf_texadd2[3] ;
 wire \rbzero.spi_registers.buf_texadd2[4] ;
 wire \rbzero.spi_registers.buf_texadd2[5] ;
 wire \rbzero.spi_registers.buf_texadd2[6] ;
 wire \rbzero.spi_registers.buf_texadd2[7] ;
 wire \rbzero.spi_registers.buf_texadd2[8] ;
 wire \rbzero.spi_registers.buf_texadd2[9] ;
 wire \rbzero.spi_registers.buf_texadd3[0] ;
 wire \rbzero.spi_registers.buf_texadd3[10] ;
 wire \rbzero.spi_registers.buf_texadd3[11] ;
 wire \rbzero.spi_registers.buf_texadd3[12] ;
 wire \rbzero.spi_registers.buf_texadd3[13] ;
 wire \rbzero.spi_registers.buf_texadd3[14] ;
 wire \rbzero.spi_registers.buf_texadd3[15] ;
 wire \rbzero.spi_registers.buf_texadd3[16] ;
 wire \rbzero.spi_registers.buf_texadd3[17] ;
 wire \rbzero.spi_registers.buf_texadd3[18] ;
 wire \rbzero.spi_registers.buf_texadd3[19] ;
 wire \rbzero.spi_registers.buf_texadd3[1] ;
 wire \rbzero.spi_registers.buf_texadd3[20] ;
 wire \rbzero.spi_registers.buf_texadd3[21] ;
 wire \rbzero.spi_registers.buf_texadd3[22] ;
 wire \rbzero.spi_registers.buf_texadd3[23] ;
 wire \rbzero.spi_registers.buf_texadd3[2] ;
 wire \rbzero.spi_registers.buf_texadd3[3] ;
 wire \rbzero.spi_registers.buf_texadd3[4] ;
 wire \rbzero.spi_registers.buf_texadd3[5] ;
 wire \rbzero.spi_registers.buf_texadd3[6] ;
 wire \rbzero.spi_registers.buf_texadd3[7] ;
 wire \rbzero.spi_registers.buf_texadd3[8] ;
 wire \rbzero.spi_registers.buf_texadd3[9] ;
 wire \rbzero.spi_registers.buf_vinf ;
 wire \rbzero.spi_registers.buf_vshift[0] ;
 wire \rbzero.spi_registers.buf_vshift[1] ;
 wire \rbzero.spi_registers.buf_vshift[2] ;
 wire \rbzero.spi_registers.buf_vshift[3] ;
 wire \rbzero.spi_registers.buf_vshift[4] ;
 wire \rbzero.spi_registers.buf_vshift[5] ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.trace_state[0] ;
 wire \rbzero.trace_state[1] ;
 wire \rbzero.trace_state[2] ;
 wire \rbzero.trace_state[3] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \reg_gpout[0] ;
 wire \reg_gpout[1] ;
 wire \reg_gpout[2] ;
 wire \reg_gpout[3] ;
 wire \reg_gpout[4] ;
 wire \reg_gpout[5] ;
 wire reg_hsync;
 wire \reg_rgb[14] ;
 wire \reg_rgb[15] ;
 wire \reg_rgb[22] ;
 wire \reg_rgb[23] ;
 wire \reg_rgb[6] ;
 wire \reg_rgb[7] ;
 wire reg_vsync;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_05616_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_05781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_05892_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_08025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_08025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_08279_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_08873_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_09286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_09286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_10205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_10205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_10205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_10329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_10329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_10329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_10329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net3772));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net4050));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net4532));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net4779));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net4779));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net6146));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net6146));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_05051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_08195_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_08479_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_09284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_10454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_10454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net3222));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net3222));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net4090));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_04978_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_06045_));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_980 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_994 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__buf_4 _10598_ (.A(net4049),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_8 _10599_ (.A(net4050),
    .X(_04160_));
 sky130_fd_sc_hd__buf_4 _10600_ (.A(net4004),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_4 _10601_ (.A(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(net3992),
    .X(_04163_));
 sky130_fd_sc_hd__buf_2 _10603_ (.A(net4052),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_4 _10604_ (.A(net4053),
    .X(_04165_));
 sky130_fd_sc_hd__and3b_2 _10605_ (.A_N(_04162_),
    .B(net3993),
    .C(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__xor2_4 _10606_ (.A(net47),
    .B(net48),
    .X(_04167_));
 sky130_fd_sc_hd__and3_2 _10607_ (.A(_04160_),
    .B(_04166_),
    .C(net89),
    .X(_04168_));
 sky130_fd_sc_hd__buf_4 _10608_ (.A(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_4 _10609_ (.A(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(net2686),
    .A1(net51),
    .S(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(net2687),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(net7026),
    .A1(net2686),
    .S(_04170_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10613_ (.A(net2648),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(net6902),
    .A1(net7026),
    .S(_04170_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _10615_ (.A(net2263),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(net6516),
    .A1(net6902),
    .S(_04170_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _10617_ (.A(net1836),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(net2427),
    .A1(net6516),
    .S(_04170_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _10619_ (.A(net6518),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(net5824),
    .A1(net2427),
    .S(_04170_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(net5826),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(net5828),
    .A1(net5824),
    .S(_04170_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(net5830),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(net2820),
    .A1(net5828),
    .S(_04170_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(net2575),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(net7272),
    .A1(net2820),
    .S(_04170_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(net2821),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(net7161),
    .A1(net7272),
    .S(_04170_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(net2751),
    .X(_01577_));
 sky130_fd_sc_hd__clkbuf_4 _10630_ (.A(_04169_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(net7153),
    .A1(net7161),
    .S(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(net2572),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(net2602),
    .A1(net7153),
    .S(_04181_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10634_ (.A(net7155),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(net6910),
    .A1(net7181),
    .S(_04181_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _10636_ (.A(net2603),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(net6371),
    .A1(net6910),
    .S(_04181_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _10638_ (.A(net2138),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(net2066),
    .A1(net6371),
    .S(_04181_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _10640_ (.A(net6373),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(net2469),
    .A1(net6818),
    .S(_04181_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _10642_ (.A(net6820),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(net2405),
    .A1(net6906),
    .S(_04181_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(net6908),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(net7006),
    .A1(net2405),
    .S(_04181_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(net7008),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(net6564),
    .A1(net7006),
    .S(_04181_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(net2380),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(net2224),
    .A1(net6564),
    .S(_04181_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(net6566),
    .X(_01567_));
 sky130_fd_sc_hd__clkbuf_4 _10651_ (.A(_04169_),
    .X(_04192_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(net6688),
    .A1(net6782),
    .S(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _10653_ (.A(net2225),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(net2298),
    .A1(net6688),
    .S(_04192_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(net6690),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(net6848),
    .A1(net7044),
    .S(_04192_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _10657_ (.A(net2299),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(net5821),
    .A1(net6848),
    .S(_04192_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10659_ (.A(net2083),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(net1762),
    .A1(net5821),
    .S(_04192_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _10661_ (.A(net5823),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(net5798),
    .A1(net1762),
    .S(_04192_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(net5800),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(net5811),
    .A1(net5798),
    .S(_04192_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(net5813),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(net2518),
    .A1(net5811),
    .S(_04192_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(net2153),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(net6626),
    .A1(net2518),
    .S(_04192_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(net2519),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(net2568),
    .A1(net6626),
    .S(_04192_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(net6628),
    .X(_01557_));
 sky130_fd_sc_hd__clkbuf_4 _10672_ (.A(_04169_),
    .X(_04203_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(net7056),
    .A1(net7141),
    .S(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _10674_ (.A(net2569),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(net6760),
    .A1(net7056),
    .S(_04203_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _10676_ (.A(net2344),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _10677_ (.A0(net2635),
    .A1(net6760),
    .S(_04203_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _10678_ (.A(net6762),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(net6419),
    .A1(net7175),
    .S(_04203_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10680_ (.A(net2636),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(net5981),
    .A1(net6419),
    .S(_04203_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _10682_ (.A(net1180),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(net5914),
    .A1(net5981),
    .S(_04203_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _10684_ (.A(net5983),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(net2556),
    .A1(net5914),
    .S(_04203_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10686_ (.A(net5916),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(net2855),
    .A1(net7241),
    .S(_04203_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10688_ (.A(net2779),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(net7209),
    .A1(net2855),
    .S(_04203_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10690_ (.A(net2856),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(net6942),
    .A1(net7209),
    .S(_04203_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _10692_ (.A(net2485),
    .X(_01547_));
 sky130_fd_sc_hd__clkbuf_4 _10693_ (.A(_04169_),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(net6642),
    .A1(net6942),
    .S(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(net2374),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(net2328),
    .A1(net6642),
    .S(_04214_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(net6644),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(net2007),
    .A1(net6786),
    .S(_04214_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(net6788),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(net6359),
    .A1(net6852),
    .S(_04214_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10701_ (.A(net2008),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(net2827),
    .A1(net6359),
    .S(_04214_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _10703_ (.A(net6361),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(net7197),
    .A1(net7280),
    .S(_04214_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _10705_ (.A(net2828),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(net2702),
    .A1(net7197),
    .S(_04214_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(net7199),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(net6520),
    .A1(net7266),
    .S(_04214_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(net2703),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(net2728),
    .A1(net6520),
    .S(_04214_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(net6522),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(net2085),
    .A1(net7169),
    .S(_04214_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(net7171),
    .X(_01537_));
 sky130_fd_sc_hd__clkbuf_4 _10714_ (.A(_04169_),
    .X(_04225_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(net6880),
    .A1(net2085),
    .S(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _10716_ (.A(net6882),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(net5927),
    .A1(net1683),
    .S(_04225_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _10718_ (.A(net5929),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(net2699),
    .A1(net5976),
    .S(_04225_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _10720_ (.A(net2260),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(net6445),
    .A1(net2699),
    .S(_04225_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10722_ (.A(net2700),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(net1900),
    .A1(net6445),
    .S(_04225_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _10724_ (.A(net6447),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(net2221),
    .A1(net6868),
    .S(_04225_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(net6870),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(net6898),
    .A1(net7073),
    .S(_04225_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(net2222),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(net2382),
    .A1(net6898),
    .S(_04225_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(net6900),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(net7089),
    .A1(net2382),
    .S(_04225_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(net7091),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(net5857),
    .A1(net1458),
    .S(_04225_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _10734_ (.A(net5859),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_4 _10735_ (.A(_04169_),
    .X(_04236_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(net5886),
    .A1(net5857),
    .S(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(net5888),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(net7249),
    .A1(net5886),
    .S(_04236_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(net2724),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(net7278),
    .A1(net7249),
    .S(_04236_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(net2754),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(net6453),
    .A1(net2753),
    .S(_04236_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _10743_ (.A(net6455),
    .X(_01523_));
 sky130_fd_sc_hd__clkinv_8 _10744_ (.A(_04167_),
    .Y(_04241_));
 sky130_fd_sc_hd__or3b_4 _10745_ (.A(_04241_),
    .B(_04160_),
    .C_N(_04166_),
    .X(_04242_));
 sky130_fd_sc_hd__buf_4 _10746_ (.A(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_4 _10747_ (.A(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(net51),
    .A1(net2367),
    .S(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(net2368),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(net2367),
    .A1(net5942),
    .S(_04244_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(net2338),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(net5804),
    .A1(net1932),
    .S(_04244_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(net5806),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(net7018),
    .A1(net7004),
    .S(_04244_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(net1954),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(net7004),
    .A1(net2101),
    .S(_04244_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(net2102),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(net2101),
    .A1(net7121),
    .S(_04244_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(net1473),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(net7121),
    .A1(net7060),
    .S(_04244_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(net2680),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(net7060),
    .A1(net2756),
    .S(_04244_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(net7062),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(net7282),
    .A1(net7243),
    .S(_04244_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(net2757),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(net7243),
    .A1(net6395),
    .S(_04244_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(net2419),
    .X(_01513_));
 sky130_fd_sc_hd__clkbuf_4 _10768_ (.A(_04243_),
    .X(_04255_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(net6395),
    .A1(net1723),
    .S(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _10770_ (.A(net6397),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(net6652),
    .A1(net1976),
    .S(_04255_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _10772_ (.A(net6654),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(net7079),
    .A1(net2848),
    .S(_04255_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(net7081),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(net7292),
    .A1(net7193),
    .S(_04255_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(net2849),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(net7193),
    .A1(net6489),
    .S(_04255_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(net2690),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(net6489),
    .A1(net2499),
    .S(_04255_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(net6491),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(net7233),
    .A1(net7203),
    .S(_04255_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(net2500),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(net7203),
    .A1(net7191),
    .S(_04255_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(net2170),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(net7191),
    .A1(net6714),
    .S(_04255_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(net2623),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(net6714),
    .A1(net6465),
    .S(_04255_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(net1733),
    .X(_01503_));
 sky130_fd_sc_hd__clkbuf_4 _10789_ (.A(_04243_),
    .X(_04266_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(net6465),
    .A1(net2304),
    .S(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10791_ (.A(net6467),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10792_ (.A0(net6772),
    .A1(net2421),
    .S(_04266_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _10793_ (.A(net6774),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(net6936),
    .A1(net6704),
    .S(_04266_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10795_ (.A(net2422),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(net6704),
    .A1(net2759),
    .S(_04266_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _10797_ (.A(net6706),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(net7207),
    .A1(net6578),
    .S(_04266_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10799_ (.A(net2760),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(net6578),
    .A1(net2307),
    .S(_04266_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(net6580),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(net7173),
    .A1(net6828),
    .S(_04266_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(net2308),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(net6828),
    .A1(net2644),
    .S(_04266_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(net6830),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(net7163),
    .A1(net2845),
    .S(_04266_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(net7165),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(net7290),
    .A1(net6407),
    .S(_04266_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(net2846),
    .X(_01493_));
 sky130_fd_sc_hd__clkbuf_4 _10810_ (.A(_04243_),
    .X(_04277_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(net6407),
    .A1(net2445),
    .S(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _10812_ (.A(net6409),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10813_ (.A0(net6944),
    .A1(net2641),
    .S(_04277_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_1 _10814_ (.A(net6946),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(net7149),
    .A1(net2668),
    .S(_04277_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _10816_ (.A(net7151),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(net7284),
    .A1(net6796),
    .S(_04277_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _10818_ (.A(net2669),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(net6796),
    .A1(net6744),
    .S(_04277_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _10820_ (.A(net2061),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(net6744),
    .A1(net6604),
    .S(_04277_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(net1760),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(net6604),
    .A1(net2902),
    .S(_04277_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(net6606),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(net7309),
    .A1(net7262),
    .S(_04277_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(net2903),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(net7262),
    .A1(net6712),
    .S(_04277_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(net2852),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(net6712),
    .A1(net6403),
    .S(_04277_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(net2055),
    .X(_01483_));
 sky130_fd_sc_hd__clkbuf_4 _10831_ (.A(_04243_),
    .X(_04288_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(net6403),
    .A1(net1777),
    .S(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _10833_ (.A(net6405),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10834_ (.A0(net6632),
    .A1(net2475),
    .S(_04288_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _10835_ (.A(net6634),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(net7036),
    .A1(net6674),
    .S(_04288_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _10837_ (.A(net2476),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(net6674),
    .A1(net2376),
    .S(_04288_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _10839_ (.A(net6676),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(net6866),
    .A1(net6500),
    .S(_04288_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10841_ (.A(net2377),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(net6500),
    .A1(net2559),
    .S(_04288_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _10843_ (.A(net6502),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(net7221),
    .A1(net7069),
    .S(_04288_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _10845_ (.A(net2560),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(net7069),
    .A1(net7058),
    .S(_04288_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(net2041),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(net7058),
    .A1(net6702),
    .S(_04288_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _10849_ (.A(net2011),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _10850_ (.A0(net6702),
    .A1(net6437),
    .S(_04288_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _10851_ (.A(net1974),
    .X(_01473_));
 sky130_fd_sc_hd__clkbuf_4 _10852_ (.A(_04243_),
    .X(_04299_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(net6437),
    .A1(net2063),
    .S(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(net6439),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(net6698),
    .A1(net2458),
    .S(_04299_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(net6700),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(net7085),
    .A1(net6992),
    .S(_04299_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(net2459),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(net6992),
    .A1(net6531),
    .S(_04299_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(net2144),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(net6531),
    .A1(net2107),
    .S(_04299_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(net6533),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(net6824),
    .A1(net2292),
    .S(_04299_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(net6826),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(net7115),
    .A1(net2695),
    .S(_04299_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _10866_ (.A(net7117),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(net7235),
    .A1(net2682),
    .S(_04299_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _10868_ (.A(net7237),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(net7247),
    .A1(net7066),
    .S(_04299_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _10870_ (.A(net2683),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(net7066),
    .A1(net2714),
    .S(_04299_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _10872_ (.A(net2386),
    .X(_01463_));
 sky130_fd_sc_hd__clkbuf_4 _10873_ (.A(_04243_),
    .X(_04310_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(net7300),
    .A1(net6922),
    .S(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(net2715),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(net6922),
    .A1(net5911),
    .S(_04310_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(net2164),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(net5911),
    .A1(net5775),
    .S(_04310_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(net5913),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(net5775),
    .A1(net1488),
    .S(_04310_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(net5777),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(net2747),
    .A1(net52),
    .S(_04236_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(net2748),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(net6916),
    .A1(net2747),
    .S(_04236_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _10885_ (.A(net2721),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(net2057),
    .A1(net6916),
    .S(_04236_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _10887_ (.A(net6918),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(net2781),
    .A1(net6988),
    .S(_04236_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _10889_ (.A(net6990),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10890_ (.A0(net7167),
    .A1(net7177),
    .S(_04236_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _10891_ (.A(net2782),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _10892_ (.A0(net6411),
    .A1(net7167),
    .S(_04236_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _10893_ (.A(net2626),
    .X(_01453_));
 sky130_fd_sc_hd__clkbuf_4 _10894_ (.A(_04169_),
    .X(_04321_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(net2861),
    .A1(net6411),
    .S(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(net6413),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(net2496),
    .A1(net7304),
    .S(_04321_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(net7306),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(net7157),
    .A1(net2496),
    .S(_04321_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(net7159),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(net6904),
    .A1(net7157),
    .S(_04321_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(net2453),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(net5989),
    .A1(net6904),
    .S(_04321_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(net2335),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(net5893),
    .A1(net5989),
    .S(_04321_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(net5991),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(net2632),
    .A1(net5893),
    .S(_04321_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(net5895),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(net2762),
    .A1(net7229),
    .S(_04321_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(net7231),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(net7075),
    .A1(net2762),
    .S(_04321_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(net7077),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(net2253),
    .A1(net7075),
    .S(_04321_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(net2254),
    .X(_01443_));
 sky130_fd_sc_hd__clkbuf_4 _10915_ (.A(_04168_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_4 _10916_ (.A(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__mux2_1 _10917_ (.A0(net5931),
    .A1(net2253),
    .S(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _10918_ (.A(net933),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(net5844),
    .A1(net5931),
    .S(_04333_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _10920_ (.A(net5933),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(net2708),
    .A1(net5844),
    .S(_04333_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _10922_ (.A(net5846),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10923_ (.A0(net7127),
    .A1(net2708),
    .S(_04333_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _10924_ (.A(net2709),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10925_ (.A0(net6930),
    .A1(net7127),
    .S(_04333_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _10926_ (.A(net2462),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(net6752),
    .A1(net6930),
    .S(_04333_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _10928_ (.A(net2210),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10929_ (.A0(net2830),
    .A1(net6752),
    .S(_04333_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _10930_ (.A(net6754),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(net7101),
    .A1(net7288),
    .S(_04333_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _10932_ (.A(net2831),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10933_ (.A0(net2674),
    .A1(net7101),
    .S(_04333_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _10934_ (.A(net7103),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(net6367),
    .A1(net7227),
    .S(_04333_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(net2675),
    .X(_01433_));
 sky130_fd_sc_hd__clkbuf_4 _10937_ (.A(_04332_),
    .X(_04344_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(net2737),
    .A1(net6367),
    .S(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _10939_ (.A(net6369),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(net7034),
    .A1(net7213),
    .S(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _10941_ (.A(net2738),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(net6551),
    .A1(net7034),
    .S(_04344_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _10943_ (.A(net2046),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(net2125),
    .A1(net6551),
    .S(_04344_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _10945_ (.A(net6553),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10946_ (.A0(net5897),
    .A1(net6890),
    .S(_04344_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _10947_ (.A(net2126),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(net5854),
    .A1(net5897),
    .S(_04344_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _10949_ (.A(net5899),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10950_ (.A0(net2234),
    .A1(net5854),
    .S(_04344_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _10951_ (.A(net5856),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10952_ (.A0(net6582),
    .A1(net2234),
    .S(_04344_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _10953_ (.A(net2235),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10954_ (.A0(net1697),
    .A1(net6582),
    .S(_04344_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _10955_ (.A(net6584),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(net6433),
    .A1(net6850),
    .S(_04344_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _10957_ (.A(net1698),
    .X(_01423_));
 sky130_fd_sc_hd__clkbuf_4 _10958_ (.A(_04332_),
    .X(_04355_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(net2490),
    .A1(net6433),
    .S(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _10960_ (.A(net6435),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(net6982),
    .A1(net7183),
    .S(_04355_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _10962_ (.A(net2491),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10963_ (.A0(net6836),
    .A1(net6982),
    .S(_04355_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _10964_ (.A(net1866),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(net6512),
    .A1(net6836),
    .S(_04355_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _10966_ (.A(net1822),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10967_ (.A0(net2765),
    .A1(net6512),
    .S(_04355_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _10968_ (.A(net6514),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10969_ (.A0(net6894),
    .A1(net7133),
    .S(_04355_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _10970_ (.A(net2766),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(net2638),
    .A1(net6894),
    .S(_04355_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _10972_ (.A(net6896),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(net6856),
    .A1(net7109),
    .S(_04355_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _10974_ (.A(net2639),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10975_ (.A0(net2357),
    .A1(net6856),
    .S(_04355_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _10976_ (.A(net6858),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(net6415),
    .A1(net7052),
    .S(_04355_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _10978_ (.A(net2358),
    .X(_01413_));
 sky130_fd_sc_hd__clkbuf_4 _10979_ (.A(_04332_),
    .X(_04366_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(net1771),
    .A1(net6415),
    .S(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _10981_ (.A(net6417),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(net2134),
    .A1(net6646),
    .S(_04366_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(net6648),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(net6636),
    .A1(net6876),
    .S(_04366_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(net2135),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(net2004),
    .A1(net6636),
    .S(_04366_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _10987_ (.A(net6638),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(net6768),
    .A1(net6986),
    .S(_04366_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _10989_ (.A(net2005),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(net6527),
    .A1(net6768),
    .S(_04366_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _10991_ (.A(net1742),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(net2876),
    .A1(net6527),
    .S(_04366_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _10993_ (.A(net6529),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(net7022),
    .A1(net7286),
    .S(_04366_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _10995_ (.A(net2877),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(net2478),
    .A1(net7022),
    .S(_04366_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _10997_ (.A(net7024),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(net6343),
    .A1(net7105),
    .S(_04366_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _10999_ (.A(net2479),
    .X(_01403_));
 sky130_fd_sc_hd__clkbuf_4 _11000_ (.A(_04332_),
    .X(_04377_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(net2514),
    .A1(net6343),
    .S(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _11002_ (.A(net6345),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(net2599),
    .A1(net6958),
    .S(_04377_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(net6960),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(net2325),
    .A1(net7129),
    .S(_04377_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(net7131),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(net6778),
    .A1(net7145),
    .S(_04377_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(net2326),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(net5879),
    .A1(net6778),
    .S(_04377_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(net1980),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(net5831),
    .A1(net5879),
    .S(_04377_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _11012_ (.A(net5881),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(net2442),
    .A1(net5831),
    .S(_04377_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _11014_ (.A(net5833),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(net6481),
    .A1(net2442),
    .S(_04377_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _11016_ (.A(net6483),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(net52),
    .A1(net2771),
    .S(_04310_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _11018_ (.A(net2772),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(net2771),
    .A1(net6485),
    .S(_04310_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _11020_ (.A(net1983),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(net6485),
    .A1(net2671),
    .S(_04310_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _11022_ (.A(net6487),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(net7260),
    .A1(net7012),
    .S(_04310_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _11024_ (.A(net2672),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(net7012),
    .A1(net6998),
    .S(_04310_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _11026_ (.A(net2132),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(net6998),
    .A1(net2439),
    .S(_04310_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _11028_ (.A(net7000),
    .X(_01389_));
 sky130_fd_sc_hd__clkbuf_4 _11029_ (.A(_04243_),
    .X(_04392_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(net7064),
    .A1(net6543),
    .S(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _11031_ (.A(net2440),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(net6543),
    .A1(net2659),
    .S(_04392_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _11033_ (.A(net6545),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(net7099),
    .A1(net6684),
    .S(_04392_),
    .X(_04395_));
 sky130_fd_sc_hd__clkbuf_1 _11035_ (.A(net2660),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(net6684),
    .A1(net2897),
    .S(_04392_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _11037_ (.A(net6686),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(net7296),
    .A1(net6802),
    .S(_04392_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _11039_ (.A(net2898),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(net6802),
    .A1(net6383),
    .S(_04392_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _11041_ (.A(net1898),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _11042_ (.A0(net6383),
    .A1(net1950),
    .S(_04392_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _11043_ (.A(net6385),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _11044_ (.A0(net6932),
    .A1(net6878),
    .S(_04392_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _11045_ (.A(net1951),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _11046_ (.A0(net6878),
    .A1(net6618),
    .S(_04392_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _11047_ (.A(net1996),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _11048_ (.A0(net6618),
    .A1(net2662),
    .S(_04392_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _11049_ (.A(net6620),
    .X(_01379_));
 sky130_fd_sc_hd__buf_4 _11050_ (.A(_04242_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_4 _11051_ (.A(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(net7245),
    .A1(net6574),
    .S(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _11053_ (.A(net2663),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(net6574),
    .A1(net2550),
    .S(_04404_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(net6576),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(net6994),
    .A1(net2538),
    .S(_04404_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(net6996),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(net7143),
    .A1(net7095),
    .S(_04404_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(net2539),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(net7095),
    .A1(net6940),
    .S(_04404_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(net2266),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(net6940),
    .A1(net6449),
    .S(_04404_),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(net2219),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(net6449),
    .A1(net1765),
    .S(_04404_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(net6451),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(net6678),
    .A1(net2424),
    .S(_04404_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(net6680),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(net7113),
    .A1(net6962),
    .S(_04404_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(net2425),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(net6962),
    .A1(net2870),
    .S(_04404_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _11071_ (.A(net6964),
    .X(_01369_));
 sky130_fd_sc_hd__clkbuf_4 _11072_ (.A(_04403_),
    .X(_04415_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(net7302),
    .A1(net6610),
    .S(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(net2871),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(net6610),
    .A1(net2237),
    .S(_04415_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(net6612),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(net7028),
    .A1(net5985),
    .S(_04415_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(net2238),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(net5985),
    .A1(net5834),
    .S(_04415_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(net5987),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(net5834),
    .A1(net2024),
    .S(_04415_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _11082_ (.A(net5836),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(net2024),
    .A1(net6316),
    .S(_04415_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _11084_ (.A(net2025),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(net6316),
    .A1(net2313),
    .S(_04415_),
    .X(_04422_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(net6318),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(net6924),
    .A1(net6914),
    .S(_04415_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _11088_ (.A(net2314),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(net6914),
    .A1(net6770),
    .S(_04415_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(net2403),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(net6770),
    .A1(net6457),
    .S(_04415_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _11092_ (.A(net2049),
    .X(_01359_));
 sky130_fd_sc_hd__clkbuf_4 _11093_ (.A(_04403_),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(net6457),
    .A1(net2527),
    .S(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(net6459),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(net7032),
    .A1(net6666),
    .S(_04426_),
    .X(_04428_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(net2528),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(net6666),
    .A1(net2128),
    .S(_04426_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(net6668),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(net7083),
    .A1(net6844),
    .S(_04426_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(net2129),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(net6844),
    .A1(net6664),
    .S(_04426_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _11103_ (.A(net2361),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(net6664),
    .A1(net6379),
    .S(_04426_),
    .X(_04432_));
 sky130_fd_sc_hd__clkbuf_1 _11105_ (.A(net1675),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(net6379),
    .A1(net2740),
    .S(_04426_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _11107_ (.A(net6381),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(net7274),
    .A1(net6716),
    .S(_04426_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _11109_ (.A(net2741),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(net6716),
    .A1(net2717),
    .S(_04426_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(net6718),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(net7255),
    .A1(net7217),
    .S(_04426_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _11113_ (.A(net2718),
    .X(_01349_));
 sky130_fd_sc_hd__clkbuf_4 _11114_ (.A(_04403_),
    .X(_04437_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(net7217),
    .A1(net6670),
    .S(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(net2666),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(net6670),
    .A1(net1935),
    .S(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(net6672),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(net6966),
    .A1(net2271),
    .S(_04437_),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(net6968),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(net7050),
    .A1(net6892),
    .S(_04437_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(net2272),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _11123_ (.A0(net6892),
    .A1(net6640),
    .S(_04437_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _11124_ (.A(net1986),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(net6640),
    .A1(net6391),
    .S(_04437_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _11126_ (.A(net1889),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(net6391),
    .A1(net1750),
    .S(_04437_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(net6393),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(net7016),
    .A1(net6980),
    .S(_04437_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(net1751),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _11131_ (.A0(net6980),
    .A1(net6656),
    .S(_04437_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _11132_ (.A(net2117),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(net6656),
    .A1(net2521),
    .S(_04437_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _11134_ (.A(net6658),
    .X(_01339_));
 sky130_fd_sc_hd__buf_4 _11135_ (.A(_04403_),
    .X(_04448_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(net7111),
    .A1(net6792),
    .S(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(net2522),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(net6792),
    .A1(net2616),
    .S(_04448_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _11139_ (.A(net6794),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _11140_ (.A0(net7093),
    .A1(net7071),
    .S(_04448_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_1 _11141_ (.A(net2617),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(net7071),
    .A1(net6756),
    .S(_04448_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(net1927),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(net6756),
    .A1(net6570),
    .S(_04448_),
    .X(_04453_));
 sky130_fd_sc_hd__clkbuf_1 _11145_ (.A(net2350),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(net6570),
    .A1(net750),
    .S(_04448_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _11147_ (.A(net6572),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(net750),
    .A1(net5920),
    .S(_04448_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(net5922),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(net5920),
    .A1(net5935),
    .S(_04448_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(net5937),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(net2449),
    .A1(net53),
    .S(_04377_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _11153_ (.A(net2450),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(net6547),
    .A1(net2449),
    .S(_04377_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(net2244),
    .X(_01329_));
 sky130_fd_sc_hd__clkbuf_4 _11156_ (.A(_04332_),
    .X(_04459_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(net5848),
    .A1(net6547),
    .S(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(net1519),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(net5814),
    .A1(net5848),
    .S(_04459_),
    .X(_04461_));
 sky130_fd_sc_hd__clkbuf_1 _11160_ (.A(net5850),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(net2140),
    .A1(net5814),
    .S(_04459_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _11162_ (.A(net5816),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(net2212),
    .A1(net6884),
    .S(_04459_),
    .X(_04463_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(net6886),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(net2578),
    .A1(net7119),
    .S(_04459_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_1 _11166_ (.A(net2566),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(net6441),
    .A1(net2578),
    .S(_04459_),
    .X(_04465_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(net2579),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(net1485),
    .A1(net6441),
    .S(_04459_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(net6443),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(net2149),
    .A1(net6594),
    .S(_04459_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(net6596),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(net2743),
    .A1(net6764),
    .S(_04459_),
    .X(_04468_));
 sky130_fd_sc_hd__clkbuf_1 _11174_ (.A(net6766),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(net6814),
    .A1(net7239),
    .S(_04459_),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(net2744),
    .X(_01319_));
 sky130_fd_sc_hd__clkbuf_4 _11177_ (.A(_04332_),
    .X(_04470_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(net2249),
    .A1(net6814),
    .S(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _11179_ (.A(net6816),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(net7042),
    .A1(net7046),
    .S(_04470_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_1 _11181_ (.A(net2250),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(net6972),
    .A1(net7042),
    .S(_04470_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _11183_ (.A(net2323),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(net2544),
    .A1(net6972),
    .S(_04470_),
    .X(_04474_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(net6974),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(net6842),
    .A1(net7215),
    .S(_04470_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _11187_ (.A(net2545),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(net6387),
    .A1(net6842),
    .S(_04470_),
    .X(_04476_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(net2201),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(net1372),
    .A1(net6387),
    .S(_04470_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _11191_ (.A(net6389),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(net2188),
    .A1(net6425),
    .S(_04470_),
    .X(_04478_));
 sky130_fd_sc_hd__clkbuf_1 _11193_ (.A(net6427),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(net5904),
    .A1(net6750),
    .S(_04470_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _11195_ (.A(net2189),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(net5868),
    .A1(net5904),
    .S(_04470_),
    .X(_04480_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(net5906),
    .X(_01309_));
 sky130_fd_sc_hd__clkbuf_4 _11198_ (.A(_04332_),
    .X(_04481_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(net1856),
    .A1(net5868),
    .S(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(net5870),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(net1923),
    .A1(net6736),
    .S(_04481_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _11202_ (.A(net6738),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(net2173),
    .A1(net7225),
    .S(_04481_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(net2174),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(net7097),
    .A1(net2173),
    .S(_04481_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(net1757),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(net7107),
    .A1(net7097),
    .S(_04481_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(net2597),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(net6421),
    .A1(net7107),
    .S(_04481_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(net2588),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(net2227),
    .A1(net6421),
    .S(_04481_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(net6423),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(net6790),
    .A1(net6912),
    .S(_04481_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(net2228),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(net6776),
    .A1(net6790),
    .S(_04481_),
    .X(_04490_));
 sky130_fd_sc_hd__clkbuf_1 _11216_ (.A(net2207),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(net6493),
    .A1(net6776),
    .S(_04481_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(net1810),
    .X(_01299_));
 sky130_fd_sc_hd__clkbuf_4 _11219_ (.A(_04332_),
    .X(_04492_));
 sky130_fd_sc_hd__mux2_1 _11220_ (.A0(net2508),
    .A1(net6493),
    .S(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _11221_ (.A(net6495),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _11222_ (.A0(net7054),
    .A1(net7201),
    .S(_04492_),
    .X(_04494_));
 sky130_fd_sc_hd__clkbuf_1 _11223_ (.A(net2509),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _11224_ (.A0(net5872),
    .A1(net7054),
    .S(_04492_),
    .X(_04495_));
 sky130_fd_sc_hd__clkbuf_1 _11225_ (.A(net2186),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(net5865),
    .A1(net5872),
    .S(_04492_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_1 _11227_ (.A(net5874),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(net2197),
    .A1(net5865),
    .S(_04492_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_1 _11229_ (.A(net5867),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(net6504),
    .A1(net2197),
    .S(_04492_),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _11231_ (.A(net2198),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(net5962),
    .A1(net6504),
    .S(_04492_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_1 _11233_ (.A(net1384),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(net5900),
    .A1(net5962),
    .S(_04492_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(net5964),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(net2412),
    .A1(net5900),
    .S(_04492_),
    .X(_04501_));
 sky130_fd_sc_hd__clkbuf_1 _11237_ (.A(net5902),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(net6539),
    .A1(net2412),
    .S(_04492_),
    .X(_04502_));
 sky130_fd_sc_hd__clkbuf_1 _11239_ (.A(net2413),
    .X(_01289_));
 sky130_fd_sc_hd__clkbuf_4 _11240_ (.A(_04332_),
    .X(_04503_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(net2796),
    .A1(net6539),
    .S(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _11242_ (.A(net6541),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(net6926),
    .A1(net7251),
    .S(_04503_),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_1 _11244_ (.A(net2797),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _11245_ (.A0(net6708),
    .A1(net6926),
    .S(_04503_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _11246_ (.A(net2167),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(net1880),
    .A1(net6708),
    .S(_04503_),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_1 _11248_ (.A(net6710),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(net6696),
    .A1(net6758),
    .S(_04503_),
    .X(_04508_));
 sky130_fd_sc_hd__clkbuf_1 _11250_ (.A(net1881),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(net6375),
    .A1(net6696),
    .S(_04503_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(net1801),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _11253_ (.A0(net2866),
    .A1(net6375),
    .S(_04503_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _11254_ (.A(net6377),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(net6938),
    .A1(net7253),
    .S(_04503_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_1 _11256_ (.A(net2867),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(net6862),
    .A1(net6938),
    .S(_04503_),
    .X(_04512_));
 sky130_fd_sc_hd__clkbuf_1 _11258_ (.A(net2585),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(net2881),
    .A1(net6862),
    .S(_04503_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _11260_ (.A(net6864),
    .X(_01279_));
 sky130_fd_sc_hd__clkbuf_4 _11261_ (.A(_04168_),
    .X(_04514_));
 sky130_fd_sc_hd__mux2_1 _11262_ (.A0(net7187),
    .A1(net7298),
    .S(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_1 _11263_ (.A(net2882),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _11264_ (.A0(net2858),
    .A1(net7187),
    .S(_04514_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _11265_ (.A(net7189),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _11266_ (.A0(net6860),
    .A1(net7268),
    .S(_04514_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_1 _11267_ (.A(net2859),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(net6810),
    .A1(net6860),
    .S(_04514_),
    .X(_04518_));
 sky130_fd_sc_hd__clkbuf_1 _11269_ (.A(net2320),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _11270_ (.A0(net2653),
    .A1(net6810),
    .S(_04514_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _11271_ (.A(net6812),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(net6337),
    .A1(net7002),
    .S(_04514_),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_1 _11273_ (.A(net2654),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _11274_ (.A0(net2436),
    .A1(net6337),
    .S(_04514_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_1 _11275_ (.A(net6339),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _11276_ (.A0(net6780),
    .A1(net7020),
    .S(_04514_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _11277_ (.A(net2437),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _11278_ (.A0(net5890),
    .A1(net6780),
    .S(_04514_),
    .X(_04523_));
 sky130_fd_sc_hd__clkbuf_1 _11279_ (.A(net2105),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(net5841),
    .A1(net5890),
    .S(_04514_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_1 _11281_ (.A(net5892),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(net2037),
    .A1(net5841),
    .S(_04169_),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_1 _11283_ (.A(net5843),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _11284_ (.A0(net6473),
    .A1(net2037),
    .S(_04169_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_1 _11285_ (.A(net6475),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _11286_ (.A0(net53),
    .A1(net2034),
    .S(_04448_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _11287_ (.A(net2035),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(net2034),
    .A1(net7087),
    .S(_04448_),
    .X(_04528_));
 sky130_fd_sc_hd__clkbuf_1 _11289_ (.A(net1930),
    .X(_01172_));
 sky130_fd_sc_hd__clkbuf_4 _11290_ (.A(_04403_),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _11291_ (.A0(net7087),
    .A1(net6692),
    .S(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__clkbuf_1 _11292_ (.A(net2416),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(net6692),
    .A1(net6506),
    .S(_04529_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_1 _11294_ (.A(net1907),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(net6506),
    .A1(net5953),
    .S(_04529_),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_1 _11296_ (.A(net1462),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(net5953),
    .A1(net5817),
    .S(_04529_),
    .X(_04533_));
 sky130_fd_sc_hd__clkbuf_1 _11298_ (.A(net5955),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(net5817),
    .A1(net2289),
    .S(_04529_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_1 _11300_ (.A(net5819),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(net2289),
    .A1(net7038),
    .S(_04529_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(net2290),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(net7038),
    .A1(net2613),
    .S(_04529_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _11304_ (.A(net7040),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(net7294),
    .A1(net6846),
    .S(_04529_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(net2614),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _11307_ (.A0(net6846),
    .A1(net6614),
    .S(_04529_),
    .X(_04538_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(net2147),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(net6614),
    .A1(net2799),
    .S(_04529_),
    .X(_04539_));
 sky130_fd_sc_hd__clkbuf_1 _11310_ (.A(net6616),
    .X(_01162_));
 sky130_fd_sc_hd__clkbuf_4 _11311_ (.A(_04403_),
    .X(_04540_));
 sky130_fd_sc_hd__mux2_1 _11312_ (.A0(net7270),
    .A1(net6742),
    .S(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_1 _11313_ (.A(net2800),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _11314_ (.A0(net6742),
    .A1(net6399),
    .S(_04540_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _11315_ (.A(net1816),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _11316_ (.A0(net6399),
    .A1(net2346),
    .S(_04540_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _11317_ (.A(net6401),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _11318_ (.A0(net7135),
    .A1(net7123),
    .S(_04540_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_1 _11319_ (.A(net2347),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _11320_ (.A0(net7123),
    .A1(net6976),
    .S(_04540_),
    .X(_04545_));
 sky130_fd_sc_hd__clkbuf_1 _11321_ (.A(net2503),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _11322_ (.A0(net6976),
    .A1(net6469),
    .S(_04540_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _11323_ (.A(net1962),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(net6469),
    .A1(net1753),
    .S(_04540_),
    .X(_04547_));
 sky130_fd_sc_hd__clkbuf_1 _11325_ (.A(net6471),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _11326_ (.A0(net6724),
    .A1(net2316),
    .S(_04540_),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_1 _11327_ (.A(net6726),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(net7179),
    .A1(net7014),
    .S(_04540_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_1 _11329_ (.A(net2317),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(net7014),
    .A1(net6728),
    .S(_04540_),
    .X(_04550_));
 sky130_fd_sc_hd__clkbuf_1 _11331_ (.A(net2531),
    .X(_01152_));
 sky130_fd_sc_hd__clkbuf_4 _11332_ (.A(_04403_),
    .X(_04551_));
 sky130_fd_sc_hd__mux2_1 _11333_ (.A0(net6728),
    .A1(net6592),
    .S(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _11334_ (.A(net2391),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _11335_ (.A0(net6592),
    .A1(net6429),
    .S(_04551_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_1 _11336_ (.A(net1825),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _11337_ (.A0(net6429),
    .A1(net2399),
    .S(_04551_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_1 _11338_ (.A(net6431),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _11339_ (.A0(net7030),
    .A1(net6888),
    .S(_04551_),
    .X(_04555_));
 sky130_fd_sc_hd__clkbuf_1 _11340_ (.A(net2400),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _11341_ (.A0(net6888),
    .A1(net6746),
    .S(_04551_),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _11342_ (.A(net2582),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _11343_ (.A0(net6746),
    .A1(net2051),
    .S(_04551_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_1 _11344_ (.A(net6748),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _11345_ (.A0(net6956),
    .A1(net6535),
    .S(_04551_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _11346_ (.A(net2052),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _11347_ (.A0(net6535),
    .A1(net2331),
    .S(_04551_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _11348_ (.A(net6537),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _11349_ (.A0(net6838),
    .A1(net2027),
    .S(_04551_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _11350_ (.A(net6840),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _11351_ (.A0(net6872),
    .A1(net2619),
    .S(_04551_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _11352_ (.A(net6874),
    .X(_01142_));
 sky130_fd_sc_hd__clkbuf_4 _11353_ (.A(_04403_),
    .X(_04562_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(net7223),
    .A1(net6822),
    .S(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _11355_ (.A(net2620),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _11356_ (.A0(net6822),
    .A1(net6477),
    .S(_04562_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _11357_ (.A(net1895),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _11358_ (.A0(net6477),
    .A1(net2295),
    .S(_04562_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _11359_ (.A(net6479),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _11360_ (.A0(net6832),
    .A1(net2430),
    .S(_04562_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_1 _11361_ (.A(net6834),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _11362_ (.A0(net6934),
    .A1(net6804),
    .S(_04562_),
    .X(_04567_));
 sky130_fd_sc_hd__clkbuf_1 _11363_ (.A(net2431),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _11364_ (.A0(net6804),
    .A1(net6508),
    .S(_04562_),
    .X(_04568_));
 sky130_fd_sc_hd__clkbuf_1 _11365_ (.A(net2278),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _11366_ (.A0(net6508),
    .A1(net2804),
    .S(_04562_),
    .X(_04569_));
 sky130_fd_sc_hd__clkbuf_1 _11367_ (.A(net6510),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(net7258),
    .A1(net6806),
    .S(_04562_),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_1 _11369_ (.A(net2805),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _11370_ (.A0(net6806),
    .A1(net2030),
    .S(_04562_),
    .X(_04571_));
 sky130_fd_sc_hd__clkbuf_1 _11371_ (.A(net6808),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _11372_ (.A0(net6948),
    .A1(net2711),
    .S(_04562_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_1 _11373_ (.A(net6950),
    .X(_01132_));
 sky130_fd_sc_hd__clkbuf_4 _11374_ (.A(_04403_),
    .X(_04573_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(net7125),
    .A1(net7048),
    .S(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__clkbuf_1 _11376_ (.A(net2712),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(net7048),
    .A1(net6351),
    .S(_04573_),
    .X(_04575_));
 sky130_fd_sc_hd__clkbuf_1 _11378_ (.A(net2204),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(net6351),
    .A1(net2656),
    .S(_04573_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_1 _11380_ (.A(net6353),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(net7211),
    .A1(net6970),
    .S(_04573_),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_1 _11382_ (.A(net2657),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(net6970),
    .A1(net6952),
    .S(_04573_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _11384_ (.A(net2512),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _11385_ (.A0(net6952),
    .A1(net2816),
    .S(_04573_),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _11386_ (.A(net6954),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(net7185),
    .A1(net6978),
    .S(_04573_),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_1 _11388_ (.A(net2817),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(net6978),
    .A1(net6732),
    .S(_04573_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_1 _11390_ (.A(net2609),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(net6732),
    .A1(net2734),
    .S(_04573_),
    .X(_04582_));
 sky130_fd_sc_hd__clkbuf_1 _11392_ (.A(net6734),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _11393_ (.A0(net7137),
    .A1(net2809),
    .S(_04573_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _11394_ (.A(net7139),
    .X(_01122_));
 sky130_fd_sc_hd__clkbuf_4 _11395_ (.A(_04242_),
    .X(_04584_));
 sky130_fd_sc_hd__mux2_1 _11396_ (.A0(net7276),
    .A1(net7219),
    .S(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _11397_ (.A(net2810),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _11398_ (.A0(net7219),
    .A1(net6333),
    .S(_04584_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _11399_ (.A(net2693),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _11400_ (.A0(net6333),
    .A1(net1620),
    .S(_04584_),
    .X(_04587_));
 sky130_fd_sc_hd__clkbuf_1 _11401_ (.A(net6335),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _11402_ (.A0(net6598),
    .A1(net2215),
    .S(_04584_),
    .X(_04588_));
 sky130_fd_sc_hd__buf_1 _11403_ (.A(net6600),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _11404_ (.A0(net7010),
    .A1(net6984),
    .S(_04584_),
    .X(_04589_));
 sky130_fd_sc_hd__clkbuf_1 _11405_ (.A(net2216),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _11406_ (.A0(net6984),
    .A1(net6461),
    .S(_04584_),
    .X(_04590_));
 sky130_fd_sc_hd__clkbuf_1 _11407_ (.A(net2409),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _11408_ (.A0(net6461),
    .A1(net2793),
    .S(_04584_),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_1 _11409_ (.A(net6463),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _11410_ (.A0(net7264),
    .A1(net6798),
    .S(_04584_),
    .X(_04592_));
 sky130_fd_sc_hd__clkbuf_1 _11411_ (.A(net2794),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _11412_ (.A0(net6798),
    .A1(net2370),
    .S(_04584_),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _11413_ (.A(net6800),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _11414_ (.A0(net6920),
    .A1(net5924),
    .S(_04584_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _11415_ (.A(net2371),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _11416_ (.A0(net5924),
    .A1(net5767),
    .S(_04243_),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_1 _11417_ (.A(net5926),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _11418_ (.A0(net5767),
    .A1(net1521),
    .S(_04243_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _11419_ (.A(net5769),
    .X(_01110_));
 sky130_fd_sc_hd__clkbuf_8 _11420_ (.A(_04241_),
    .X(_04597_));
 sky130_fd_sc_hd__buf_8 _11421_ (.A(_04597_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 _11422_ (.A(net4036),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_4 _11423_ (.A(net4037),
    .X(_04599_));
 sky130_fd_sc_hd__inv_2 _11424_ (.A(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__inv_2 _11425_ (.A(net3993),
    .Y(_04601_));
 sky130_fd_sc_hd__buf_4 _11426_ (.A(net4009),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_4 _11427_ (.A(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_4 _11428_ (.A(net3760),
    .X(_04604_));
 sky130_fd_sc_hd__inv_2 _11429_ (.A(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__inv_2 _11430_ (.A(net3908),
    .Y(_04606_));
 sky130_fd_sc_hd__nor2_1 _11431_ (.A(_04605_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__or2_2 _11432_ (.A(net4052),
    .B(_04599_),
    .X(_04608_));
 sky130_fd_sc_hd__o31a_1 _11433_ (.A1(_04164_),
    .A2(_04603_),
    .A3(_04607_),
    .B1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__xnor2_1 _11434_ (.A(_04161_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__or2_1 _11435_ (.A(_04601_),
    .B(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__nor2_1 _11436_ (.A(net4009),
    .B(_04607_),
    .Y(_04612_));
 sky130_fd_sc_hd__inv_2 _11437_ (.A(net4009),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_2 _11438_ (.A(_04604_),
    .B(net3908),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_1 _11439_ (.A(net4010),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__or2_1 _11440_ (.A(_04612_),
    .B(_04615_),
    .X(_04616_));
 sky130_fd_sc_hd__or4_1 _11441_ (.A(_04165_),
    .B(_04600_),
    .C(_04611_),
    .D(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__buf_6 _11442_ (.A(_04617_),
    .X(net73));
 sky130_fd_sc_hd__inv_2 _11443_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .Y(_04618_));
 sky130_fd_sc_hd__or2_1 _11444_ (.A(net3506),
    .B(net3534),
    .X(_04619_));
 sky130_fd_sc_hd__inv_2 _11445_ (.A(net4103),
    .Y(_04620_));
 sky130_fd_sc_hd__nand2_2 _11446_ (.A(net4104),
    .B(net89),
    .Y(_04621_));
 sky130_fd_sc_hd__inv_2 _11447_ (.A(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__buf_4 _11448_ (.A(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__buf_4 _11449_ (.A(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__o31ai_1 _11450_ (.A1(net3402),
    .A2(net2982),
    .A3(net3507),
    .B1(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__clkbuf_4 _11451_ (.A(net4930),
    .X(_04626_));
 sky130_fd_sc_hd__clkbuf_2 _11452_ (.A(net4026),
    .X(_04627_));
 sky130_fd_sc_hd__or4bb_2 _11453_ (.A(net4909),
    .B(net2982),
    .C_N(_04626_),
    .D_N(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__or2b_1 _11454_ (.A(net2982),
    .B_N(net4909),
    .X(_04629_));
 sky130_fd_sc_hd__or3b_1 _11455_ (.A(net4910),
    .B(_04626_),
    .C_N(_04627_),
    .X(_04630_));
 sky130_fd_sc_hd__nand2_1 _11456_ (.A(_04628_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__clkbuf_8 _11457_ (.A(_04621_),
    .X(_04632_));
 sky130_fd_sc_hd__buf_4 _11458_ (.A(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__o32ai_1 _11459_ (.A1(net7582),
    .A2(net3403),
    .A3(_04631_),
    .B1(_04633_),
    .B2(_04628_),
    .Y(_00001_));
 sky130_fd_sc_hd__or2_2 _11460_ (.A(_04162_),
    .B(_04611_),
    .X(_04634_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11461_ (.A(_04634_),
    .X(net72));
 sky130_fd_sc_hd__buf_4 _11462_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _11463_ (.A(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__a31o_1 _11464_ (.A1(net4947),
    .A2(_04628_),
    .A3(_04630_),
    .B1(net3403),
    .X(_00000_));
 sky130_fd_sc_hd__buf_4 _11465_ (.A(_04599_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_4 _11466_ (.A(net7317),
    .X(_04638_));
 sky130_fd_sc_hd__buf_4 _11467_ (.A(net6496),
    .X(_04639_));
 sky130_fd_sc_hd__nor2_4 _11468_ (.A(_04638_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__and2_1 _11469_ (.A(_04638_),
    .B(_04639_),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_4 _11470_ (.A(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__a22o_1 _11471_ (.A1(\rbzero.spi_registers.texadd3[14] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[14] ),
    .X(_04643_));
 sky130_fd_sc_hd__nor2b_4 _11472_ (.A(_04639_),
    .B_N(_04638_),
    .Y(_04644_));
 sky130_fd_sc_hd__a22o_1 _11473_ (.A1(\rbzero.spi_registers.texadd3[13] ),
    .A2(_04640_),
    .B1(_04644_),
    .B2(\rbzero.spi_registers.texadd1[13] ),
    .X(_04645_));
 sky130_fd_sc_hd__clkbuf_4 _11474_ (.A(net4086),
    .X(_04646_));
 sky130_fd_sc_hd__mux4_1 _11475_ (.A0(\rbzero.spi_registers.texadd3[12] ),
    .A1(\rbzero.spi_registers.texadd1[12] ),
    .A2(\rbzero.spi_registers.texadd0[12] ),
    .A3(\rbzero.spi_registers.texadd2[12] ),
    .S0(_04638_),
    .S1(_04639_),
    .X(_04647_));
 sky130_fd_sc_hd__and2_1 _11476_ (.A(_04646_),
    .B(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__mux4_1 _11477_ (.A0(\rbzero.spi_registers.texadd3[11] ),
    .A1(\rbzero.spi_registers.texadd1[11] ),
    .A2(\rbzero.spi_registers.texadd0[11] ),
    .A3(\rbzero.spi_registers.texadd2[11] ),
    .S0(_04638_),
    .S1(_04639_),
    .X(_04649_));
 sky130_fd_sc_hd__nand2_1 _11478_ (.A(\rbzero.texu_hot[5] ),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__mux4_1 _11479_ (.A0(\rbzero.spi_registers.texadd3[10] ),
    .A1(\rbzero.spi_registers.texadd1[10] ),
    .A2(\rbzero.spi_registers.texadd0[10] ),
    .A3(\rbzero.spi_registers.texadd2[10] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04651_));
 sky130_fd_sc_hd__nand2_1 _11480_ (.A(\rbzero.texu_hot[4] ),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__mux4_1 _11481_ (.A0(\rbzero.spi_registers.texadd3[9] ),
    .A1(\rbzero.spi_registers.texadd1[9] ),
    .A2(\rbzero.spi_registers.texadd0[9] ),
    .A3(\rbzero.spi_registers.texadd2[9] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04653_));
 sky130_fd_sc_hd__nand2_1 _11482_ (.A(\rbzero.texu_hot[3] ),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__mux4_1 _11483_ (.A0(\rbzero.spi_registers.texadd3[8] ),
    .A1(\rbzero.spi_registers.texadd1[8] ),
    .A2(\rbzero.spi_registers.texadd0[8] ),
    .A3(\rbzero.spi_registers.texadd2[8] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04655_));
 sky130_fd_sc_hd__nand2_1 _11484_ (.A(\rbzero.texu_hot[2] ),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__mux4_1 _11485_ (.A0(\rbzero.spi_registers.texadd3[7] ),
    .A1(\rbzero.spi_registers.texadd1[7] ),
    .A2(\rbzero.spi_registers.texadd0[7] ),
    .A3(\rbzero.spi_registers.texadd2[7] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _11486_ (.A(\rbzero.texu_hot[1] ),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__mux4_1 _11487_ (.A0(\rbzero.spi_registers.texadd3[6] ),
    .A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(\rbzero.spi_registers.texadd0[6] ),
    .A3(\rbzero.spi_registers.texadd2[6] ),
    .S0(\rbzero.wall_hot[1] ),
    .S1(\rbzero.wall_hot[0] ),
    .X(_04659_));
 sky130_fd_sc_hd__nand2_1 _11488_ (.A(\rbzero.texu_hot[0] ),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__or2_1 _11489_ (.A(\rbzero.texu_hot[1] ),
    .B(_04657_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2_1 _11490_ (.A(_04658_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__or2_1 _11491_ (.A(_04660_),
    .B(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__or2_1 _11492_ (.A(\rbzero.texu_hot[2] ),
    .B(_04655_),
    .X(_04664_));
 sky130_fd_sc_hd__nand2_1 _11493_ (.A(_04656_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__a21o_1 _11494_ (.A1(_04658_),
    .A2(_04663_),
    .B1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__or2_1 _11495_ (.A(\rbzero.texu_hot[3] ),
    .B(_04653_),
    .X(_04667_));
 sky130_fd_sc_hd__nand2_1 _11496_ (.A(_04654_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__a21o_1 _11497_ (.A1(_04656_),
    .A2(_04666_),
    .B1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__or2_1 _11498_ (.A(\rbzero.texu_hot[4] ),
    .B(_04651_),
    .X(_04670_));
 sky130_fd_sc_hd__nand2_1 _11499_ (.A(_04652_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__a21o_1 _11500_ (.A1(_04654_),
    .A2(_04669_),
    .B1(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__or2_1 _11501_ (.A(\rbzero.texu_hot[5] ),
    .B(_04649_),
    .X(_04673_));
 sky130_fd_sc_hd__nand2_1 _11502_ (.A(_04650_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__a21o_1 _11503_ (.A1(_04652_),
    .A2(_04672_),
    .B1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__nor2_1 _11504_ (.A(_04646_),
    .B(_04647_),
    .Y(_04676_));
 sky130_fd_sc_hd__or2_1 _11505_ (.A(_04648_),
    .B(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__a21oi_1 _11506_ (.A1(_04650_),
    .A2(_04675_),
    .B1(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__inv_2 _11507_ (.A(_04642_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand2b_4 _11508_ (.A_N(_04638_),
    .B(_04639_),
    .Y(_04680_));
 sky130_fd_sc_hd__inv_2 _11509_ (.A(_04645_),
    .Y(_04681_));
 sky130_fd_sc_hd__o221a_1 _11510_ (.A1(\rbzero.spi_registers.texadd2[13] ),
    .A2(_04679_),
    .B1(_04680_),
    .B2(\rbzero.spi_registers.texadd0[13] ),
    .C1(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__o21a_1 _11511_ (.A1(_04648_),
    .A2(_04678_),
    .B1(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__or2_1 _11512_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_04680_),
    .X(_04684_));
 sky130_fd_sc_hd__or3b_1 _11513_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .B(_04639_),
    .C_N(_04638_),
    .X(_04685_));
 sky130_fd_sc_hd__a22oi_2 _11514_ (.A1(\rbzero.spi_registers.texadd3[14] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[14] ),
    .Y(_04686_));
 sky130_fd_sc_hd__o2111a_1 _11515_ (.A1(_04645_),
    .A2(_04683_),
    .B1(_04684_),
    .C1(_04685_),
    .D1(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__mux4_1 _11516_ (.A0(\rbzero.spi_registers.texadd3[15] ),
    .A1(\rbzero.spi_registers.texadd1[15] ),
    .A2(\rbzero.spi_registers.texadd0[15] ),
    .A3(\rbzero.spi_registers.texadd2[15] ),
    .S0(_04638_),
    .S1(_04639_),
    .X(_04688_));
 sky130_fd_sc_hd__o21ai_1 _11517_ (.A1(_04643_),
    .A2(_04687_),
    .B1(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__mux4_1 _11518_ (.A0(\rbzero.spi_registers.texadd3[16] ),
    .A1(\rbzero.spi_registers.texadd1[16] ),
    .A2(\rbzero.spi_registers.texadd0[16] ),
    .A3(\rbzero.spi_registers.texadd2[16] ),
    .S0(_04638_),
    .S1(_04639_),
    .X(_04690_));
 sky130_fd_sc_hd__nor2b_1 _11519_ (.A(_04689_),
    .B_N(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__buf_4 _11520_ (.A(net7318),
    .X(_04692_));
 sky130_fd_sc_hd__buf_4 _11521_ (.A(net6497),
    .X(_04693_));
 sky130_fd_sc_hd__mux4_2 _11522_ (.A0(\rbzero.spi_registers.texadd3[17] ),
    .A1(\rbzero.spi_registers.texadd1[17] ),
    .A2(\rbzero.spi_registers.texadd0[17] ),
    .A3(\rbzero.spi_registers.texadd2[17] ),
    .S0(_04692_),
    .S1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__mux4_1 _11523_ (.A0(\rbzero.spi_registers.texadd3[18] ),
    .A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(\rbzero.spi_registers.texadd0[18] ),
    .A3(\rbzero.spi_registers.texadd2[18] ),
    .S0(_04692_),
    .S1(_04693_),
    .X(_04695_));
 sky130_fd_sc_hd__and3_1 _11524_ (.A(_04691_),
    .B(_04694_),
    .C(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__mux4_2 _11525_ (.A0(\rbzero.spi_registers.texadd3[19] ),
    .A1(\rbzero.spi_registers.texadd1[19] ),
    .A2(\rbzero.spi_registers.texadd0[19] ),
    .A3(\rbzero.spi_registers.texadd2[19] ),
    .S0(_04692_),
    .S1(_04693_),
    .X(_04697_));
 sky130_fd_sc_hd__mux4_1 _11526_ (.A0(\rbzero.spi_registers.texadd3[20] ),
    .A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(\rbzero.spi_registers.texadd0[20] ),
    .A3(\rbzero.spi_registers.texadd2[20] ),
    .S0(_04692_),
    .S1(_04693_),
    .X(_04698_));
 sky130_fd_sc_hd__and3_1 _11527_ (.A(_04696_),
    .B(_04697_),
    .C(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__mux4_1 _11528_ (.A0(\rbzero.spi_registers.texadd3[21] ),
    .A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(\rbzero.spi_registers.texadd0[21] ),
    .A3(\rbzero.spi_registers.texadd2[21] ),
    .S0(_04692_),
    .S1(_04693_),
    .X(_04700_));
 sky130_fd_sc_hd__nand2_1 _11529_ (.A(_04699_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__o21ba_1 _11530_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_04693_),
    .B1_N(_04692_),
    .X(_04702_));
 sky130_fd_sc_hd__a221o_1 _11531_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(_04693_),
    .B1(_04644_),
    .B2(\rbzero.spi_registers.texadd1[22] ),
    .C1(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__o21ai_1 _11532_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_04680_),
    .B1(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__and3_1 _11533_ (.A(_04160_),
    .B(_04701_),
    .C(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__or2_1 _11534_ (.A(_04701_),
    .B(_04704_),
    .X(_04706_));
 sky130_fd_sc_hd__and2b_1 _11535_ (.A_N(_04692_),
    .B(\rbzero.spi_registers.texadd3[23] ),
    .X(_04707_));
 sky130_fd_sc_hd__a221o_1 _11536_ (.A1(\rbzero.spi_registers.texadd2[23] ),
    .A2(_04642_),
    .B1(_04644_),
    .B2(\rbzero.spi_registers.texadd1[23] ),
    .C1(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__nor2b_2 _11537_ (.A(_04692_),
    .B_N(_04693_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21o_1 _11538_ (.A1(\rbzero.spi_registers.texadd0[23] ),
    .A2(_04709_),
    .B1(_04159_),
    .X(_04710_));
 sky130_fd_sc_hd__a21oi_1 _11539_ (.A1(_04680_),
    .A2(_04708_),
    .B1(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__xnor2_1 _11540_ (.A(_04706_),
    .B(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__inv_2 _11541_ (.A(net4891),
    .Y(_04713_));
 sky130_fd_sc_hd__buf_4 _11542_ (.A(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__o21a_1 _11543_ (.A1(_04705_),
    .A2(_04712_),
    .B1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__or2_1 _11544_ (.A(_04699_),
    .B(_04700_),
    .X(_04716_));
 sky130_fd_sc_hd__nand2_1 _11545_ (.A(_04701_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__buf_4 _11546_ (.A(net4891),
    .X(_04718_));
 sky130_fd_sc_hd__inv_2 _11547_ (.A(net3868),
    .Y(_04719_));
 sky130_fd_sc_hd__nand2_1 _11548_ (.A(_04718_),
    .B(net3869),
    .Y(_04720_));
 sky130_fd_sc_hd__inv_2 _11549_ (.A(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__a21oi_1 _11550_ (.A1(_04696_),
    .A2(_04697_),
    .B1(_04698_),
    .Y(_04722_));
 sky130_fd_sc_hd__or2_1 _11551_ (.A(_04699_),
    .B(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__clkbuf_4 _11552_ (.A(net3869),
    .X(_04724_));
 sky130_fd_sc_hd__nor2_2 _11553_ (.A(_04714_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__buf_4 _11554_ (.A(net6049),
    .X(_04726_));
 sky130_fd_sc_hd__buf_4 _11555_ (.A(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__a221o_1 _11556_ (.A1(_04717_),
    .A2(_04721_),
    .B1(_04723_),
    .B2(_04725_),
    .C1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__or2_1 _11557_ (.A(_04696_),
    .B(_04697_),
    .X(_04729_));
 sky130_fd_sc_hd__nand2_1 _11558_ (.A(_04696_),
    .B(_04697_),
    .Y(_04730_));
 sky130_fd_sc_hd__a21o_1 _11559_ (.A1(_04691_),
    .A2(_04694_),
    .B1(_04695_),
    .X(_04731_));
 sky130_fd_sc_hd__nor2_1 _11560_ (.A(_04724_),
    .B(_04696_),
    .Y(_04732_));
 sky130_fd_sc_hd__a32o_1 _11561_ (.A1(_04724_),
    .A2(_04729_),
    .A3(_04730_),
    .B1(_04731_),
    .B2(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__or2_1 _11562_ (.A(_04691_),
    .B(_04694_),
    .X(_04734_));
 sky130_fd_sc_hd__nand2_1 _11563_ (.A(_04691_),
    .B(_04694_),
    .Y(_04735_));
 sky130_fd_sc_hd__and2b_1 _11564_ (.A_N(_04690_),
    .B(_04689_),
    .X(_04736_));
 sky130_fd_sc_hd__o31ai_1 _11565_ (.A1(_04724_),
    .A2(_04736_),
    .A3(_04691_),
    .B1(_04718_),
    .Y(_04737_));
 sky130_fd_sc_hd__a31o_1 _11566_ (.A1(_04724_),
    .A2(_04734_),
    .A3(_04735_),
    .B1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__o211a_1 _11567_ (.A1(_04718_),
    .A2(_04733_),
    .B1(_04738_),
    .C1(_04727_),
    .X(_04739_));
 sky130_fd_sc_hd__o21bai_2 _11568_ (.A1(_04715_),
    .A2(_04728_),
    .B1_N(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__or3_1 _11569_ (.A(_04643_),
    .B(_04687_),
    .C(_04688_),
    .X(_04741_));
 sky130_fd_sc_hd__nor2_1 _11570_ (.A(_04714_),
    .B(_04683_),
    .Y(_04742_));
 sky130_fd_sc_hd__o31a_1 _11571_ (.A1(_04648_),
    .A2(_04678_),
    .A3(_04682_),
    .B1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__a311o_1 _11572_ (.A1(_04714_),
    .A2(_04689_),
    .A3(_04741_),
    .B1(_04743_),
    .C1(_04160_),
    .X(_04744_));
 sky130_fd_sc_hd__and3_1 _11573_ (.A(_04677_),
    .B(_04650_),
    .C(_04675_),
    .X(_04745_));
 sky130_fd_sc_hd__a311o_1 _11574_ (.A1(_04686_),
    .A2(_04684_),
    .A3(_04685_),
    .B1(_04645_),
    .C1(_04683_),
    .X(_04746_));
 sky130_fd_sc_hd__or3b_1 _11575_ (.A(_04718_),
    .B(_04687_),
    .C_N(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__o311a_1 _11576_ (.A1(_04714_),
    .A2(_04678_),
    .A3(_04745_),
    .B1(_04747_),
    .C1(_04160_),
    .X(_04748_));
 sky130_fd_sc_hd__nor2_1 _11577_ (.A(_04727_),
    .B(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__nand3_1 _11578_ (.A(_04671_),
    .B(_04654_),
    .C(_04669_),
    .Y(_04750_));
 sky130_fd_sc_hd__nand3_1 _11579_ (.A(_04674_),
    .B(_04652_),
    .C(_04672_),
    .Y(_04751_));
 sky130_fd_sc_hd__and3_1 _11580_ (.A(_04724_),
    .B(_04675_),
    .C(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__a311o_1 _11581_ (.A1(_04160_),
    .A2(_04672_),
    .A3(_04750_),
    .B1(_04752_),
    .C1(_04718_),
    .X(_04753_));
 sky130_fd_sc_hd__nand3_1 _11582_ (.A(_04656_),
    .B(_04666_),
    .C(_04668_),
    .Y(_04754_));
 sky130_fd_sc_hd__and3_1 _11583_ (.A(_04724_),
    .B(_04669_),
    .C(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__nand3_1 _11584_ (.A(_04665_),
    .B(_04658_),
    .C(_04663_),
    .Y(_04756_));
 sky130_fd_sc_hd__a31o_1 _11585_ (.A1(_04159_),
    .A2(_04666_),
    .A3(_04756_),
    .B1(_04714_),
    .X(_04757_));
 sky130_fd_sc_hd__o21a_1 _11586_ (.A1(_04755_),
    .A2(_04757_),
    .B1(_04727_),
    .X(_04758_));
 sky130_fd_sc_hd__clkbuf_4 _11587_ (.A(_04604_),
    .X(_04759_));
 sky130_fd_sc_hd__buf_4 _11588_ (.A(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__a221o_1 _11589_ (.A1(_04744_),
    .A2(_04749_),
    .B1(_04753_),
    .B2(_04758_),
    .C1(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__a21o_1 _11590_ (.A1(\rbzero.spi_registers.texadd1[3] ),
    .A2(_04644_),
    .B1(_04709_),
    .X(_04762_));
 sky130_fd_sc_hd__a22o_1 _11591_ (.A1(\rbzero.spi_registers.texadd3[3] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[3] ),
    .X(_04763_));
 sky130_fd_sc_hd__o221a_1 _11592_ (.A1(\rbzero.spi_registers.texadd0[3] ),
    .A2(_04680_),
    .B1(_04762_),
    .B2(_04763_),
    .C1(_04724_),
    .X(_04764_));
 sky130_fd_sc_hd__a21o_1 _11593_ (.A1(\rbzero.spi_registers.texadd1[2] ),
    .A2(_04644_),
    .B1(_04709_),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_1 _11594_ (.A1(\rbzero.spi_registers.texadd3[2] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[2] ),
    .X(_04766_));
 sky130_fd_sc_hd__o221a_1 _11595_ (.A1(\rbzero.spi_registers.texadd0[2] ),
    .A2(_04680_),
    .B1(_04765_),
    .B2(_04766_),
    .C1(_04159_),
    .X(_04767_));
 sky130_fd_sc_hd__o31a_1 _11596_ (.A1(_04718_),
    .A2(_04764_),
    .A3(_04767_),
    .B1(_04727_),
    .X(_04768_));
 sky130_fd_sc_hd__a22o_1 _11597_ (.A1(\rbzero.spi_registers.texadd3[0] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[0] ),
    .X(_04769_));
 sky130_fd_sc_hd__a21o_1 _11598_ (.A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(_04644_),
    .B1(_04709_),
    .X(_04770_));
 sky130_fd_sc_hd__o221a_1 _11599_ (.A1(\rbzero.spi_registers.texadd0[0] ),
    .A2(_04680_),
    .B1(_04769_),
    .B2(_04770_),
    .C1(_04159_),
    .X(_04771_));
 sky130_fd_sc_hd__a22o_1 _11600_ (.A1(\rbzero.spi_registers.texadd3[1] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[1] ),
    .X(_04772_));
 sky130_fd_sc_hd__a21o_1 _11601_ (.A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(_04644_),
    .B1(_04709_),
    .X(_04773_));
 sky130_fd_sc_hd__o221a_1 _11602_ (.A1(\rbzero.spi_registers.texadd0[1] ),
    .A2(_04680_),
    .B1(_04772_),
    .B2(_04773_),
    .C1(_04724_),
    .X(_04774_));
 sky130_fd_sc_hd__or3_1 _11603_ (.A(_04714_),
    .B(_04771_),
    .C(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__clkbuf_4 _11604_ (.A(net6025),
    .X(_04776_));
 sky130_fd_sc_hd__buf_4 _11605_ (.A(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__nand2_1 _11606_ (.A(_04660_),
    .B(_04662_),
    .Y(_04778_));
 sky130_fd_sc_hd__or2_1 _11607_ (.A(\rbzero.texu_hot[0] ),
    .B(_04659_),
    .X(_04779_));
 sky130_fd_sc_hd__and3_1 _11608_ (.A(_04159_),
    .B(_04660_),
    .C(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__a31o_1 _11609_ (.A1(_04724_),
    .A2(_04663_),
    .A3(_04778_),
    .B1(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__a22o_1 _11610_ (.A1(\rbzero.spi_registers.texadd1[5] ),
    .A2(_04644_),
    .B1(_04709_),
    .B2(\rbzero.spi_registers.texadd0[5] ),
    .X(_04782_));
 sky130_fd_sc_hd__a221o_1 _11611_ (.A1(\rbzero.spi_registers.texadd3[5] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[5] ),
    .C1(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__a22o_1 _11612_ (.A1(\rbzero.spi_registers.texadd1[4] ),
    .A2(_04644_),
    .B1(_04709_),
    .B2(\rbzero.spi_registers.texadd0[4] ),
    .X(_04784_));
 sky130_fd_sc_hd__a22o_1 _11613_ (.A1(\rbzero.spi_registers.texadd3[4] ),
    .A2(_04640_),
    .B1(_04642_),
    .B2(\rbzero.spi_registers.texadd2[4] ),
    .X(_04785_));
 sky130_fd_sc_hd__o21a_1 _11614_ (.A1(_04784_),
    .A2(_04785_),
    .B1(_04725_),
    .X(_04786_));
 sky130_fd_sc_hd__a221o_1 _11615_ (.A1(_04714_),
    .A2(_04781_),
    .B1(_04783_),
    .B2(_04721_),
    .C1(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__and2b_1 _11616_ (.A_N(_04727_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__a211o_1 _11617_ (.A1(_04768_),
    .A2(_04775_),
    .B1(_04777_),
    .C1(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__or2_2 _11618_ (.A(_04759_),
    .B(_04776_),
    .X(_04790_));
 sky130_fd_sc_hd__and3_1 _11619_ (.A(_04637_),
    .B(_04614_),
    .C(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__a31o_1 _11620_ (.A1(_04761_),
    .A2(_04789_),
    .A3(_04791_),
    .B1(_04613_),
    .X(_04792_));
 sky130_fd_sc_hd__a41o_1 _11621_ (.A1(_04637_),
    .A2(_04605_),
    .A3(_04606_),
    .A4(_04740_),
    .B1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__a21oi_1 _11622_ (.A1(_04614_),
    .A2(_04790_),
    .B1(_04160_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _11623_ (.A(_04714_),
    .B(_04160_),
    .Y(_04795_));
 sky130_fd_sc_hd__o21ai_1 _11624_ (.A1(_04727_),
    .A2(_04721_),
    .B1(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__o31a_1 _11625_ (.A1(_04727_),
    .A2(_04718_),
    .A3(_04794_),
    .B1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__o21ai_1 _11626_ (.A1(_04614_),
    .A2(_04797_),
    .B1(_04613_),
    .Y(_04798_));
 sky130_fd_sc_hd__and3b_1 _11627_ (.A_N(net73),
    .B(_04793_),
    .C(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__buf_2 _11628_ (.A(_04799_),
    .X(net74));
 sky130_fd_sc_hd__buf_1 _11629_ (.A(clknet_leaf_66_i_clk),
    .X(_04800_));
 sky130_fd_sc_hd__inv_2 _11630__1 (.A(clknet_1_0__leaf__04800_),
    .Y(net140));
 sky130_fd_sc_hd__buf_4 _11631_ (.A(net4971),
    .X(_04801_));
 sky130_fd_sc_hd__buf_4 _11632_ (.A(net4972),
    .X(_04802_));
 sky130_fd_sc_hd__or3_1 _11633_ (.A(net4020),
    .B(net3897),
    .C(net3964),
    .X(_04803_));
 sky130_fd_sc_hd__clkbuf_1 _11634_ (.A(net4099),
    .X(_04804_));
 sky130_fd_sc_hd__clkbuf_1 _11635_ (.A(net4032),
    .X(_04805_));
 sky130_fd_sc_hd__or2_1 _11636_ (.A(net4033),
    .B(net4013),
    .X(_04806_));
 sky130_fd_sc_hd__or2_1 _11637_ (.A(net4059),
    .B(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__or2_1 _11638_ (.A(_04803_),
    .B(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__or4b_1 _11639_ (.A(net3936),
    .B(net3929),
    .C(net4001),
    .D_N(net3),
    .X(_04809_));
 sky130_fd_sc_hd__and3_1 _11640_ (.A(net3987),
    .B(net2986),
    .C(net3868),
    .X(_04810_));
 sky130_fd_sc_hd__clkbuf_2 _11641_ (.A(net3988),
    .X(_04811_));
 sky130_fd_sc_hd__and2_1 _11642_ (.A(net6025),
    .B(net3989),
    .X(_04812_));
 sky130_fd_sc_hd__or2_1 _11643_ (.A(net3760),
    .B(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__o211a_1 _11644_ (.A1(net4009),
    .A2(net3761),
    .B1(net4052),
    .C1(net4037),
    .X(_04814_));
 sky130_fd_sc_hd__a21oi_1 _11645_ (.A1(net4004),
    .A2(_04814_),
    .B1(net3992),
    .Y(_04815_));
 sky130_fd_sc_hd__a211oi_2 _11646_ (.A1(_04802_),
    .A2(_04808_),
    .B1(_04809_),
    .C1(net7362),
    .Y(_04816_));
 sky130_fd_sc_hd__inv_2 _11647_ (.A(net2),
    .Y(_04817_));
 sky130_fd_sc_hd__nand2_4 _11648_ (.A(net4909),
    .B(net6168),
    .Y(_04818_));
 sky130_fd_sc_hd__nand2_1 _11649_ (.A(net4930),
    .B(net4026),
    .Y(_04819_));
 sky130_fd_sc_hd__o21a_1 _11650_ (.A1(_04818_),
    .A2(net3535),
    .B1(net2),
    .X(_04820_));
 sky130_fd_sc_hd__inv_2 _11651_ (.A(net4001),
    .Y(_04821_));
 sky130_fd_sc_hd__inv_2 _11652_ (.A(net3893),
    .Y(_04822_));
 sky130_fd_sc_hd__inv_2 _11653_ (.A(net4090),
    .Y(_04823_));
 sky130_fd_sc_hd__a22o_1 _11654_ (.A1(_04801_),
    .A2(_04822_),
    .B1(_04823_),
    .B2(_04602_),
    .X(_04824_));
 sky130_fd_sc_hd__a221o_1 _11655_ (.A1(_04821_),
    .A2(net3279),
    .B1(net4090),
    .B2(net4010),
    .C1(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__inv_2 _11656_ (.A(net3921),
    .Y(_04826_));
 sky130_fd_sc_hd__inv_2 _11657_ (.A(net3279),
    .Y(_04827_));
 sky130_fd_sc_hd__inv_2 _11658_ (.A(net3995),
    .Y(_04828_));
 sky130_fd_sc_hd__a22o_1 _11659_ (.A1(net4001),
    .A2(_04827_),
    .B1(net3996),
    .B2(_04759_),
    .X(_04829_));
 sky130_fd_sc_hd__a221o_1 _11660_ (.A1(_04826_),
    .A2(_04599_),
    .B1(_04605_),
    .B2(net3995),
    .C1(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__buf_4 _11661_ (.A(net6330),
    .X(_04831_));
 sky130_fd_sc_hd__xor2_1 _11662_ (.A(_04831_),
    .B(net3917),
    .X(_04832_));
 sky130_fd_sc_hd__xor2_1 _11663_ (.A(net4059),
    .B(net4387),
    .X(_04833_));
 sky130_fd_sc_hd__xor2_1 _11664_ (.A(net3853),
    .B(net4052),
    .X(_04834_));
 sky130_fd_sc_hd__a221o_1 _11665_ (.A1(net3921),
    .A2(_04600_),
    .B1(_04606_),
    .B2(net3821),
    .C1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__inv_2 _11666_ (.A(net4971),
    .Y(_04836_));
 sky130_fd_sc_hd__inv_2 _11667_ (.A(net3821),
    .Y(_04837_));
 sky130_fd_sc_hd__xor2_1 _11668_ (.A(net4033),
    .B(net3880),
    .X(_04838_));
 sky130_fd_sc_hd__a221o_1 _11669_ (.A1(_04836_),
    .A2(net3893),
    .B1(_04837_),
    .B2(_04776_),
    .C1(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__or4_1 _11670_ (.A(_04832_),
    .B(_04833_),
    .C(_04835_),
    .D(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__or3_1 _11671_ (.A(net4091),
    .B(_04830_),
    .C(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__inv_2 _11672_ (.A(net4092),
    .Y(_04842_));
 sky130_fd_sc_hd__inv_2 _11673_ (.A(net3964),
    .Y(_04843_));
 sky130_fd_sc_hd__xnor2_1 _11674_ (.A(net4020),
    .B(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_04844_));
 sky130_fd_sc_hd__o221a_1 _11675_ (.A1(_04843_),
    .A2(net4063),
    .B1(net3028),
    .B2(_04714_),
    .C1(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__inv_2 _11676_ (.A(net4105),
    .Y(_04846_));
 sky130_fd_sc_hd__inv_2 _11677_ (.A(net3028),
    .Y(_04847_));
 sky130_fd_sc_hd__xnor2_1 _11678_ (.A(net3008),
    .B(net4049),
    .Y(_04848_));
 sky130_fd_sc_hd__o221a_1 _11679_ (.A1(_04846_),
    .A2(_04726_),
    .B1(net2986),
    .B2(_04847_),
    .C1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__xor2_1 _11680_ (.A(net3897),
    .B(net4358),
    .X(_04850_));
 sky130_fd_sc_hd__a221oi_1 _11681_ (.A1(_04843_),
    .A2(net4063),
    .B1(_04846_),
    .B2(_04726_),
    .C1(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__nor2_1 _11682_ (.A(_04599_),
    .B(_04602_),
    .Y(_04852_));
 sky130_fd_sc_hd__or3b_1 _11683_ (.A(_04164_),
    .B(_04790_),
    .C_N(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__or3_1 _11684_ (.A(_04726_),
    .B(net4891),
    .C(net3868),
    .X(_04854_));
 sky130_fd_sc_hd__or2_1 _11685_ (.A(_04853_),
    .B(net2987),
    .X(_04855_));
 sky130_fd_sc_hd__or3_1 _11686_ (.A(net4001),
    .B(net4972),
    .C(_04808_),
    .X(_04856_));
 sky130_fd_sc_hd__or3b_1 _11687_ (.A(net3936),
    .B(net3992),
    .C_N(net1),
    .X(_04857_));
 sky130_fd_sc_hd__a221o_2 _11688_ (.A1(_04161_),
    .A2(_04855_),
    .B1(_04856_),
    .B2(net3929),
    .C1(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__a41o_1 _11689_ (.A1(_04842_),
    .A2(net4064),
    .A3(_04849_),
    .A4(_04851_),
    .B1(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__inv_2 _11690_ (.A(net2705),
    .Y(_04860_));
 sky130_fd_sc_hd__xor2_1 _11691_ (.A(net2677),
    .B(_04776_),
    .X(_04861_));
 sky130_fd_sc_hd__a221o_1 _11692_ (.A1(_04821_),
    .A2(net2823),
    .B1(_04860_),
    .B2(_04759_),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__inv_2 _11693_ (.A(net2043),
    .Y(_04863_));
 sky130_fd_sc_hd__or2_1 _11694_ (.A(net4033),
    .B(net2905),
    .X(_04864_));
 sky130_fd_sc_hd__nand2_1 _11695_ (.A(net4033),
    .B(net2905),
    .Y(_04865_));
 sky130_fd_sc_hd__nand2_1 _11696_ (.A(_04801_),
    .B(net2536),
    .Y(_04866_));
 sky130_fd_sc_hd__or2_1 _11697_ (.A(net4971),
    .B(net2536),
    .X(_04867_));
 sky130_fd_sc_hd__inv_2 _11698_ (.A(net2917),
    .Y(_04868_));
 sky130_fd_sc_hd__a22o_1 _11699_ (.A1(net2043),
    .A2(_04600_),
    .B1(_04602_),
    .B2(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__a221o_1 _11700_ (.A1(_04864_),
    .A2(_04865_),
    .B1(_04866_),
    .B2(_04867_),
    .C1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__a221o_1 _11701_ (.A1(_04863_),
    .A2(_04599_),
    .B1(net4010),
    .B2(net2917),
    .C1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__or2_1 _11702_ (.A(net2839),
    .B(_04164_),
    .X(_04872_));
 sky130_fd_sc_hd__nand2_1 _11703_ (.A(net2839),
    .B(_04164_),
    .Y(_04873_));
 sky130_fd_sc_hd__or2_1 _11704_ (.A(_04831_),
    .B(net2925),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _11705_ (.A(_04831_),
    .B(net2925),
    .Y(_04875_));
 sky130_fd_sc_hd__inv_2 _11706_ (.A(net2823),
    .Y(_04876_));
 sky130_fd_sc_hd__xor2_1 _11707_ (.A(net4059),
    .B(net2864),
    .X(_04877_));
 sky130_fd_sc_hd__a221o_1 _11708_ (.A1(net4001),
    .A2(_04876_),
    .B1(net2705),
    .B2(_04605_),
    .C1(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__a221o_1 _11709_ (.A1(_04872_),
    .A2(_04873_),
    .B1(_04874_),
    .B2(_04875_),
    .C1(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__or3_1 _11710_ (.A(_04862_),
    .B(_04871_),
    .C(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__inv_2 _11711_ (.A(net4059),
    .Y(_04881_));
 sky130_fd_sc_hd__a22o_1 _11712_ (.A1(_04821_),
    .A2(net2726),
    .B1(net2789),
    .B2(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__inv_2 _11713_ (.A(net2791),
    .Y(_04883_));
 sky130_fd_sc_hd__xnor2_1 _11714_ (.A(net4033),
    .B(net2879),
    .Y(_04884_));
 sky130_fd_sc_hd__o221a_1 _11715_ (.A1(_04801_),
    .A2(_04883_),
    .B1(net2789),
    .B2(_04881_),
    .C1(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__inv_2 _11716_ (.A(net2802),
    .Y(_04886_));
 sky130_fd_sc_hd__or4_1 _11717_ (.A(net2791),
    .B(net2789),
    .C(net2879),
    .D(net2802),
    .X(_04887_));
 sky130_fd_sc_hd__o21a_1 _11718_ (.A1(net1506),
    .A2(_04887_),
    .B1(_04821_),
    .X(_04888_));
 sky130_fd_sc_hd__clkinv_4 _11719_ (.A(net4013),
    .Y(_04889_));
 sky130_fd_sc_hd__o22a_1 _11720_ (.A1(_04836_),
    .A2(net2791),
    .B1(net2802),
    .B2(net4014),
    .X(_04890_));
 sky130_fd_sc_hd__o221a_1 _11721_ (.A1(_04831_),
    .A2(_04886_),
    .B1(_04888_),
    .B2(net2726),
    .C1(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__and3b_1 _11722_ (.A_N(_04882_),
    .B(_04885_),
    .C(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__inv_2 _11723_ (.A(net3619),
    .Y(_04893_));
 sky130_fd_sc_hd__inv_2 _11724_ (.A(net2895),
    .Y(_04894_));
 sky130_fd_sc_hd__inv_2 _11725_ (.A(net2774),
    .Y(_04895_));
 sky130_fd_sc_hd__xnor2_1 _11726_ (.A(net2825),
    .B(_04602_),
    .Y(_04896_));
 sky130_fd_sc_hd__o221a_1 _11727_ (.A1(_04894_),
    .A2(_04759_),
    .B1(_04776_),
    .B2(_04895_),
    .C1(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__inv_2 _11728_ (.A(net4345),
    .Y(_04898_));
 sky130_fd_sc_hd__or4_1 _11729_ (.A(net4345),
    .B(net2825),
    .C(net2895),
    .D(net2774),
    .X(_04899_));
 sky130_fd_sc_hd__o21a_1 _11730_ (.A1(net1185),
    .A2(_04899_),
    .B1(net3620),
    .X(_04900_));
 sky130_fd_sc_hd__o22a_1 _11731_ (.A1(net4345),
    .A2(_04600_),
    .B1(_04606_),
    .B2(net2774),
    .X(_04901_));
 sky130_fd_sc_hd__o221a_1 _11732_ (.A1(_04898_),
    .A2(_04599_),
    .B1(_04900_),
    .B2(_04164_),
    .C1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__nand2_1 _11733_ (.A(_04897_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__a221o_1 _11734_ (.A1(net3620),
    .A2(_04164_),
    .B1(_04759_),
    .B2(_04894_),
    .C1(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _11735_ (.A(_04892_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__and2_1 _11736_ (.A(_04803_),
    .B(net2987),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_1 _11737_ (.A(net4092),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__a21oi_1 _11738_ (.A1(_04880_),
    .A2(_04905_),
    .B1(net4093),
    .Y(_04908_));
 sky130_fd_sc_hd__inv_2 _11739_ (.A(net42),
    .Y(_04909_));
 sky130_fd_sc_hd__nand2_2 _11740_ (.A(net1257),
    .B(net2158),
    .Y(_04910_));
 sky130_fd_sc_hd__xnor2_2 _11741_ (.A(net1500),
    .B(net2968),
    .Y(_04911_));
 sky130_fd_sc_hd__xnor2_4 _11742_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__or2_1 _11743_ (.A(net1257),
    .B(net2158),
    .X(_04913_));
 sky130_fd_sc_hd__nand2_1 _11744_ (.A(_04910_),
    .B(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__or2_1 _11745_ (.A(net1060),
    .B(net1915),
    .X(_04915_));
 sky130_fd_sc_hd__nand2_1 _11746_ (.A(net1060),
    .B(net1915),
    .Y(_04916_));
 sky130_fd_sc_hd__a21boi_1 _11747_ (.A1(net2931),
    .A2(_04915_),
    .B1_N(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__nand2_1 _11748_ (.A(net785),
    .B(net2467),
    .Y(_04918_));
 sky130_fd_sc_hd__or2_1 _11749_ (.A(net785),
    .B(net2467),
    .X(_04919_));
 sky130_fd_sc_hd__nand3_1 _11750_ (.A(net2909),
    .B(_04918_),
    .C(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__a21o_1 _11751_ (.A1(_04918_),
    .A2(_04919_),
    .B1(net2909),
    .X(_04921_));
 sky130_fd_sc_hd__nand2_1 _11752_ (.A(_04920_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_1 _11753_ (.A(net757),
    .B(net2194),
    .Y(_04923_));
 sky130_fd_sc_hd__or2_1 _11754_ (.A(net757),
    .B(net2194),
    .X(_04924_));
 sky130_fd_sc_hd__nand3_1 _11755_ (.A(net1504),
    .B(_04923_),
    .C(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__nand3_1 _11756_ (.A(_04922_),
    .B(_04923_),
    .C(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__a21o_1 _11757_ (.A1(_04923_),
    .A2(_04924_),
    .B1(net1504),
    .X(_04927_));
 sky130_fd_sc_hd__nand2_1 _11758_ (.A(_04925_),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__and2_1 _11759_ (.A(net923),
    .B(net1569),
    .X(_04929_));
 sky130_fd_sc_hd__nor2_1 _11760_ (.A(net923),
    .B(net1569),
    .Y(_04930_));
 sky130_fd_sc_hd__nor2_1 _11761_ (.A(_04929_),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__a21oi_1 _11762_ (.A1(net2776),
    .A2(_04931_),
    .B1(_04929_),
    .Y(_04932_));
 sky130_fd_sc_hd__xnor2_1 _11763_ (.A(_04928_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2_1 _11764_ (.A(net869),
    .B(net1529),
    .Y(_04934_));
 sky130_fd_sc_hd__or2_1 _11765_ (.A(net869),
    .B(net1529),
    .X(_04935_));
 sky130_fd_sc_hd__nand3_1 _11766_ (.A(net1583),
    .B(_04934_),
    .C(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__xnor2_1 _11767_ (.A(net2776),
    .B(_04931_),
    .Y(_04937_));
 sky130_fd_sc_hd__a21oi_1 _11768_ (.A1(_04934_),
    .A2(_04936_),
    .B1(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21o_1 _11769_ (.A1(_04934_),
    .A2(_04935_),
    .B1(net1583),
    .X(_04939_));
 sky130_fd_sc_hd__nand2_1 _11770_ (.A(_04936_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__or2_1 _11771_ (.A(net1010),
    .B(net1650),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _11772_ (.A(net1010),
    .B(net1650),
    .Y(_04942_));
 sky130_fd_sc_hd__a21boi_1 _11773_ (.A1(net1886),
    .A2(_04941_),
    .B1_N(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__nor2_1 _11774_ (.A(_04940_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__xnor2_1 _11775_ (.A(_04940_),
    .B(_04943_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _11776_ (.A(_04942_),
    .B(_04941_),
    .Y(_04946_));
 sky130_fd_sc_hd__xor2_1 _11777_ (.A(net1886),
    .B(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__o211a_1 _11778_ (.A1(net1072),
    .A2(net1456),
    .B1(net1166),
    .C1(net700),
    .X(_04948_));
 sky130_fd_sc_hd__a22o_1 _11779_ (.A1(net924),
    .A2(net1364),
    .B1(net1456),
    .B2(net1072),
    .X(_04949_));
 sky130_fd_sc_hd__nor2_1 _11780_ (.A(_04948_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nor2_1 _11781_ (.A(net924),
    .B(net1364),
    .Y(_04951_));
 sky130_fd_sc_hd__or3_2 _11782_ (.A(_04947_),
    .B(_04950_),
    .C(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__nor2_2 _11783_ (.A(_04945_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__and3_1 _11784_ (.A(_04937_),
    .B(_04934_),
    .C(_04936_),
    .X(_04954_));
 sky130_fd_sc_hd__or2_1 _11785_ (.A(_04938_),
    .B(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__inv_2 _11786_ (.A(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__o21a_1 _11787_ (.A1(_04944_),
    .A2(_04953_),
    .B1(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__nor2_1 _11788_ (.A(_04938_),
    .B(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__nor2_1 _11789_ (.A(_04933_),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__o21bai_1 _11790_ (.A1(_04928_),
    .A2(_04932_),
    .B1_N(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__a21oi_1 _11791_ (.A1(_04923_),
    .A2(_04925_),
    .B1(_04922_),
    .Y(_04961_));
 sky130_fd_sc_hd__a21o_1 _11792_ (.A1(_04926_),
    .A2(_04960_),
    .B1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_04915_),
    .B(_04916_),
    .Y(_04963_));
 sky130_fd_sc_hd__xor2_1 _11794_ (.A(net2931),
    .B(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__nand3_1 _11795_ (.A(_04964_),
    .B(_04918_),
    .C(_04920_),
    .Y(_04965_));
 sky130_fd_sc_hd__a21oi_1 _11796_ (.A1(_04918_),
    .A2(_04920_),
    .B1(_04964_),
    .Y(_04966_));
 sky130_fd_sc_hd__a21oi_1 _11797_ (.A1(_04962_),
    .A2(_04965_),
    .B1(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21o_1 _11798_ (.A1(_04914_),
    .A2(_04917_),
    .B1(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__o21a_1 _11799_ (.A1(_04914_),
    .A2(_04917_),
    .B1(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__xnor2_4 _11800_ (.A(_04912_),
    .B(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__nor2_4 _11801_ (.A(net3026),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__and2b_1 _11802_ (.A_N(_04966_),
    .B(_04965_),
    .X(_04972_));
 sky130_fd_sc_hd__xnor2_1 _11803_ (.A(_04962_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__or2_1 _11804_ (.A(_04971_),
    .B(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__clkbuf_8 _11805_ (.A(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__and2_1 _11806_ (.A(_04933_),
    .B(_04958_),
    .X(_04976_));
 sky130_fd_sc_hd__nor3_2 _11807_ (.A(_04959_),
    .B(_04971_),
    .C(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__buf_6 _11808_ (.A(net81),
    .X(_04978_));
 sky130_fd_sc_hd__clkbuf_8 _11809_ (.A(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__and2_1 _11810_ (.A(_04945_),
    .B(_04952_),
    .X(_04980_));
 sky130_fd_sc_hd__or3_4 _11811_ (.A(_04953_),
    .B(_04971_),
    .C(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__clkbuf_8 _11812_ (.A(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__buf_2 _11813_ (.A(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_4 _11814_ (.A(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__o21ai_2 _11815_ (.A1(_04950_),
    .A2(_04951_),
    .B1(_04947_),
    .Y(_04985_));
 sky130_fd_sc_hd__o211ai_4 _11816_ (.A1(net3026),
    .A2(_04970_),
    .B1(_04985_),
    .C1(_04952_),
    .Y(_04986_));
 sky130_fd_sc_hd__buf_4 _11817_ (.A(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__buf_4 _11818_ (.A(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__buf_4 _11819_ (.A(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__nor3_4 _11821_ (.A(_04953_),
    .B(_04971_),
    .C(_04980_),
    .Y(_04991_));
 sky130_fd_sc_hd__buf_4 _11822_ (.A(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__clkbuf_8 _11823_ (.A(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__buf_4 _11824_ (.A(_04987_),
    .X(_04994_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__or2_1 _11826_ (.A(_04993_),
    .B(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__nor3_1 _11827_ (.A(_04956_),
    .B(_04944_),
    .C(_04953_),
    .Y(_04997_));
 sky130_fd_sc_hd__or3_1 _11828_ (.A(_04957_),
    .B(_04971_),
    .C(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__clkbuf_8 _11829_ (.A(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__buf_4 _11830_ (.A(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__o211a_1 _11831_ (.A1(_04984_),
    .A2(_04990_),
    .B1(_04996_),
    .C1(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__clkbuf_8 _11832_ (.A(_04992_),
    .X(_05002_));
 sky130_fd_sc_hd__buf_4 _11833_ (.A(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__buf_4 _11834_ (.A(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _11835_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04989_),
    .X(_05005_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04988_),
    .X(_05006_));
 sky130_fd_sc_hd__or2_1 _11837_ (.A(_04983_),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__nor3_2 _11838_ (.A(_04957_),
    .B(_04971_),
    .C(_04997_),
    .Y(_05008_));
 sky130_fd_sc_hd__buf_6 _11839_ (.A(net80),
    .X(_05009_));
 sky130_fd_sc_hd__buf_4 _11840_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__o211a_1 _11841_ (.A1(_05004_),
    .A2(_05005_),
    .B1(_05007_),
    .C1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04988_),
    .X(_05012_));
 sky130_fd_sc_hd__or2_1 _11843_ (.A(_04983_),
    .B(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__clkbuf_8 _11844_ (.A(_04987_),
    .X(_05014_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__o21a_1 _11846_ (.A1(_05003_),
    .A2(_05015_),
    .B1(_04999_),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04994_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04994_),
    .X(_05018_));
 sky130_fd_sc_hd__clkbuf_8 _11849_ (.A(_04982_),
    .X(_05019_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(_05017_),
    .A1(_05018_),
    .S(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__or3_1 _11851_ (.A(_04959_),
    .B(_04971_),
    .C(_04976_),
    .X(_05021_));
 sky130_fd_sc_hd__buf_4 _11852_ (.A(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__clkbuf_8 _11853_ (.A(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__a221o_1 _11854_ (.A1(_05013_),
    .A2(_05016_),
    .B1(_05020_),
    .B2(_05010_),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__and2b_1 _11855_ (.A_N(_04961_),
    .B(_04926_),
    .X(_05025_));
 sky130_fd_sc_hd__xnor2_1 _11856_ (.A(_04960_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__or2_4 _11857_ (.A(_04971_),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_8 _11858_ (.A(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__o311a_1 _11859_ (.A1(_04979_),
    .A2(_05001_),
    .A3(_05011_),
    .B1(_05024_),
    .C1(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__clkbuf_8 _11860_ (.A(_05022_),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04989_),
    .X(_05031_));
 sky130_fd_sc_hd__mux2_1 _11862_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04988_),
    .X(_05032_));
 sky130_fd_sc_hd__or2_1 _11863_ (.A(_05003_),
    .B(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__buf_4 _11864_ (.A(_04999_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_8 _11865_ (.A(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__o211a_1 _11866_ (.A1(_04984_),
    .A2(_05031_),
    .B1(_05033_),
    .C1(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__buf_4 _11867_ (.A(_05014_),
    .X(_05037_));
 sky130_fd_sc_hd__mux2_1 _11868_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_05014_),
    .X(_05039_));
 sky130_fd_sc_hd__or2_1 _11870_ (.A(_04983_),
    .B(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__o211a_1 _11871_ (.A1(_05004_),
    .A2(_05038_),
    .B1(_05040_),
    .C1(_05010_),
    .X(_05041_));
 sky130_fd_sc_hd__mux2_1 _11872_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_05014_),
    .X(_05042_));
 sky130_fd_sc_hd__or2_1 _11873_ (.A(_04983_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_05014_),
    .X(_05044_));
 sky130_fd_sc_hd__o21a_1 _11875_ (.A1(_05003_),
    .A2(_05044_),
    .B1(_04999_),
    .X(_05045_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04988_),
    .X(_05046_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04988_),
    .X(_05047_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(_05046_),
    .A1(_05047_),
    .S(_05019_),
    .X(_05048_));
 sky130_fd_sc_hd__a221o_1 _11879_ (.A1(_05043_),
    .A2(_05045_),
    .B1(_05048_),
    .B2(_05010_),
    .C1(_04978_),
    .X(_05049_));
 sky130_fd_sc_hd__nor2_2 _11880_ (.A(_04971_),
    .B(_05026_),
    .Y(_05050_));
 sky130_fd_sc_hd__clkbuf_8 _11881_ (.A(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__o311a_1 _11882_ (.A1(_05030_),
    .A2(_05036_),
    .A3(_05041_),
    .B1(_05049_),
    .C1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__or3_1 _11883_ (.A(_04975_),
    .B(_05029_),
    .C(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__mux2_1 _11884_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_05037_),
    .X(_05054_));
 sky130_fd_sc_hd__or2_1 _11885_ (.A(_04984_),
    .B(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_05037_),
    .X(_05056_));
 sky130_fd_sc_hd__o21a_1 _11887_ (.A1(_05004_),
    .A2(_05056_),
    .B1(_05035_),
    .X(_05057_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_05037_),
    .X(_05058_));
 sky130_fd_sc_hd__mux2_1 _11889_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_05037_),
    .X(_05059_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(_05058_),
    .A1(_05059_),
    .S(_04984_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_8 _11891_ (.A(_05008_),
    .X(_05061_));
 sky130_fd_sc_hd__buf_4 _11892_ (.A(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__a221o_1 _11893_ (.A1(_05055_),
    .A2(_05057_),
    .B1(_05060_),
    .B2(_05062_),
    .C1(_05030_),
    .X(_05063_));
 sky130_fd_sc_hd__mux2_1 _11894_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_05037_),
    .X(_05064_));
 sky130_fd_sc_hd__mux2_1 _11895_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_05037_),
    .X(_05065_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(_05064_),
    .A1(_05065_),
    .S(_05004_),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _11897_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_05037_),
    .X(_05067_));
 sky130_fd_sc_hd__buf_4 _11898_ (.A(_04982_),
    .X(_05068_));
 sky130_fd_sc_hd__clkbuf_8 _11899_ (.A(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__buf_4 _11900_ (.A(_04986_),
    .X(_05070_));
 sky130_fd_sc_hd__buf_4 _11901_ (.A(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_8 _11902_ (.A(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__mux2_1 _11903_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__or2_1 _11904_ (.A(_05069_),
    .B(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__o211a_1 _11905_ (.A1(_05004_),
    .A2(_05067_),
    .B1(_05074_),
    .C1(_05035_),
    .X(_05075_));
 sky130_fd_sc_hd__a211o_1 _11906_ (.A1(_05062_),
    .A2(_05066_),
    .B1(_05075_),
    .C1(_04979_),
    .X(_05076_));
 sky130_fd_sc_hd__buf_4 _11907_ (.A(_04986_),
    .X(_05077_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _11909_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_05077_),
    .X(_05079_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(_05078_),
    .A1(_05079_),
    .S(_04992_),
    .X(_05080_));
 sky130_fd_sc_hd__mux2_1 _11911_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_05077_),
    .X(_05081_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_05077_),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(_05081_),
    .A1(_05082_),
    .S(_04992_),
    .X(_05083_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(_05080_),
    .A1(_05083_),
    .S(_05009_),
    .X(_05084_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_05077_),
    .X(_05085_));
 sky130_fd_sc_hd__mux2_1 _11916_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_05077_),
    .X(_05086_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(_05085_),
    .A1(_05086_),
    .S(_04992_),
    .X(_05087_));
 sky130_fd_sc_hd__mux2_1 _11918_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_05077_),
    .X(_05088_));
 sky130_fd_sc_hd__mux2_1 _11919_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04987_),
    .X(_05089_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(_05088_),
    .A1(_05089_),
    .S(_04982_),
    .X(_05090_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(_05087_),
    .A1(_05090_),
    .S(_05009_),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_1 _11922_ (.A0(_05084_),
    .A1(_05091_),
    .S(_05023_),
    .X(_05092_));
 sky130_fd_sc_hd__a21bo_1 _11923_ (.A1(_05051_),
    .A2(_05092_),
    .B1_N(_04975_),
    .X(_05093_));
 sky130_fd_sc_hd__a31o_1 _11924_ (.A1(_05028_),
    .A2(_05063_),
    .A3(_05076_),
    .B1(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__inv_2 _11925_ (.A(net3218),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(net3378),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__o211a_1 _11927_ (.A1(net3026),
    .A2(_04970_),
    .B1(_04985_),
    .C1(_04952_),
    .X(_05097_));
 sky130_fd_sc_hd__or3_1 _11928_ (.A(_05008_),
    .B(_05002_),
    .C(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__nand2_1 _11929_ (.A(net4303),
    .B(net4271),
    .Y(_05099_));
 sky130_fd_sc_hd__nand2_1 _11930_ (.A(net4254),
    .B(net4280),
    .Y(_05100_));
 sky130_fd_sc_hd__or4_1 _11931_ (.A(net4303),
    .B(net4271),
    .C(_05022_),
    .D(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__o41a_1 _11932_ (.A1(net4254),
    .A2(net4280),
    .A3(_04977_),
    .A4(_05099_),
    .B1(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__a21oi_1 _11933_ (.A1(_05098_),
    .A2(_05102_),
    .B1(net4239),
    .Y(_05103_));
 sky130_fd_sc_hd__or2_1 _11934_ (.A(net3014),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__inv_2 _11935_ (.A(net3014),
    .Y(_05105_));
 sky130_fd_sc_hd__a41o_1 _11936_ (.A1(net4239),
    .A2(_05000_),
    .A3(_04984_),
    .A4(_05037_),
    .B1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__nand2_1 _11937_ (.A(_05104_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__and3_1 _11938_ (.A(_04999_),
    .B(_04982_),
    .C(_05022_),
    .X(_05108_));
 sky130_fd_sc_hd__and3_1 _11939_ (.A(net7670),
    .B(net7677),
    .C(net7671),
    .X(_05109_));
 sky130_fd_sc_hd__nor3_1 _11940_ (.A(net4280),
    .B(net4303),
    .C(net4271),
    .Y(_05110_));
 sky130_fd_sc_hd__a31o_1 _11941_ (.A1(_05008_),
    .A2(_04992_),
    .A3(_04977_),
    .B1(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__o21ba_1 _11942_ (.A1(_05108_),
    .A2(_05109_),
    .B1_N(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__and3_1 _11943_ (.A(net3378),
    .B(net3218),
    .C(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__xnor2_1 _11944_ (.A(net3014),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__or2_1 _11945_ (.A(net3378),
    .B(_05095_),
    .X(_05115_));
 sky130_fd_sc_hd__mux2_1 _11946_ (.A0(_05107_),
    .A1(_05114_),
    .S(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__a31o_1 _11947_ (.A1(_05105_),
    .A2(net3378),
    .A3(_05095_),
    .B1(_04909_),
    .X(_05117_));
 sky130_fd_sc_hd__a21oi_1 _11948_ (.A1(_05096_),
    .A2(_05116_),
    .B1(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__a31o_1 _11949_ (.A1(_04909_),
    .A2(_05053_),
    .A3(_05094_),
    .B1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a21oi_4 _11950_ (.A1(_04161_),
    .A2(_04608_),
    .B1(net3992),
    .Y(_05120_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(net3144),
    .A1(net915),
    .S(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__inv_2 _11952_ (.A(net1673),
    .Y(_05122_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(net3016),
    .B(net1603),
    .Y(_05123_));
 sky130_fd_sc_hd__nand2_1 _11954_ (.A(_05122_),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__or2_1 _11955_ (.A(net1600),
    .B(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__or3_1 _11956_ (.A(net1793),
    .B(net2993),
    .C(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__and2_1 _11957_ (.A(net2955),
    .B(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__or2_2 _11958_ (.A(net3040),
    .B(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__xor2_1 _11959_ (.A(net2069),
    .B(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__a21oi_2 _11960_ (.A1(net2069),
    .A2(_05128_),
    .B1(net2869),
    .Y(_05130_));
 sky130_fd_sc_hd__and3_1 _11961_ (.A(net2869),
    .B(net2069),
    .C(_05128_),
    .X(_05131_));
 sky130_fd_sc_hd__nand2_1 _11962_ (.A(net3040),
    .B(_05127_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand2_1 _11963_ (.A(_05128_),
    .B(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__nor2_1 _11964_ (.A(net2955),
    .B(_05126_),
    .Y(_05134_));
 sky130_fd_sc_hd__nor2_1 _11965_ (.A(_05127_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_1 _11966_ (.A1(net2993),
    .A2(_05125_),
    .B1(net1793),
    .Y(_05136_));
 sky130_fd_sc_hd__nand2_1 _11967_ (.A(_05126_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__xnor2_1 _11968_ (.A(net2993),
    .B(_05125_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _11969_ (.A(net1600),
    .B(_05124_),
    .Y(_05139_));
 sky130_fd_sc_hd__nand2_1 _11970_ (.A(_05125_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__or2_1 _11971_ (.A(_04776_),
    .B(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__o21a_1 _11972_ (.A1(net3016),
    .A2(net3868),
    .B1(net2986),
    .X(_05142_));
 sky130_fd_sc_hd__and3_1 _11973_ (.A(net3016),
    .B(net1603),
    .C(\gpout0.hpos[0] ),
    .X(_05143_));
 sky130_fd_sc_hd__or2_1 _11974_ (.A(_05122_),
    .B(_05123_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_1 _11975_ (.A(_05124_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__o32a_1 _11976_ (.A1(_05123_),
    .A2(_05142_),
    .A3(_05143_),
    .B1(_05145_),
    .B2(net3987),
    .X(_05146_));
 sky130_fd_sc_hd__a221o_1 _11977_ (.A1(net1673),
    .A2(_04726_),
    .B1(_04776_),
    .B2(_05140_),
    .C1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__a22o_1 _11978_ (.A1(_05141_),
    .A2(_05147_),
    .B1(_05138_),
    .B2(_04604_),
    .X(_05148_));
 sky130_fd_sc_hd__o221a_1 _11979_ (.A1(_04604_),
    .A2(_05138_),
    .B1(_05137_),
    .B2(_04602_),
    .C1(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__a221o_1 _11980_ (.A1(_04602_),
    .A2(_05137_),
    .B1(_05135_),
    .B2(_04598_),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__o221a_1 _11981_ (.A1(_04598_),
    .A2(_05135_),
    .B1(_05133_),
    .B2(net4041),
    .C1(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__a221o_1 _11982_ (.A1(net4041),
    .A2(_05133_),
    .B1(_05129_),
    .B2(_04161_),
    .C1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__o221a_1 _11983_ (.A1(_04161_),
    .A2(_05129_),
    .B1(_05130_),
    .B2(_05131_),
    .C1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__a21o_1 _11984_ (.A1(net3040),
    .A2(net2955),
    .B1(net2069),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_1 _11985_ (.A(net2869),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_1 _11986_ (.A(net3992),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__nand3_1 _11987_ (.A(net2069),
    .B(net3040),
    .C(net2955),
    .Y(_05157_));
 sky130_fd_sc_hd__and2_1 _11988_ (.A(_05154_),
    .B(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__xnor2_1 _11989_ (.A(net3040),
    .B(net2955),
    .Y(_05159_));
 sky130_fd_sc_hd__inv_2 _11990_ (.A(net1793),
    .Y(_05160_));
 sky130_fd_sc_hd__inv_2 _11991_ (.A(net2993),
    .Y(_05161_));
 sky130_fd_sc_hd__inv_2 _11992_ (.A(net1600),
    .Y(_05162_));
 sky130_fd_sc_hd__inv_2 _11993_ (.A(net3016),
    .Y(_05163_));
 sky130_fd_sc_hd__a211oi_1 _11994_ (.A1(net3016),
    .A2(_04713_),
    .B1(_04719_),
    .C1(net1603),
    .Y(_05164_));
 sky130_fd_sc_hd__a221o_1 _11995_ (.A1(_05122_),
    .A2(net3987),
    .B1(net2986),
    .B2(_05163_),
    .C1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__o221a_1 _11996_ (.A1(_05122_),
    .A2(net3987),
    .B1(net3908),
    .B2(_05162_),
    .C1(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__a221o_1 _11997_ (.A1(_05161_),
    .A2(_04604_),
    .B1(_04776_),
    .B2(_05162_),
    .C1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__o221a_1 _11998_ (.A1(_05160_),
    .A2(net4009),
    .B1(_04604_),
    .B2(_05161_),
    .C1(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__a221o_1 _11999_ (.A1(net2955),
    .A2(_04598_),
    .B1(_04602_),
    .B2(_05160_),
    .C1(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__o221a_1 _12000_ (.A1(net2955),
    .A2(_04598_),
    .B1(_05159_),
    .B2(net4041),
    .C1(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__a221o_1 _12001_ (.A1(net4004),
    .A2(_05158_),
    .B1(_05159_),
    .B2(net4041),
    .C1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__o21ai_1 _12002_ (.A1(_04161_),
    .A2(_05158_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nor2_1 _12003_ (.A(net3992),
    .B(_05155_),
    .Y(_05173_));
 sky130_fd_sc_hd__a221o_1 _12004_ (.A1(net2869),
    .A2(_05154_),
    .B1(_05156_),
    .B2(_05172_),
    .C1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o21a_2 _12005_ (.A1(net3992),
    .A2(_05153_),
    .B1(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__or2b_1 _12006_ (.A(net694),
    .B_N(_05130_),
    .X(_05176_));
 sky130_fd_sc_hd__buf_4 _12007_ (.A(_04993_),
    .X(_05177_));
 sky130_fd_sc_hd__and4_1 _12008_ (.A(_05037_),
    .B(_05027_),
    .C(_04974_),
    .D(_05108_),
    .X(_05178_));
 sky130_fd_sc_hd__or3b_1 _12009_ (.A(_05177_),
    .B(_05120_),
    .C_N(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__o21ai_1 _12010_ (.A1(_05175_),
    .A2(_05176_),
    .B1(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__inv_2 _12011_ (.A(net3026),
    .Y(_05181_));
 sky130_fd_sc_hd__o211a_1 _12012_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04981_),
    .B1(_04987_),
    .C1(net1113),
    .X(_05182_));
 sky130_fd_sc_hd__a221o_1 _12013_ (.A1(net1524),
    .A2(_04998_),
    .B1(_04982_),
    .B2(\rbzero.floor_leak[1] ),
    .C1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__o221a_1 _12014_ (.A1(net1524),
    .A2(_04999_),
    .B1(_05022_),
    .B2(net1326),
    .C1(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__a221o_1 _12015_ (.A1(net1326),
    .A2(_05022_),
    .B1(_05027_),
    .B2(net1402),
    .C1(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__o221a_1 _12016_ (.A1(net1402),
    .A2(_05027_),
    .B1(_04975_),
    .B2(net4076),
    .C1(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__a221o_1 _12017_ (.A1(net4076),
    .A2(_04975_),
    .B1(_05180_),
    .B2(_05181_),
    .C1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_1 _12018_ (.A0(_05119_),
    .A1(_05121_),
    .S(net4077),
    .X(_05188_));
 sky130_fd_sc_hd__inv_2 _12019_ (.A(_04858_),
    .Y(_05189_));
 sky130_fd_sc_hd__o22a_1 _12020_ (.A1(net4065),
    .A2(net4094),
    .B1(_05188_),
    .B2(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__o22a_1 _12021_ (.A1(_04627_),
    .A2(_04817_),
    .B1(_04820_),
    .B2(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__nand2_1 _12022_ (.A(net4033),
    .B(_04831_),
    .Y(_05192_));
 sky130_fd_sc_hd__buf_1 _12023_ (.A(net4059),
    .X(_05193_));
 sky130_fd_sc_hd__buf_4 _12024_ (.A(net4033),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_2 _12025_ (.A(net4060),
    .B(net4034),
    .Y(_05195_));
 sky130_fd_sc_hd__or2_1 _12026_ (.A(net4059),
    .B(net4033),
    .X(_05196_));
 sky130_fd_sc_hd__or2b_1 _12027_ (.A(net3989),
    .B_N(_04803_),
    .X(_05197_));
 sky130_fd_sc_hd__a41o_1 _12028_ (.A1(_04806_),
    .A2(_05192_),
    .A3(_05195_),
    .A4(_05196_),
    .B1(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__o21a_1 _12029_ (.A1(net4041),
    .A2(net4004),
    .B1(net3992),
    .X(_05199_));
 sky130_fd_sc_hd__and3_1 _12030_ (.A(net4001),
    .B(net4972),
    .C(net4059),
    .X(_05200_));
 sky130_fd_sc_hd__a21o_4 _12031_ (.A1(net6041),
    .A2(_05200_),
    .B1(net6220),
    .X(_05201_));
 sky130_fd_sc_hd__a211oi_1 _12032_ (.A1(_04816_),
    .A2(_05198_),
    .B1(net4043),
    .C1(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__o21a_1 _12033_ (.A1(net83),
    .A2(_05191_),
    .B1(net4044),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_8 _12034_ (.A(net45),
    .X(_05204_));
 sky130_fd_sc_hd__mux2_4 _12035_ (.A0(\reg_rgb[6] ),
    .A1(_05203_),
    .S(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__clkbuf_1 _12036_ (.A(_05205_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _12037_ (.A0(net826),
    .A1(net7325),
    .S(_05120_),
    .X(_05206_));
 sky130_fd_sc_hd__buf_6 _12038_ (.A(net42),
    .X(_05207_));
 sky130_fd_sc_hd__a21oi_1 _12039_ (.A1(net3014),
    .A2(_05103_),
    .B1(_05115_),
    .Y(_05208_));
 sky130_fd_sc_hd__and2_1 _12040_ (.A(net3378),
    .B(_05095_),
    .X(_05209_));
 sky130_fd_sc_hd__a211o_1 _12041_ (.A1(_05105_),
    .A2(_05113_),
    .B1(_05208_),
    .C1(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__o21ai_1 _12042_ (.A1(net4254),
    .A2(_05051_),
    .B1(_05209_),
    .Y(_05211_));
 sky130_fd_sc_hd__a21o_1 _12043_ (.A1(net4254),
    .A2(_05051_),
    .B1(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__a31o_1 _12044_ (.A1(_05207_),
    .A2(_05210_),
    .A3(_05212_),
    .B1(net4077),
    .X(_05213_));
 sky130_fd_sc_hd__mux2_1 _12045_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_05072_),
    .X(_05214_));
 sky130_fd_sc_hd__mux2_1 _12046_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_05071_),
    .X(_05215_));
 sky130_fd_sc_hd__or2_1 _12047_ (.A(_05002_),
    .B(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__o211a_1 _12048_ (.A1(_05069_),
    .A2(_05214_),
    .B1(_05216_),
    .C1(_05061_),
    .X(_05217_));
 sky130_fd_sc_hd__clkbuf_8 _12049_ (.A(_05070_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_8 _12050_ (.A(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__mux2_1 _12051_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_05071_),
    .X(_05221_));
 sky130_fd_sc_hd__or2_1 _12053_ (.A(_05002_),
    .B(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__o211a_1 _12054_ (.A1(_05069_),
    .A2(_05220_),
    .B1(_05222_),
    .C1(_05034_),
    .X(_05223_));
 sky130_fd_sc_hd__mux2_1 _12055_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_05077_),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _12056_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_05077_),
    .X(_05225_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(_05224_),
    .A1(_05225_),
    .S(_05002_),
    .X(_05226_));
 sky130_fd_sc_hd__mux2_1 _12058_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_05071_),
    .X(_05227_));
 sky130_fd_sc_hd__or2_1 _12059_ (.A(_05002_),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__buf_4 _12060_ (.A(_04982_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_8 _12061_ (.A(_05070_),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__o21a_1 _12063_ (.A1(_05229_),
    .A2(_05231_),
    .B1(net80),
    .X(_05232_));
 sky130_fd_sc_hd__a221o_1 _12064_ (.A1(_05034_),
    .A2(_05226_),
    .B1(_05228_),
    .B2(_05232_),
    .C1(_05022_),
    .X(_05233_));
 sky130_fd_sc_hd__o31a_1 _12065_ (.A1(_04978_),
    .A2(_05217_),
    .A3(_05223_),
    .B1(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__buf_4 _12066_ (.A(_05002_),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_1 _12067_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_05072_),
    .X(_05236_));
 sky130_fd_sc_hd__mux2_1 _12068_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_05077_),
    .X(_05237_));
 sky130_fd_sc_hd__or2_1 _12069_ (.A(_05068_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__o211a_1 _12070_ (.A1(_05235_),
    .A2(_05236_),
    .B1(_05238_),
    .C1(_05034_),
    .X(_05239_));
 sky130_fd_sc_hd__mux2_1 _12071_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_05072_),
    .X(_05240_));
 sky130_fd_sc_hd__mux2_1 _12072_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_05071_),
    .X(_05241_));
 sky130_fd_sc_hd__or2_1 _12073_ (.A(_05068_),
    .B(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__o211a_1 _12074_ (.A1(_05235_),
    .A2(_05240_),
    .B1(_05242_),
    .C1(_05061_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_8 _12075_ (.A(_04999_),
    .X(_05244_));
 sky130_fd_sc_hd__mux2_1 _12076_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(_05071_),
    .X(_05245_));
 sky130_fd_sc_hd__mux2_1 _12077_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_05071_),
    .X(_05246_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(_05245_),
    .A1(_05246_),
    .S(_05002_),
    .X(_05247_));
 sky130_fd_sc_hd__buf_4 _12079_ (.A(_04992_),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_1 _12080_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_05230_),
    .X(_05249_));
 sky130_fd_sc_hd__mux2_1 _12081_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_05070_),
    .X(_05250_));
 sky130_fd_sc_hd__or2_1 _12082_ (.A(_04982_),
    .B(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__o211a_1 _12083_ (.A1(_05248_),
    .A2(_05249_),
    .B1(_05251_),
    .C1(_05009_),
    .X(_05252_));
 sky130_fd_sc_hd__a211o_1 _12084_ (.A1(_05244_),
    .A2(_05247_),
    .B1(_05252_),
    .C1(_05022_),
    .X(_05253_));
 sky130_fd_sc_hd__o31a_1 _12085_ (.A1(_04978_),
    .A2(_05239_),
    .A3(_05243_),
    .B1(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__mux2_1 _12086_ (.A0(_05234_),
    .A1(_05254_),
    .S(_05028_),
    .X(_05255_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_05014_),
    .X(_05256_));
 sky130_fd_sc_hd__mux2_1 _12088_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_05014_),
    .X(_05257_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(_05256_),
    .A1(_05257_),
    .S(_05003_),
    .X(_05258_));
 sky130_fd_sc_hd__mux2_1 _12090_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_05219_),
    .X(_05259_));
 sky130_fd_sc_hd__or2_1 _12091_ (.A(_05235_),
    .B(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__clkbuf_8 _12092_ (.A(_05229_),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_8 _12093_ (.A(_05070_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_8 _12094_ (.A(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__mux2_1 _12095_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__o21a_1 _12096_ (.A1(_05261_),
    .A2(_05264_),
    .B1(_05034_),
    .X(_05265_));
 sky130_fd_sc_hd__a221o_1 _12097_ (.A1(_05010_),
    .A2(_05258_),
    .B1(_05260_),
    .B2(_05265_),
    .C1(_05030_),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_1 _12098_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_05072_),
    .X(_05267_));
 sky130_fd_sc_hd__or2_1 _12099_ (.A(_05235_),
    .B(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _12100_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_05263_),
    .X(_05269_));
 sky130_fd_sc_hd__o21a_1 _12101_ (.A1(_05261_),
    .A2(_05269_),
    .B1(_05034_),
    .X(_05270_));
 sky130_fd_sc_hd__mux2_1 _12102_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_05072_),
    .X(_05271_));
 sky130_fd_sc_hd__mux2_1 _12103_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_05072_),
    .X(_05272_));
 sky130_fd_sc_hd__mux2_1 _12104_ (.A0(_05271_),
    .A1(_05272_),
    .S(_05235_),
    .X(_05273_));
 sky130_fd_sc_hd__a221o_1 _12105_ (.A1(_05268_),
    .A2(_05270_),
    .B1(_05273_),
    .B2(_05010_),
    .C1(_04978_),
    .X(_05274_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_05219_),
    .X(_05275_));
 sky130_fd_sc_hd__mux2_1 _12107_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_05071_),
    .X(_05276_));
 sky130_fd_sc_hd__or2_1 _12108_ (.A(_05002_),
    .B(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__o211a_1 _12109_ (.A1(_05069_),
    .A2(_05275_),
    .B1(_05277_),
    .C1(_05034_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_8 _12110_ (.A(_04993_),
    .X(_05279_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_05263_),
    .X(_05280_));
 sky130_fd_sc_hd__mux2_1 _12112_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_05218_),
    .X(_05281_));
 sky130_fd_sc_hd__or2_1 _12113_ (.A(_05068_),
    .B(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__o211a_1 _12114_ (.A1(_05279_),
    .A2(_05280_),
    .B1(_05282_),
    .C1(_05061_),
    .X(_05283_));
 sky130_fd_sc_hd__mux2_1 _12115_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_05230_),
    .X(_05284_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_05230_),
    .X(_05285_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(_05284_),
    .A1(_05285_),
    .S(_05068_),
    .X(_05286_));
 sky130_fd_sc_hd__mux2_1 _12118_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_05262_),
    .X(_05287_));
 sky130_fd_sc_hd__mux2_1 _12119_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_05070_),
    .X(_05288_));
 sky130_fd_sc_hd__or2_1 _12120_ (.A(_04992_),
    .B(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__o211a_1 _12121_ (.A1(_05019_),
    .A2(_05287_),
    .B1(_05289_),
    .C1(_05009_),
    .X(_05290_));
 sky130_fd_sc_hd__a211o_1 _12122_ (.A1(_05244_),
    .A2(_05286_),
    .B1(_05290_),
    .C1(_05023_),
    .X(_05291_));
 sky130_fd_sc_hd__o311a_1 _12123_ (.A1(_04978_),
    .A2(_05278_),
    .A3(_05283_),
    .B1(_05291_),
    .C1(_05050_),
    .X(_05292_));
 sky130_fd_sc_hd__a31o_1 _12124_ (.A1(_05028_),
    .A2(_05266_),
    .A3(_05274_),
    .B1(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__mux2_2 _12125_ (.A0(_05255_),
    .A1(_05293_),
    .S(_04975_),
    .X(_05294_));
 sky130_fd_sc_hd__nor2_1 _12126_ (.A(_05207_),
    .B(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__o2bb2a_1 _12127_ (.A1_N(net4077),
    .A2_N(_05206_),
    .B1(_05213_),
    .B2(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__inv_2 _12128_ (.A(_04892_),
    .Y(_05297_));
 sky130_fd_sc_hd__and4_1 _12129_ (.A(_04164_),
    .B(_04637_),
    .C(_04603_),
    .D(_04607_),
    .X(_05298_));
 sky130_fd_sc_hd__buf_4 _12130_ (.A(_04831_),
    .X(_05299_));
 sky130_fd_sc_hd__xnor2_1 _12131_ (.A(net4058),
    .B(_04602_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(_04806_),
    .B(_05192_),
    .Y(_05301_));
 sky130_fd_sc_hd__a32o_1 _12133_ (.A1(net4059),
    .A2(_04759_),
    .A3(_05301_),
    .B1(_04606_),
    .B2(net4014),
    .X(_05302_));
 sky130_fd_sc_hd__a32o_1 _12134_ (.A1(_05194_),
    .A2(_05299_),
    .A3(_05200_),
    .B1(_05300_),
    .B2(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__a22o_1 _12135_ (.A1(net4033),
    .A2(_04759_),
    .B1(_04606_),
    .B2(net4014),
    .X(_05304_));
 sky130_fd_sc_hd__a21o_1 _12136_ (.A1(_04831_),
    .A2(_04776_),
    .B1(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__o21bai_1 _12137_ (.A1(_05194_),
    .A2(_04759_),
    .B1_N(_05300_),
    .Y(_05306_));
 sky130_fd_sc_hd__o32a_1 _12138_ (.A1(_04599_),
    .A2(_05305_),
    .A3(_05306_),
    .B1(_04807_),
    .B2(net4001),
    .X(_05307_));
 sky130_fd_sc_hd__nor2_1 _12139_ (.A(net4972),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__or4b_2 _12140_ (.A(_05298_),
    .B(_05303_),
    .C(_05308_),
    .D_N(_04853_),
    .X(_05309_));
 sky130_fd_sc_hd__xnor2_1 _12141_ (.A(net4059),
    .B(_04776_),
    .Y(_05310_));
 sky130_fd_sc_hd__a22o_1 _12142_ (.A1(net4033),
    .A2(_04599_),
    .B1(_04759_),
    .B2(_04831_),
    .X(_05311_));
 sky130_fd_sc_hd__a221o_1 _12143_ (.A1(_04836_),
    .A2(net4010),
    .B1(_04605_),
    .B2(net4014),
    .C1(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__a2bb2o_1 _12144_ (.A1_N(_05194_),
    .A2_N(_04599_),
    .B1(_04602_),
    .B2(_04801_),
    .X(_05313_));
 sky130_fd_sc_hd__or3_1 _12145_ (.A(_05310_),
    .B(_05312_),
    .C(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__or4_1 _12146_ (.A(net4001),
    .B(_04831_),
    .C(_04164_),
    .D(_04600_),
    .X(_05315_));
 sky130_fd_sc_hd__or3b_1 _12147_ (.A(_04790_),
    .B(net4059),
    .C_N(_05194_),
    .X(_05316_));
 sky130_fd_sc_hd__or4_1 _12148_ (.A(_04836_),
    .B(_04603_),
    .C(_05315_),
    .D(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _12149_ (.A(_05314_),
    .B(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(_04880_),
    .B(_04904_),
    .Y(_05319_));
 sky130_fd_sc_hd__a31o_1 _12151_ (.A1(_05297_),
    .A2(_05309_),
    .A3(_05318_),
    .B1(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__a31oi_1 _12152_ (.A1(net4092),
    .A2(_04906_),
    .A3(_05320_),
    .B1(net4065),
    .Y(_05321_));
 sky130_fd_sc_hd__a21oi_1 _12153_ (.A1(_04858_),
    .A2(_05296_),
    .B1(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__o22a_1 _12154_ (.A1(_04626_),
    .A2(_04817_),
    .B1(_04820_),
    .B2(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__nand2_1 _12155_ (.A(net4037),
    .B(net4009),
    .Y(_05324_));
 sky130_fd_sc_hd__o22a_1 _12156_ (.A1(net4037),
    .A2(_04615_),
    .B1(_05324_),
    .B2(_04614_),
    .X(_05325_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(net4037),
    .A1(_05325_),
    .S(net3989),
    .X(_05326_));
 sky130_fd_sc_hd__o21ai_1 _12158_ (.A1(net4009),
    .A2(net3761),
    .B1(net4070),
    .Y(_05327_));
 sky130_fd_sc_hd__and2b_1 _12159_ (.A_N(net4052),
    .B(net4071),
    .X(_05328_));
 sky130_fd_sc_hd__or2_2 _12160_ (.A(_04814_),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__or3_1 _12161_ (.A(net4037),
    .B(net4009),
    .C(net3761),
    .X(_05330_));
 sky130_fd_sc_hd__nor2_1 _12162_ (.A(net3908),
    .B(_04811_),
    .Y(_05331_));
 sky130_fd_sc_hd__or2_1 _12163_ (.A(_04812_),
    .B(net3909),
    .X(_05332_));
 sky130_fd_sc_hd__nor2_1 _12164_ (.A(_04604_),
    .B(net3910),
    .Y(_05333_));
 sky130_fd_sc_hd__a21o_1 _12165_ (.A1(net4071),
    .A2(_05330_),
    .B1(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__or3_1 _12166_ (.A(_05326_),
    .B(_05329_),
    .C(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__inv_2 _12167_ (.A(_05329_),
    .Y(_05336_));
 sky130_fd_sc_hd__and2_1 _12168_ (.A(_05324_),
    .B(net4072),
    .X(_05337_));
 sky130_fd_sc_hd__a21oi_1 _12169_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_04814_),
    .Y(_05338_));
 sky130_fd_sc_hd__xnor2_1 _12170_ (.A(net4004),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__o21bai_1 _12171_ (.A1(_05335_),
    .A2(_05339_),
    .B1_N(_05326_),
    .Y(_05340_));
 sky130_fd_sc_hd__a21o_2 _12172_ (.A1(_05335_),
    .A2(_05339_),
    .B1(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__nor2_1 _12173_ (.A(_04612_),
    .B(_04615_),
    .Y(_05342_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(net4009),
    .A1(_05342_),
    .S(_04811_),
    .X(_05343_));
 sky130_fd_sc_hd__or3b_1 _12175_ (.A(_04815_),
    .B(net4005),
    .C_N(_05335_),
    .X(_05344_));
 sky130_fd_sc_hd__or3_1 _12176_ (.A(_04605_),
    .B(net3910),
    .C(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__or2_1 _12177_ (.A(_05343_),
    .B(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__nor2_1 _12178_ (.A(_05341_),
    .B(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__mux2_2 _12179_ (.A0(net4010),
    .A1(_04616_),
    .S(net3989),
    .X(_05348_));
 sky130_fd_sc_hd__nor3_1 _12180_ (.A(_04604_),
    .B(net3910),
    .C(_05344_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _12181_ (.A(_05348_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__nor2_1 _12182_ (.A(_05341_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__o21ba_1 _12183_ (.A1(net4038),
    .A2(net4072),
    .B1_N(_05337_),
    .X(_05352_));
 sky130_fd_sc_hd__xnor2_2 _12184_ (.A(_05329_),
    .B(net4073),
    .Y(_05353_));
 sky130_fd_sc_hd__nand2_1 _12185_ (.A(_04604_),
    .B(_04812_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_1 _12186_ (.A(net3761),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__or2b_1 _12187_ (.A(_05344_),
    .B_N(net3910),
    .X(_05356_));
 sky130_fd_sc_hd__nor2_1 _12188_ (.A(net3762),
    .B(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__inv_2 _12189_ (.A(_05339_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand2_2 _12190_ (.A(_05326_),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__nand2_1 _12191_ (.A(_05343_),
    .B(_05349_),
    .Y(_05360_));
 sky130_fd_sc_hd__and2b_1 _12192_ (.A_N(_05356_),
    .B(net3762),
    .X(_05361_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_05343_),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__and4b_1 _12194_ (.A_N(_05357_),
    .B(_05360_),
    .C(_05346_),
    .D(_05362_),
    .X(_05363_));
 sky130_fd_sc_hd__nor2_1 _12195_ (.A(_05359_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__nor2_1 _12196_ (.A(_05348_),
    .B(_05345_),
    .Y(_05365_));
 sky130_fd_sc_hd__a211o_1 _12197_ (.A1(_05343_),
    .A2(_05357_),
    .B1(_05364_),
    .C1(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_05348_),
    .B(_05361_),
    .Y(_05367_));
 sky130_fd_sc_hd__nor2_1 _12199_ (.A(_05341_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__and3b_1 _12200_ (.A_N(_05341_),
    .B(_05348_),
    .C(_05357_),
    .X(_05369_));
 sky130_fd_sc_hd__a211o_1 _12201_ (.A1(_05353_),
    .A2(_05366_),
    .B1(_05368_),
    .C1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__or3_2 _12202_ (.A(_05347_),
    .B(_05351_),
    .C(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__nor2_2 _12203_ (.A(_05341_),
    .B(_05362_),
    .Y(_05372_));
 sky130_fd_sc_hd__and2b_2 _12204_ (.A_N(_05341_),
    .B(_05365_),
    .X(_05373_));
 sky130_fd_sc_hd__and3b_2 _12205_ (.A_N(_05341_),
    .B(_05343_),
    .C(_05357_),
    .X(_05374_));
 sky130_fd_sc_hd__a22o_1 _12206_ (.A1(\rbzero.debug_overlay.facingY[-3] ),
    .A2(_05373_),
    .B1(_05374_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .X(_05375_));
 sky130_fd_sc_hd__or2_2 _12207_ (.A(_05353_),
    .B(_05359_),
    .X(_05376_));
 sky130_fd_sc_hd__nor2_2 _12208_ (.A(_05362_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__and3b_2 _12209_ (.A_N(_05376_),
    .B(_05348_),
    .C(_05357_),
    .X(_05378_));
 sky130_fd_sc_hd__nor2_2 _12210_ (.A(_05346_),
    .B(_05376_),
    .Y(_05379_));
 sky130_fd_sc_hd__a22o_1 _12211_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_05378_),
    .B1(_05379_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .X(_05380_));
 sky130_fd_sc_hd__nor2_2 _12212_ (.A(_05341_),
    .B(_05360_),
    .Y(_05381_));
 sky130_fd_sc_hd__nor2_2 _12213_ (.A(_05360_),
    .B(_05376_),
    .Y(_05382_));
 sky130_fd_sc_hd__nor2_2 _12214_ (.A(_05367_),
    .B(_05359_),
    .Y(_05383_));
 sky130_fd_sc_hd__nor2_2 _12215_ (.A(_05350_),
    .B(_05359_),
    .Y(_05384_));
 sky130_fd_sc_hd__a22o_1 _12216_ (.A1(\rbzero.debug_overlay.facingY[-4] ),
    .A2(_05383_),
    .B1(_05384_),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .X(_05385_));
 sky130_fd_sc_hd__a221o_1 _12217_ (.A1(\rbzero.debug_overlay.facingY[-1] ),
    .A2(_05381_),
    .B1(_05382_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .C1(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__a211o_1 _12218_ (.A1(\rbzero.debug_overlay.facingY[-8] ),
    .A2(_05377_),
    .B1(_05380_),
    .C1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__a211o_1 _12219_ (.A1(net3857),
    .A2(_05372_),
    .B1(_05375_),
    .C1(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__a21oi_1 _12220_ (.A1(net3876),
    .A2(_05371_),
    .B1(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__or3_1 _12221_ (.A(_04881_),
    .B(_04806_),
    .C(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__buf_2 _12222_ (.A(net4625),
    .X(_05391_));
 sky130_fd_sc_hd__a22o_1 _12223_ (.A1(net3699),
    .A2(_05374_),
    .B1(_05372_),
    .B2(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_4 _12224_ (.A(net4620),
    .X(_05393_));
 sky130_fd_sc_hd__a22o_1 _12225_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_05382_),
    .B1(_05378_),
    .B2(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_05394_));
 sky130_fd_sc_hd__a221o_1 _12226_ (.A1(_05393_),
    .A2(_05377_),
    .B1(_05379_),
    .B2(\rbzero.debug_overlay.vplaneY[-7] ),
    .C1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_4 _12227_ (.A(net4549),
    .X(_05396_));
 sky130_fd_sc_hd__a221o_1 _12228_ (.A1(net3807),
    .A2(_05383_),
    .B1(_05384_),
    .B2(_05396_),
    .C1(_04889_),
    .X(_05397_));
 sky130_fd_sc_hd__a211o_1 _12229_ (.A1(\rbzero.debug_overlay.vplaneY[-3] ),
    .A2(_05373_),
    .B1(_05395_),
    .C1(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__a211o_1 _12230_ (.A1(_05391_),
    .A2(_05381_),
    .B1(_05392_),
    .C1(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__a21oi_1 _12231_ (.A1(net4708),
    .A2(_05371_),
    .B1(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__clkbuf_4 _12232_ (.A(net4772),
    .X(_05401_));
 sky130_fd_sc_hd__a22o_1 _12233_ (.A1(net3241),
    .A2(_05374_),
    .B1(_05372_),
    .B2(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_4 _12234_ (.A(net4656),
    .X(_05403_));
 sky130_fd_sc_hd__a22o_1 _12235_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_05382_),
    .B1(_05378_),
    .B2(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_05404_));
 sky130_fd_sc_hd__a221o_1 _12236_ (.A1(_05403_),
    .A2(_05377_),
    .B1(_05379_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_1 _12237_ (.A(net3837),
    .X(_05406_));
 sky130_fd_sc_hd__a221o_1 _12238_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(_05383_),
    .B1(_05384_),
    .B2(net3838),
    .C1(_04831_),
    .X(_05407_));
 sky130_fd_sc_hd__a211o_1 _12239_ (.A1(\rbzero.debug_overlay.vplaneX[-3] ),
    .A2(_05373_),
    .B1(_05405_),
    .C1(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__a211o_1 _12240_ (.A1(_05401_),
    .A2(_05381_),
    .B1(_05402_),
    .C1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__a21oi_1 _12241_ (.A1(net4666),
    .A2(_05371_),
    .B1(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__or3_2 _12242_ (.A(_05195_),
    .B(_05400_),
    .C(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__a22o_1 _12243_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(_05374_),
    .B1(_05372_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .X(_05412_));
 sky130_fd_sc_hd__a22o_1 _12244_ (.A1(\rbzero.debug_overlay.facingX[-8] ),
    .A2(_05377_),
    .B1(_05378_),
    .B2(\rbzero.debug_overlay.facingX[-6] ),
    .X(_05413_));
 sky130_fd_sc_hd__a22o_1 _12245_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_05383_),
    .B1(_05384_),
    .B2(\rbzero.debug_overlay.facingX[-5] ),
    .X(_05414_));
 sky130_fd_sc_hd__a221o_1 _12246_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_05373_),
    .B1(_05379_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .C1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__a211o_1 _12247_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(_05382_),
    .B1(_05413_),
    .C1(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__a211o_1 _12248_ (.A1(net3786),
    .A2(_05381_),
    .B1(_05412_),
    .C1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__a21oi_2 _12249_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_05371_),
    .B1(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a211o_1 _12250_ (.A1(_05194_),
    .A2(_05418_),
    .B1(net4014),
    .C1(_05193_),
    .X(_05419_));
 sky130_fd_sc_hd__a22o_1 _12251_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_05374_),
    .B1(_05372_),
    .B2(net3917),
    .X(_05420_));
 sky130_fd_sc_hd__a22o_1 _12252_ (.A1(net3024),
    .A2(_05377_),
    .B1(_05382_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .X(_05421_));
 sky130_fd_sc_hd__a22o_1 _12253_ (.A1(net2942),
    .A2(_05378_),
    .B1(_05379_),
    .B2(net2940),
    .X(_05422_));
 sky130_fd_sc_hd__a22o_1 _12254_ (.A1(net3880),
    .A2(_05347_),
    .B1(_05351_),
    .B2(net3893),
    .X(_05423_));
 sky130_fd_sc_hd__a221o_1 _12255_ (.A1(net4063),
    .A2(_05373_),
    .B1(_05368_),
    .B2(net3279),
    .C1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__and2_1 _12256_ (.A(_05365_),
    .B(_05353_),
    .X(_05425_));
 sky130_fd_sc_hd__a22o_1 _12257_ (.A1(net3003),
    .A2(_05383_),
    .B1(_05425_),
    .B2(net3952),
    .X(_05426_));
 sky130_fd_sc_hd__a22o_1 _12258_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_05369_),
    .B1(_05384_),
    .B2(\rbzero.debug_overlay.playerY[-5] ),
    .X(_05427_));
 sky130_fd_sc_hd__or4_1 _12259_ (.A(_04889_),
    .B(_05196_),
    .C(_05426_),
    .D(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__or4_1 _12260_ (.A(_05421_),
    .B(_05422_),
    .C(_05424_),
    .D(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__a211oi_1 _12261_ (.A1(net4288),
    .A2(_05381_),
    .B1(_05420_),
    .C1(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__a31o_1 _12262_ (.A1(_05390_),
    .A2(_05411_),
    .A3(_05419_),
    .B1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__a22o_1 _12263_ (.A1(net3028),
    .A2(_05374_),
    .B1(_05372_),
    .B2(net3821),
    .X(_05432_));
 sky130_fd_sc_hd__a22o_1 _12264_ (.A1(net4306),
    .A2(_05377_),
    .B1(_05378_),
    .B2(net4338),
    .X(_05433_));
 sky130_fd_sc_hd__a22o_1 _12265_ (.A1(net7369),
    .A2(_05382_),
    .B1(_05379_),
    .B2(net2933),
    .X(_05434_));
 sky130_fd_sc_hd__a22o_1 _12266_ (.A1(net3008),
    .A2(_05373_),
    .B1(_05381_),
    .B2(net4218),
    .X(_05435_));
 sky130_fd_sc_hd__a221o_1 _12267_ (.A1(net3853),
    .A2(_05368_),
    .B1(_05347_),
    .B2(net3995),
    .C1(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__a221o_1 _12268_ (.A1(net7427),
    .A2(_05383_),
    .B1(_05425_),
    .B2(\rbzero.debug_overlay.playerX[5] ),
    .C1(_04807_),
    .X(_05437_));
 sky130_fd_sc_hd__a221o_1 _12269_ (.A1(net3921),
    .A2(_05351_),
    .B1(_05384_),
    .B2(net2935),
    .C1(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__or4_1 _12270_ (.A(_05433_),
    .B(_05434_),
    .C(_05436_),
    .D(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__a211oi_1 _12271_ (.A1(net4090),
    .A2(_05369_),
    .B1(_05432_),
    .C1(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__a211o_1 _12272_ (.A1(_04807_),
    .A2(_05431_),
    .B1(_05440_),
    .C1(_05197_),
    .X(_05441_));
 sky130_fd_sc_hd__a2111oi_1 _12273_ (.A1(_04614_),
    .A2(_04790_),
    .B1(_04161_),
    .C1(_04601_),
    .D1(_04608_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand4_1 _12274_ (.A(_05342_),
    .B(_05197_),
    .C(_05333_),
    .D(net85),
    .Y(_05443_));
 sky130_fd_sc_hd__a311oi_1 _12275_ (.A1(_04816_),
    .A2(_05441_),
    .A3(_05443_),
    .B1(net4043),
    .C1(_05201_),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_1 _12276_ (.A1(net83),
    .A2(_05323_),
    .B1(net4006),
    .Y(_05445_));
 sky130_fd_sc_hd__clkinv_4 _12277_ (.A(net4007),
    .Y(_05446_));
 sky130_fd_sc_hd__mux2_4 _12278_ (.A0(\reg_rgb[7] ),
    .A1(_05446_),
    .S(_05204_),
    .X(_05447_));
 sky130_fd_sc_hd__clkbuf_1 _12279_ (.A(_05447_),
    .X(net71));
 sky130_fd_sc_hd__a21o_1 _12280_ (.A1(net4532),
    .A2(_05111_),
    .B1(_05095_),
    .X(_05448_));
 sky130_fd_sc_hd__o2111a_1 _12281_ (.A1(net4239),
    .A2(_05102_),
    .B1(_05097_),
    .C1(_05004_),
    .D1(_05010_),
    .X(_05449_));
 sky130_fd_sc_hd__o21ai_1 _12282_ (.A1(_05106_),
    .A2(_05449_),
    .B1(_05104_),
    .Y(_05450_));
 sky130_fd_sc_hd__o2bb2a_1 _12283_ (.A1_N(net3378),
    .A2_N(_05448_),
    .B1(_05450_),
    .B2(_05115_),
    .X(_05451_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_05219_),
    .X(_05452_));
 sky130_fd_sc_hd__mux2_1 _12285_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_05071_),
    .X(_05453_));
 sky130_fd_sc_hd__or2_1 _12286_ (.A(_05248_),
    .B(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__o211a_1 _12287_ (.A1(_05069_),
    .A2(_05452_),
    .B1(_05454_),
    .C1(_05034_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_8 _12288_ (.A(_04987_),
    .X(_05456_));
 sky130_fd_sc_hd__buf_4 _12289_ (.A(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__mux2_1 _12291_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_05230_),
    .X(_05459_));
 sky130_fd_sc_hd__or2_1 _12292_ (.A(_05229_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__buf_4 _12293_ (.A(_05009_),
    .X(_05461_));
 sky130_fd_sc_hd__o211a_1 _12294_ (.A1(_05279_),
    .A2(_05458_),
    .B1(_05460_),
    .C1(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_05262_),
    .X(_05463_));
 sky130_fd_sc_hd__or2_1 _12296_ (.A(_05229_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_05456_),
    .X(_05465_));
 sky130_fd_sc_hd__o21a_1 _12298_ (.A1(_04993_),
    .A2(_05465_),
    .B1(_04999_),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_05218_),
    .X(_05467_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_05218_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(_05467_),
    .A1(_05468_),
    .S(_05068_),
    .X(_05469_));
 sky130_fd_sc_hd__a221o_1 _12302_ (.A1(_05464_),
    .A2(_05466_),
    .B1(_05469_),
    .B2(_05061_),
    .C1(net81),
    .X(_05470_));
 sky130_fd_sc_hd__o311a_1 _12303_ (.A1(_05030_),
    .A2(_05455_),
    .A3(_05462_),
    .B1(_05470_),
    .C1(_05051_),
    .X(_05471_));
 sky130_fd_sc_hd__mux2_1 _12304_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_05263_),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_05230_),
    .X(_05473_));
 sky130_fd_sc_hd__or2_1 _12306_ (.A(_05248_),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__o211a_1 _12307_ (.A1(_05261_),
    .A2(_05472_),
    .B1(_05474_),
    .C1(_05244_),
    .X(_05475_));
 sky130_fd_sc_hd__buf_4 _12308_ (.A(_05456_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _12310_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_05262_),
    .X(_05478_));
 sky130_fd_sc_hd__or2_1 _12311_ (.A(_05229_),
    .B(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__o211a_1 _12312_ (.A1(_05279_),
    .A2(_05477_),
    .B1(_05479_),
    .C1(_05461_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_05456_),
    .X(_05481_));
 sky130_fd_sc_hd__or2_1 _12314_ (.A(_05019_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__buf_4 _12315_ (.A(_04987_),
    .X(_05483_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__o21a_1 _12317_ (.A1(_04993_),
    .A2(_05484_),
    .B1(_04999_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_05262_),
    .X(_05486_));
 sky130_fd_sc_hd__mux2_1 _12319_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_05262_),
    .X(_05487_));
 sky130_fd_sc_hd__mux2_1 _12320_ (.A0(_05486_),
    .A1(_05487_),
    .S(_05068_),
    .X(_05488_));
 sky130_fd_sc_hd__a221o_1 _12321_ (.A1(_05482_),
    .A2(_05485_),
    .B1(_05488_),
    .B2(_05061_),
    .C1(_05023_),
    .X(_05489_));
 sky130_fd_sc_hd__o311a_1 _12322_ (.A1(_04978_),
    .A2(_05475_),
    .A3(_05480_),
    .B1(_05489_),
    .C1(_05027_),
    .X(_05490_));
 sky130_fd_sc_hd__nor2_1 _12323_ (.A(_05471_),
    .B(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_05070_),
    .X(_05492_));
 sky130_fd_sc_hd__buf_4 _12325_ (.A(_04986_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__mux2_1 _12327_ (.A0(_05492_),
    .A1(_05494_),
    .S(_04992_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_05070_),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_1 _12329_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_05493_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(_05496_),
    .A1(_05497_),
    .S(_04991_),
    .X(_05498_));
 sky130_fd_sc_hd__mux2_1 _12331_ (.A0(_05495_),
    .A1(_05498_),
    .S(net80),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_05070_),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _12333_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_05493_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _12334_ (.A0(_05500_),
    .A1(_05501_),
    .S(_04992_),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _12335_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_05493_),
    .X(_05503_));
 sky130_fd_sc_hd__mux2_1 _12336_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_05493_),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _12337_ (.A0(_05503_),
    .A1(_05504_),
    .S(_04981_),
    .X(_05505_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(_05502_),
    .A1(_05505_),
    .S(net80),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _12339_ (.A0(_05499_),
    .A1(_05506_),
    .S(_05022_),
    .X(_05507_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_05070_),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _12341_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_05493_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(_05508_),
    .A1(_05509_),
    .S(_04991_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _12343_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_05493_),
    .X(_05511_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04986_),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(_05511_),
    .A1(_05512_),
    .S(_04981_),
    .X(_05513_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(_05510_),
    .A1(_05513_),
    .S(net80),
    .X(_05514_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_05493_),
    .X(_05515_));
 sky130_fd_sc_hd__mux2_1 _12348_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_05493_),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(_05515_),
    .A1(_05516_),
    .S(_04991_),
    .X(_05517_));
 sky130_fd_sc_hd__mux2_1 _12350_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_05493_),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04986_),
    .X(_05519_));
 sky130_fd_sc_hd__mux2_1 _12352_ (.A0(_05518_),
    .A1(_05519_),
    .S(_04991_),
    .X(_05520_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(_05517_),
    .A1(_05520_),
    .S(net80),
    .X(_05521_));
 sky130_fd_sc_hd__mux2_1 _12354_ (.A0(_05514_),
    .A1(_05521_),
    .S(_05022_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(_05507_),
    .A1(_05522_),
    .S(_05027_),
    .X(_05523_));
 sky130_fd_sc_hd__nand2_1 _12356_ (.A(_04975_),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_1 _12357_ (.A1(_04975_),
    .A2(_05491_),
    .B1(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__a2bb2o_1 _12358_ (.A1_N(_05117_),
    .A2_N(_05451_),
    .B1(_05525_),
    .B2(_04909_),
    .X(_05526_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(net7322),
    .A1(net1027),
    .S(_05120_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_2 _12360_ (.A0(_05526_),
    .A1(_05527_),
    .S(net4077),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(_04842_),
    .A1(_05528_),
    .S(_04858_),
    .X(_05529_));
 sky130_fd_sc_hd__o22a_1 _12362_ (.A1(net6168),
    .A2(_04817_),
    .B1(_04820_),
    .B2(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__o21a_1 _12363_ (.A1(_04816_),
    .A2(_05530_),
    .B1(net4044),
    .X(_05531_));
 sky130_fd_sc_hd__mux2_2 _12364_ (.A0(\reg_rgb[14] ),
    .A1(_05531_),
    .S(_05204_),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_1 _12365_ (.A(_05532_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _12366_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_05219_),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _12367_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_05218_),
    .X(_05534_));
 sky130_fd_sc_hd__or2_1 _12368_ (.A(_05248_),
    .B(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__o211a_1 _12369_ (.A1(_05069_),
    .A2(_05533_),
    .B1(_05535_),
    .C1(_05061_),
    .X(_05536_));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_05457_),
    .X(_05537_));
 sky130_fd_sc_hd__mux2_1 _12371_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_05230_),
    .X(_05538_));
 sky130_fd_sc_hd__or2_1 _12372_ (.A(_05248_),
    .B(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__o211a_1 _12373_ (.A1(_05261_),
    .A2(_05537_),
    .B1(_05539_),
    .C1(_05244_),
    .X(_05540_));
 sky130_fd_sc_hd__buf_4 _12374_ (.A(_05483_),
    .X(_05541_));
 sky130_fd_sc_hd__mux2_1 _12375_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_05483_),
    .X(_05543_));
 sky130_fd_sc_hd__or2_1 _12377_ (.A(_04993_),
    .B(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__o211a_1 _12378_ (.A1(_05261_),
    .A2(_05542_),
    .B1(_05544_),
    .C1(_05000_),
    .X(_05545_));
 sky130_fd_sc_hd__mux2_1 _12379_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_05483_),
    .X(_05546_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\rbzero.tex_g1[63] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_05483_),
    .X(_05547_));
 sky130_fd_sc_hd__mux2_1 _12381_ (.A0(_05546_),
    .A1(_05547_),
    .S(_05248_),
    .X(_05548_));
 sky130_fd_sc_hd__a21o_1 _12382_ (.A1(_05461_),
    .A2(_05548_),
    .B1(_05023_),
    .X(_05549_));
 sky130_fd_sc_hd__o32a_1 _12383_ (.A1(_04978_),
    .A2(_05536_),
    .A3(_05540_),
    .B1(_05545_),
    .B2(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_05457_),
    .X(_05551_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_05262_),
    .X(_05552_));
 sky130_fd_sc_hd__or2_1 _12386_ (.A(_05229_),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__o211a_1 _12387_ (.A1(_05279_),
    .A2(_05551_),
    .B1(_05553_),
    .C1(_05244_),
    .X(_05554_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_05476_),
    .X(_05555_));
 sky130_fd_sc_hd__mux2_1 _12389_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_05456_),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _12390_ (.A(_05019_),
    .B(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__o211a_1 _12391_ (.A1(_05177_),
    .A2(_05555_),
    .B1(_05557_),
    .C1(_05461_),
    .X(_05558_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_05456_),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_05456_),
    .X(_05560_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(_05559_),
    .A1(_05560_),
    .S(_05248_),
    .X(_05561_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_05483_),
    .X(_05562_));
 sky130_fd_sc_hd__mux2_1 _12396_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_04987_),
    .X(_05563_));
 sky130_fd_sc_hd__or2_1 _12397_ (.A(_04982_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__o211a_1 _12398_ (.A1(_04993_),
    .A2(_05562_),
    .B1(_05564_),
    .C1(_05009_),
    .X(_05565_));
 sky130_fd_sc_hd__a211o_1 _12399_ (.A1(_05000_),
    .A2(_05561_),
    .B1(_05565_),
    .C1(_05023_),
    .X(_05566_));
 sky130_fd_sc_hd__o31a_1 _12400_ (.A1(_04979_),
    .A2(_05554_),
    .A3(_05558_),
    .B1(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(_05550_),
    .A1(_05567_),
    .S(_05028_),
    .X(_05568_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_05263_),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_05263_),
    .X(_05570_));
 sky130_fd_sc_hd__mux2_1 _12404_ (.A0(_05569_),
    .A1(_05570_),
    .S(_05235_),
    .X(_05571_));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_05476_),
    .X(_05572_));
 sky130_fd_sc_hd__or2_1 _12406_ (.A(_05177_),
    .B(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_05541_),
    .X(_05574_));
 sky130_fd_sc_hd__o21a_1 _12408_ (.A1(_04984_),
    .A2(_05574_),
    .B1(_05000_),
    .X(_05575_));
 sky130_fd_sc_hd__a221o_1 _12409_ (.A1(_05062_),
    .A2(_05571_),
    .B1(_05573_),
    .B2(_05575_),
    .C1(_05030_),
    .X(_05576_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(_05476_),
    .X(_05577_));
 sky130_fd_sc_hd__or2_1 _12411_ (.A(_05279_),
    .B(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_05476_),
    .X(_05579_));
 sky130_fd_sc_hd__o21a_1 _12413_ (.A1(_05261_),
    .A2(_05579_),
    .B1(_05244_),
    .X(_05580_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_05457_),
    .X(_05581_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_05457_),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(_05581_),
    .A1(_05582_),
    .S(_05235_),
    .X(_05583_));
 sky130_fd_sc_hd__a221o_1 _12417_ (.A1(_05578_),
    .A2(_05580_),
    .B1(_05583_),
    .B2(_05062_),
    .C1(_04979_),
    .X(_05584_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_05476_),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_05456_),
    .X(_05586_));
 sky130_fd_sc_hd__or2_1 _12420_ (.A(_05019_),
    .B(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__o211a_1 _12421_ (.A1(_05177_),
    .A2(_05585_),
    .B1(_05587_),
    .C1(_05244_),
    .X(_05588_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_05541_),
    .X(_05589_));
 sky130_fd_sc_hd__mux2_1 _12423_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_05483_),
    .X(_05590_));
 sky130_fd_sc_hd__or2_1 _12424_ (.A(_05019_),
    .B(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__o211a_1 _12425_ (.A1(_05177_),
    .A2(_05589_),
    .B1(_05591_),
    .C1(_05461_),
    .X(_05592_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_05483_),
    .X(_05593_));
 sky130_fd_sc_hd__mux2_1 _12427_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_05483_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(_05593_),
    .A1(_05594_),
    .S(_04993_),
    .X(_05595_));
 sky130_fd_sc_hd__mux2_1 _12429_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04994_),
    .X(_05596_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04987_),
    .X(_05597_));
 sky130_fd_sc_hd__or2_1 _12431_ (.A(_04982_),
    .B(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o211a_1 _12432_ (.A1(_05003_),
    .A2(_05596_),
    .B1(_05598_),
    .C1(_05009_),
    .X(_05599_));
 sky130_fd_sc_hd__a211o_1 _12433_ (.A1(_05000_),
    .A2(_05595_),
    .B1(_05599_),
    .C1(_04978_),
    .X(_05600_));
 sky130_fd_sc_hd__o311a_1 _12434_ (.A1(_05030_),
    .A2(_05588_),
    .A3(_05592_),
    .B1(_05051_),
    .C1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__a31o_1 _12435_ (.A1(_05028_),
    .A2(_05576_),
    .A3(_05584_),
    .B1(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__mux2_2 _12436_ (.A0(_05568_),
    .A1(_05602_),
    .S(_04975_),
    .X(_05603_));
 sky130_fd_sc_hd__or3b_1 _12437_ (.A(_05105_),
    .B(_05115_),
    .C_N(_05103_),
    .X(_05604_));
 sky130_fd_sc_hd__a21oi_1 _12438_ (.A1(net4303),
    .A2(_05062_),
    .B1(_05096_),
    .Y(_05605_));
 sky130_fd_sc_hd__o21ai_1 _12439_ (.A1(net4303),
    .A2(_05062_),
    .B1(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__a31o_1 _12440_ (.A1(net42),
    .A2(_05604_),
    .A3(_05606_),
    .B1(net4077),
    .X(_05607_));
 sky130_fd_sc_hd__o21ba_1 _12441_ (.A1(_05207_),
    .A2(_05603_),
    .B1_N(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_1 _12442_ (.A0(net788),
    .A1(net7327),
    .S(_05120_),
    .X(_05609_));
 sky130_fd_sc_hd__and2_1 _12443_ (.A(net4077),
    .B(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__nor2_1 _12444_ (.A(_04892_),
    .B(_05319_),
    .Y(_05611_));
 sky130_fd_sc_hd__and4bb_1 _12445_ (.A_N(net4093),
    .B_N(_05318_),
    .C(_05611_),
    .D(_05309_),
    .X(_05612_));
 sky130_fd_sc_hd__o32a_1 _12446_ (.A1(_05189_),
    .A2(_05608_),
    .A3(_05610_),
    .B1(net4065),
    .B2(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__o22a_1 _12447_ (.A1(net4909),
    .A2(_04817_),
    .B1(_04820_),
    .B2(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__o21a_1 _12448_ (.A1(net83),
    .A2(_05614_),
    .B1(net4006),
    .X(_05615_));
 sky130_fd_sc_hd__mux2_2 _12449_ (.A0(\reg_rgb[15] ),
    .A1(_05615_),
    .S(_05204_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_05616_),
    .X(net67));
 sky130_fd_sc_hd__a31o_1 _12451_ (.A1(_05062_),
    .A2(_05004_),
    .A3(_05097_),
    .B1(_05104_),
    .X(_05617_));
 sky130_fd_sc_hd__or3b_1 _12452_ (.A(_05111_),
    .B(net3014),
    .C_N(net3378),
    .X(_05618_));
 sky130_fd_sc_hd__inv_2 _12453_ (.A(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__a221oi_1 _12454_ (.A1(net3378),
    .A2(_05448_),
    .B1(_05617_),
    .B2(_05208_),
    .C1(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_05072_),
    .X(_05621_));
 sky130_fd_sc_hd__mux2_1 _12456_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_05014_),
    .X(_05622_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(_05621_),
    .A1(_05622_),
    .S(_05003_),
    .X(_05623_));
 sky130_fd_sc_hd__mux2_1 _12458_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_05263_),
    .X(_05624_));
 sky130_fd_sc_hd__or2_1 _12459_ (.A(_05235_),
    .B(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__mux2_1 _12460_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_05457_),
    .X(_05626_));
 sky130_fd_sc_hd__o21a_1 _12461_ (.A1(_05261_),
    .A2(_05626_),
    .B1(_05244_),
    .X(_05627_));
 sky130_fd_sc_hd__a221o_1 _12462_ (.A1(_05062_),
    .A2(_05623_),
    .B1(_05625_),
    .B2(_05627_),
    .C1(_04979_),
    .X(_05628_));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_05219_),
    .X(_05629_));
 sky130_fd_sc_hd__or2_1 _12464_ (.A(_05069_),
    .B(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_05457_),
    .X(_05631_));
 sky130_fd_sc_hd__o21a_1 _12466_ (.A1(_05279_),
    .A2(_05631_),
    .B1(_05034_),
    .X(_05632_));
 sky130_fd_sc_hd__mux2_1 _12467_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_05072_),
    .X(_05633_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_05072_),
    .X(_05634_));
 sky130_fd_sc_hd__mux2_1 _12469_ (.A0(_05633_),
    .A1(_05634_),
    .S(_05069_),
    .X(_05635_));
 sky130_fd_sc_hd__a221o_1 _12470_ (.A1(_05630_),
    .A2(_05632_),
    .B1(_05635_),
    .B2(_05010_),
    .C1(_05030_),
    .X(_05636_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_05219_),
    .X(_05637_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_05218_),
    .X(_05638_));
 sky130_fd_sc_hd__or2_1 _12473_ (.A(_05248_),
    .B(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__o211a_1 _12474_ (.A1(_05069_),
    .A2(_05637_),
    .B1(_05639_),
    .C1(_05244_),
    .X(_05640_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_05457_),
    .X(_05641_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_05230_),
    .X(_05642_));
 sky130_fd_sc_hd__or2_1 _12477_ (.A(_05248_),
    .B(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__o211a_1 _12478_ (.A1(_05261_),
    .A2(_05641_),
    .B1(_05643_),
    .C1(_05461_),
    .X(_05644_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_05262_),
    .X(_05645_));
 sky130_fd_sc_hd__or2_1 _12480_ (.A(_05248_),
    .B(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__mux2_1 _12481_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_05456_),
    .X(_05647_));
 sky130_fd_sc_hd__o21a_1 _12482_ (.A1(_05019_),
    .A2(_05647_),
    .B1(_05009_),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_05218_),
    .X(_05649_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_05218_),
    .X(_05650_));
 sky130_fd_sc_hd__mux2_1 _12485_ (.A0(_05649_),
    .A1(_05650_),
    .S(_05002_),
    .X(_05651_));
 sky130_fd_sc_hd__a221o_1 _12486_ (.A1(_05646_),
    .A2(_05648_),
    .B1(_05651_),
    .B2(_05034_),
    .C1(_05023_),
    .X(_05652_));
 sky130_fd_sc_hd__o311a_1 _12487_ (.A1(_04978_),
    .A2(_05640_),
    .A3(_05644_),
    .B1(_05652_),
    .C1(_05051_),
    .X(_05653_));
 sky130_fd_sc_hd__a31o_1 _12488_ (.A1(_05028_),
    .A2(_05628_),
    .A3(_05636_),
    .B1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_05263_),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_05219_),
    .X(_05656_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(_05655_),
    .A1(_05656_),
    .S(_05069_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_05457_),
    .X(_05658_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_05262_),
    .X(_05659_));
 sky130_fd_sc_hd__or2_1 _12494_ (.A(_05229_),
    .B(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__o211a_1 _12495_ (.A1(_05279_),
    .A2(_05658_),
    .B1(_05660_),
    .C1(_05461_),
    .X(_05661_));
 sky130_fd_sc_hd__a211o_1 _12496_ (.A1(_05035_),
    .A2(_05657_),
    .B1(_05661_),
    .C1(_04979_),
    .X(_05662_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_05263_),
    .X(_05663_));
 sky130_fd_sc_hd__mux2_1 _12498_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_05219_),
    .X(_05664_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(_05663_),
    .A1(_05664_),
    .S(_05235_),
    .X(_05665_));
 sky130_fd_sc_hd__mux2_1 _12500_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_05457_),
    .X(_05666_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_05262_),
    .X(_05667_));
 sky130_fd_sc_hd__or2_1 _12502_ (.A(_05229_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__o211a_1 _12503_ (.A1(_05279_),
    .A2(_05666_),
    .B1(_05668_),
    .C1(_05461_),
    .X(_05669_));
 sky130_fd_sc_hd__a211o_1 _12504_ (.A1(_05035_),
    .A2(_05665_),
    .B1(_05669_),
    .C1(_05030_),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_05219_),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_05071_),
    .X(_05672_));
 sky130_fd_sc_hd__or2_1 _12507_ (.A(_05068_),
    .B(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__o211a_1 _12508_ (.A1(_05235_),
    .A2(_05671_),
    .B1(_05673_),
    .C1(_05061_),
    .X(_05674_));
 sky130_fd_sc_hd__mux2_1 _12509_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_05263_),
    .X(_05675_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_05230_),
    .X(_05676_));
 sky130_fd_sc_hd__or2_1 _12511_ (.A(_05229_),
    .B(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__o211a_1 _12512_ (.A1(_05279_),
    .A2(_05675_),
    .B1(_05677_),
    .C1(_05244_),
    .X(_05678_));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_05230_),
    .X(_05679_));
 sky130_fd_sc_hd__or2_1 _12514_ (.A(_05229_),
    .B(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_05456_),
    .X(_05681_));
 sky130_fd_sc_hd__o21a_1 _12516_ (.A1(_04993_),
    .A2(_05681_),
    .B1(_04999_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _12517_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_05218_),
    .X(_05683_));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_05218_),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_1 _12519_ (.A0(_05683_),
    .A1(_05684_),
    .S(_05068_),
    .X(_05685_));
 sky130_fd_sc_hd__a221o_1 _12520_ (.A1(_05680_),
    .A2(_05682_),
    .B1(_05685_),
    .B2(_05061_),
    .C1(net81),
    .X(_05686_));
 sky130_fd_sc_hd__o311a_1 _12521_ (.A1(_05023_),
    .A2(_05674_),
    .A3(_05678_),
    .B1(_05686_),
    .C1(_05051_),
    .X(_05687_));
 sky130_fd_sc_hd__a31o_1 _12522_ (.A1(_05028_),
    .A2(_05662_),
    .A3(_05670_),
    .B1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_2 _12523_ (.A0(_05654_),
    .A1(_05688_),
    .S(_04975_),
    .X(_05689_));
 sky130_fd_sc_hd__a2bb2o_1 _12524_ (.A1_N(_05117_),
    .A2_N(_05620_),
    .B1(_05689_),
    .B2(_04909_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(net4081),
    .A1(net987),
    .S(_05120_),
    .X(_05691_));
 sky130_fd_sc_hd__mux2_2 _12526_ (.A0(_05690_),
    .A1(net4082),
    .S(net4077),
    .X(_05692_));
 sky130_fd_sc_hd__o21ai_1 _12527_ (.A1(_05309_),
    .A2(_05318_),
    .B1(_05611_),
    .Y(_05693_));
 sky130_fd_sc_hd__a21o_1 _12528_ (.A1(_04906_),
    .A2(_05693_),
    .B1(_04842_),
    .X(_05694_));
 sky130_fd_sc_hd__nand2_1 _12529_ (.A(_05189_),
    .B(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__o21ai_2 _12530_ (.A1(_04818_),
    .A2(net3535),
    .B1(net2),
    .Y(_05696_));
 sky130_fd_sc_hd__o211a_1 _12531_ (.A1(_05189_),
    .A2(_05692_),
    .B1(_05695_),
    .C1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__o21a_1 _12532_ (.A1(net83),
    .A2(_05697_),
    .B1(net4044),
    .X(_05698_));
 sky130_fd_sc_hd__mux2_2 _12533_ (.A0(\reg_rgb[22] ),
    .A1(_05698_),
    .S(_05204_),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_1 _12534_ (.A(_05699_),
    .X(net68));
 sky130_fd_sc_hd__nor2_1 _12535_ (.A(net4093),
    .B(_05693_),
    .Y(_05700_));
 sky130_fd_sc_hd__mux2_1 _12536_ (.A0(net947),
    .A1(net3128),
    .S(_05120_),
    .X(_05701_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04989_),
    .X(_05702_));
 sky130_fd_sc_hd__mux2_1 _12538_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_05541_),
    .X(_05703_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(_05702_),
    .A1(_05703_),
    .S(_05261_),
    .X(_05704_));
 sky130_fd_sc_hd__mux2_1 _12540_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04989_),
    .X(_05705_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04988_),
    .X(_05706_));
 sky130_fd_sc_hd__or2_1 _12542_ (.A(_05003_),
    .B(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__o211a_1 _12543_ (.A1(_04984_),
    .A2(_05705_),
    .B1(_05707_),
    .C1(_05035_),
    .X(_05708_));
 sky130_fd_sc_hd__a211o_1 _12544_ (.A1(_05062_),
    .A2(_05704_),
    .B1(_05708_),
    .C1(_04979_),
    .X(_05709_));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_05541_),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_05541_),
    .X(_05711_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(_05710_),
    .A1(_05711_),
    .S(_05177_),
    .X(_05712_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04989_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04994_),
    .X(_05714_));
 sky130_fd_sc_hd__or2_1 _12550_ (.A(_04983_),
    .B(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__o211a_1 _12551_ (.A1(_05004_),
    .A2(_05713_),
    .B1(_05715_),
    .C1(_05010_),
    .X(_05716_));
 sky130_fd_sc_hd__a211o_1 _12552_ (.A1(_05035_),
    .A2(_05712_),
    .B1(_05716_),
    .C1(_05030_),
    .X(_05717_));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_05541_),
    .X(_05718_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04994_),
    .X(_05719_));
 sky130_fd_sc_hd__or2_1 _12555_ (.A(_04983_),
    .B(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__o211a_1 _12556_ (.A1(_05177_),
    .A2(_05718_),
    .B1(_05720_),
    .C1(_05461_),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _12557_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04989_),
    .X(_05722_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_04994_),
    .X(_05723_));
 sky130_fd_sc_hd__or2_1 _12559_ (.A(_04983_),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__o211a_1 _12560_ (.A1(_05004_),
    .A2(_05722_),
    .B1(_05724_),
    .C1(_05000_),
    .X(_05725_));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04994_),
    .X(_05726_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04994_),
    .X(_05727_));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(_05726_),
    .A1(_05727_),
    .S(_05019_),
    .X(_05728_));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04988_),
    .X(_05729_));
 sky130_fd_sc_hd__or2_1 _12565_ (.A(_04983_),
    .B(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_05014_),
    .X(_05731_));
 sky130_fd_sc_hd__o21a_1 _12567_ (.A1(_05003_),
    .A2(_05731_),
    .B1(_05009_),
    .X(_05732_));
 sky130_fd_sc_hd__a221o_1 _12568_ (.A1(_05000_),
    .A2(_05728_),
    .B1(_05730_),
    .B2(_05732_),
    .C1(_05023_),
    .X(_05733_));
 sky130_fd_sc_hd__o311a_1 _12569_ (.A1(_04979_),
    .A2(_05721_),
    .A3(_05725_),
    .B1(_05028_),
    .C1(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__a31o_1 _12570_ (.A1(_05051_),
    .A2(_05709_),
    .A3(_05717_),
    .B1(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_05476_),
    .X(_05736_));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_05476_),
    .X(_05737_));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(_05736_),
    .A1(_05737_),
    .S(_05279_),
    .X(_05738_));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_05541_),
    .X(_05739_));
 sky130_fd_sc_hd__or2_1 _12575_ (.A(_05177_),
    .B(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__mux2_1 _12576_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04989_),
    .X(_05741_));
 sky130_fd_sc_hd__o21a_1 _12577_ (.A1(_04984_),
    .A2(_05741_),
    .B1(_05000_),
    .X(_05742_));
 sky130_fd_sc_hd__a221o_1 _12578_ (.A1(_05062_),
    .A2(_05738_),
    .B1(_05740_),
    .B2(_05742_),
    .C1(_05030_),
    .X(_05743_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_05476_),
    .X(_05744_));
 sky130_fd_sc_hd__mux2_1 _12580_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_05476_),
    .X(_05745_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(_05744_),
    .A1(_05745_),
    .S(_05261_),
    .X(_05746_));
 sky130_fd_sc_hd__mux2_1 _12582_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_05541_),
    .X(_05747_));
 sky130_fd_sc_hd__or2_1 _12583_ (.A(_04984_),
    .B(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04989_),
    .X(_05749_));
 sky130_fd_sc_hd__o21a_1 _12585_ (.A1(_05004_),
    .A2(_05749_),
    .B1(_05461_),
    .X(_05750_));
 sky130_fd_sc_hd__a221o_1 _12586_ (.A1(_05035_),
    .A2(_05746_),
    .B1(_05748_),
    .B2(_05750_),
    .C1(_04979_),
    .X(_05751_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_05541_),
    .X(_05752_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_05483_),
    .X(_05753_));
 sky130_fd_sc_hd__or2_1 _12589_ (.A(_05019_),
    .B(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__o211a_1 _12590_ (.A1(_05177_),
    .A2(_05752_),
    .B1(_05754_),
    .C1(_05000_),
    .X(_05755_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04989_),
    .X(_05756_));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04994_),
    .X(_05757_));
 sky130_fd_sc_hd__or2_1 _12593_ (.A(_04983_),
    .B(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__o211a_1 _12594_ (.A1(_05177_),
    .A2(_05756_),
    .B1(_05758_),
    .C1(_05010_),
    .X(_05759_));
 sky130_fd_sc_hd__mux2_1 _12595_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04988_),
    .X(_05760_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04988_),
    .X(_05761_));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(_05760_),
    .A1(_05761_),
    .S(_04993_),
    .X(_05762_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_05014_),
    .X(_05763_));
 sky130_fd_sc_hd__mux2_1 _12599_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04987_),
    .X(_05764_));
 sky130_fd_sc_hd__or2_1 _12600_ (.A(_05068_),
    .B(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__o211a_1 _12601_ (.A1(_05003_),
    .A2(_05763_),
    .B1(_05765_),
    .C1(_05061_),
    .X(_05766_));
 sky130_fd_sc_hd__a211o_1 _12602_ (.A1(_05035_),
    .A2(_05762_),
    .B1(_05766_),
    .C1(_05023_),
    .X(_05767_));
 sky130_fd_sc_hd__o311a_1 _12603_ (.A1(_04979_),
    .A2(_05755_),
    .A3(_05759_),
    .B1(_05028_),
    .C1(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__a31o_1 _12604_ (.A1(_05051_),
    .A2(_05743_),
    .A3(_05751_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(_05735_),
    .A1(_05769_),
    .S(_04975_),
    .X(_05770_));
 sky130_fd_sc_hd__o21ai_1 _12606_ (.A1(net4239),
    .A2(_05097_),
    .B1(_05209_),
    .Y(_05771_));
 sky130_fd_sc_hd__a21o_1 _12607_ (.A1(net4239),
    .A2(_05097_),
    .B1(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__a2bb2o_1 _12608_ (.A1_N(net4239),
    .A2_N(_05102_),
    .B1(_04984_),
    .B2(_05035_),
    .X(_05773_));
 sky130_fd_sc_hd__a211o_1 _12609_ (.A1(_05208_),
    .A2(_05773_),
    .B1(_05619_),
    .C1(_05095_),
    .X(_05774_));
 sky130_fd_sc_hd__a31o_1 _12610_ (.A1(net42),
    .A2(_05772_),
    .A3(_05774_),
    .B1(net4077),
    .X(_05775_));
 sky130_fd_sc_hd__o21ba_1 _12611_ (.A1(_05207_),
    .A2(_05770_),
    .B1_N(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__a211o_1 _12612_ (.A1(net4077),
    .A2(_05701_),
    .B1(_05776_),
    .C1(_05189_),
    .X(_05777_));
 sky130_fd_sc_hd__o211a_1 _12613_ (.A1(_04858_),
    .A2(_05700_),
    .B1(_05777_),
    .C1(_05696_),
    .X(_05778_));
 sky130_fd_sc_hd__o21a_1 _12614_ (.A1(net83),
    .A2(_05778_),
    .B1(net4006),
    .X(_05779_));
 sky130_fd_sc_hd__mux2_2 _12615_ (.A0(\reg_rgb[23] ),
    .A1(_05779_),
    .S(_05204_),
    .X(_05780_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_05780_),
    .X(net69));
 sky130_fd_sc_hd__mux2_2 _12617_ (.A0(reg_vsync),
    .A1(_04620_),
    .S(_05204_),
    .X(_05781_));
 sky130_fd_sc_hd__clkbuf_2 _12618_ (.A(_05781_),
    .X(net76));
 sky130_fd_sc_hd__inv_2 _12619_ (.A(\rbzero.hsync ),
    .Y(_05782_));
 sky130_fd_sc_hd__mux2_2 _12620_ (.A0(reg_hsync),
    .A1(_05782_),
    .S(_05204_),
    .X(_05783_));
 sky130_fd_sc_hd__buf_1 _12621_ (.A(_05783_),
    .X(net64));
 sky130_fd_sc_hd__nor2_1 _12622_ (.A(net9),
    .B(net8),
    .Y(_05784_));
 sky130_fd_sc_hd__nor2_2 _12623_ (.A(net7),
    .B(net6),
    .Y(_05785_));
 sky130_fd_sc_hd__nor2_2 _12624_ (.A(net5),
    .B(net4),
    .Y(_05786_));
 sky130_fd_sc_hd__and2_1 _12625_ (.A(_05785_),
    .B(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__nand2_1 _12626_ (.A(_05784_),
    .B(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__mux4_1 _12627_ (.A0(net4045),
    .A1(net4066),
    .A2(net4083),
    .A3(net4078),
    .S0(net4),
    .S1(net7),
    .X(_05789_));
 sky130_fd_sc_hd__inv_2 _12628_ (.A(net7),
    .Y(_05790_));
 sky130_fd_sc_hd__nor2_1 _12629_ (.A(_05790_),
    .B(net8),
    .Y(_05791_));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(net4095),
    .A1(_05446_),
    .S(net4),
    .X(_05792_));
 sky130_fd_sc_hd__a22o_1 _12631_ (.A1(net8),
    .A2(_05789_),
    .B1(_05791_),
    .B2(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__and4b_1 _12632_ (.A_N(net9),
    .B(_05793_),
    .C(net5),
    .D(net6),
    .X(_05794_));
 sky130_fd_sc_hd__nor2b_2 _12633_ (.A(net4),
    .B_N(net5),
    .Y(_05795_));
 sky130_fd_sc_hd__and2b_2 _12634_ (.A_N(net5),
    .B(net4),
    .X(_05796_));
 sky130_fd_sc_hd__a22o_1 _12635_ (.A1(net54),
    .A2(_05786_),
    .B1(_05796_),
    .B2(net55),
    .X(_05797_));
 sky130_fd_sc_hd__a21o_1 _12636_ (.A1(net57),
    .A2(_05795_),
    .B1(_05797_),
    .X(_05798_));
 sky130_fd_sc_hd__and2_2 _12637_ (.A(net5),
    .B(net4),
    .X(_05799_));
 sky130_fd_sc_hd__and3_2 _12638_ (.A(clknet_leaf_69_i_clk),
    .B(_05785_),
    .C(_05795_),
    .X(_05800_));
 sky130_fd_sc_hd__a41o_2 _12639_ (.A1(net56),
    .A2(_05790_),
    .A3(net6),
    .A4(_05799_),
    .B1(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__a31o_2 _12640_ (.A1(_04241_),
    .A2(_05785_),
    .A3(_05796_),
    .B1(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__a311o_2 _12641_ (.A1(net6349),
    .A2(_05785_),
    .A3(_05799_),
    .B1(_05802_),
    .C1(_05787_),
    .X(_05803_));
 sky130_fd_sc_hd__a31o_2 _12642_ (.A1(_05790_),
    .A2(net6),
    .A3(_05798_),
    .B1(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__a22o_1 _12643_ (.A1(_05201_),
    .A2(_05786_),
    .B1(_05796_),
    .B2(net73),
    .X(_05805_));
 sky130_fd_sc_hd__and3_1 _12644_ (.A(_05790_),
    .B(net6),
    .C(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__a22o_1 _12645_ (.A1(net51),
    .A2(_05795_),
    .B1(_05799_),
    .B2(net52),
    .X(_05807_));
 sky130_fd_sc_hd__a32o_1 _12646_ (.A1(net46),
    .A2(_05785_),
    .A3(_05796_),
    .B1(_05787_),
    .B2(net43),
    .X(_05808_));
 sky130_fd_sc_hd__and3_1 _12647_ (.A(net4043),
    .B(_05785_),
    .C(_05799_),
    .X(_05809_));
 sky130_fd_sc_hd__a311o_1 _12648_ (.A1(net44),
    .A2(_05785_),
    .A3(_05795_),
    .B1(_05808_),
    .C1(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__a22o_1 _12649_ (.A1(net53),
    .A2(_05786_),
    .B1(_05796_),
    .B2(net40),
    .X(_05811_));
 sky130_fd_sc_hd__a221o_1 _12650_ (.A1(net41),
    .A2(_05795_),
    .B1(_05799_),
    .B2(_05207_),
    .C1(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__and3b_1 _12651_ (.A_N(net6),
    .B(_05812_),
    .C(net7),
    .X(_05813_));
 sky130_fd_sc_hd__a311o_1 _12652_ (.A1(_05790_),
    .A2(net6),
    .A3(_05807_),
    .B1(_05810_),
    .C1(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__o21ba_1 _12653_ (.A1(_05806_),
    .A2(_05814_),
    .B1_N(net8),
    .X(_05815_));
 sky130_fd_sc_hd__buf_4 _12654_ (.A(net4034),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_1 _12655_ (.A(net4020),
    .X(_05817_));
 sky130_fd_sc_hd__a22o_1 _12656_ (.A1(net4021),
    .A2(_05786_),
    .B1(_05796_),
    .B2(_05299_),
    .X(_05818_));
 sky130_fd_sc_hd__a221o_1 _12657_ (.A1(_05816_),
    .A2(_05795_),
    .B1(_05799_),
    .B2(net4060),
    .C1(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__a21oi_1 _12658_ (.A1(net5),
    .A2(net6),
    .B1(net7),
    .Y(_05820_));
 sky130_fd_sc_hd__a22o_1 _12659_ (.A1(net6),
    .A2(_05791_),
    .B1(_05820_),
    .B2(net8),
    .X(_05821_));
 sky130_fd_sc_hd__mux4_1 _12660_ (.A0(_04760_),
    .A1(_04603_),
    .A2(_04637_),
    .A3(_04165_),
    .S0(net4),
    .S1(net5),
    .X(_05822_));
 sky130_fd_sc_hd__a32o_1 _12661_ (.A1(net7),
    .A2(net8),
    .A3(_05819_),
    .B1(_05821_),
    .B2(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__buf_1 _12662_ (.A(net6287),
    .X(_05824_));
 sky130_fd_sc_hd__buf_4 _12663_ (.A(net6265),
    .X(_05825_));
 sky130_fd_sc_hd__a22o_1 _12664_ (.A1(net3965),
    .A2(_05795_),
    .B1(_05799_),
    .B2(_05825_),
    .X(_05826_));
 sky130_fd_sc_hd__clkbuf_1 _12665_ (.A(net6041),
    .X(_05827_));
 sky130_fd_sc_hd__clkbuf_1 _12666_ (.A(net6220),
    .X(_05828_));
 sky130_fd_sc_hd__clkbuf_1 _12667_ (.A(net5957),
    .X(_05829_));
 sky130_fd_sc_hd__a22o_1 _12668_ (.A1(_04802_),
    .A2(_05786_),
    .B1(_05796_),
    .B2(net4002),
    .X(_05830_));
 sky130_fd_sc_hd__a221o_1 _12669_ (.A1(net3930),
    .A2(_05795_),
    .B1(_05799_),
    .B2(net3937),
    .C1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(_05826_),
    .A1(_05831_),
    .S(net7),
    .X(_05832_));
 sky130_fd_sc_hd__mux2_1 _12671_ (.A0(_04162_),
    .A1(net3993),
    .S(net4),
    .X(_05833_));
 sky130_fd_sc_hd__mux4_1 _12672_ (.A0(_04159_),
    .A1(_04718_),
    .A2(_04726_),
    .A3(_04777_),
    .S0(net4),
    .S1(net5),
    .X(_05834_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(_05833_),
    .A1(_05834_),
    .S(net7),
    .X(_05835_));
 sky130_fd_sc_hd__a22o_1 _12674_ (.A1(net8),
    .A2(_05832_),
    .B1(_05835_),
    .B2(_05821_),
    .X(_05836_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(_05823_),
    .A1(_05836_),
    .S(net6),
    .X(_05837_));
 sky130_fd_sc_hd__o21a_1 _12676_ (.A1(_05815_),
    .A2(_05837_),
    .B1(net9),
    .X(_05838_));
 sky130_fd_sc_hd__a21o_2 _12677_ (.A1(_05784_),
    .A2(_05804_),
    .B1(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__o22a_2 _12678_ (.A1(net4045),
    .A2(_05788_),
    .B1(_05794_),
    .B2(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_2 _12679_ (.A0(\reg_gpout[0] ),
    .A1(clknet_1_0__leaf__05840_),
    .S(_05204_),
    .X(_05841_));
 sky130_fd_sc_hd__buf_1 _12680_ (.A(_05841_),
    .X(net58));
 sky130_fd_sc_hd__nor2_1 _12681_ (.A(net14),
    .B(net15),
    .Y(_05842_));
 sky130_fd_sc_hd__nor2_1 _12682_ (.A(net13),
    .B(net12),
    .Y(_05843_));
 sky130_fd_sc_hd__nor2_2 _12683_ (.A(net11),
    .B(net10),
    .Y(_05844_));
 sky130_fd_sc_hd__and2_1 _12684_ (.A(_05843_),
    .B(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__nand2_1 _12685_ (.A(_05842_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__mux4_1 _12686_ (.A0(net4045),
    .A1(net4066),
    .A2(net4083),
    .A3(net4078),
    .S0(net10),
    .S1(net13),
    .X(_05847_));
 sky130_fd_sc_hd__and2b_1 _12687_ (.A_N(net14),
    .B(net13),
    .X(_05848_));
 sky130_fd_sc_hd__mux2_1 _12688_ (.A0(net4095),
    .A1(_05446_),
    .S(net10),
    .X(_05849_));
 sky130_fd_sc_hd__a22o_1 _12689_ (.A1(net14),
    .A2(_05847_),
    .B1(_05848_),
    .B2(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__and4b_1 _12690_ (.A_N(net15),
    .B(_05850_),
    .C(net11),
    .D(net12),
    .X(_05851_));
 sky130_fd_sc_hd__nor2b_2 _12691_ (.A(net11),
    .B_N(net10),
    .Y(_05852_));
 sky130_fd_sc_hd__and2_2 _12692_ (.A(net11),
    .B(net10),
    .X(_05853_));
 sky130_fd_sc_hd__nor2b_2 _12693_ (.A(net10),
    .B_N(net11),
    .Y(_05854_));
 sky130_fd_sc_hd__a22o_1 _12694_ (.A1(net52),
    .A2(_05853_),
    .B1(_05854_),
    .B2(net51),
    .X(_05855_));
 sky130_fd_sc_hd__a221oi_1 _12695_ (.A1(_05201_),
    .A2(_05844_),
    .B1(_05852_),
    .B2(net73),
    .C1(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _12696_ (.A(net53),
    .B(_05844_),
    .Y(_05857_));
 sky130_fd_sc_hd__a22o_1 _12697_ (.A1(net40),
    .A2(_05852_),
    .B1(_05854_),
    .B2(net41),
    .X(_05858_));
 sky130_fd_sc_hd__a21oi_1 _12698_ (.A1(_05207_),
    .A2(_05853_),
    .B1(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__a31o_1 _12699_ (.A1(net13),
    .A2(_05857_),
    .A3(_05859_),
    .B1(net12),
    .X(_05860_));
 sky130_fd_sc_hd__o21ai_1 _12700_ (.A1(net13),
    .A2(_05856_),
    .B1(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21bo_1 _12701_ (.A1(net44),
    .A2(_05854_),
    .B1_N(_05843_),
    .X(_05862_));
 sky130_fd_sc_hd__a22o_1 _12702_ (.A1(net43),
    .A2(_05844_),
    .B1(_05852_),
    .B2(net46),
    .X(_05863_));
 sky130_fd_sc_hd__a211o_1 _12703_ (.A1(net4043),
    .A2(_05853_),
    .B1(_05862_),
    .C1(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__and4b_1 _12704_ (.A_N(net14),
    .B(net15),
    .C(_05861_),
    .D(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__a22o_1 _12705_ (.A1(net4021),
    .A2(_05844_),
    .B1(_05852_),
    .B2(_05299_),
    .X(_05866_));
 sky130_fd_sc_hd__a221o_1 _12706_ (.A1(net4060),
    .A2(_05853_),
    .B1(_05854_),
    .B2(_05816_),
    .C1(_05866_),
    .X(_05867_));
 sky130_fd_sc_hd__a21oi_1 _12707_ (.A1(net11),
    .A2(net12),
    .B1(net13),
    .Y(_05868_));
 sky130_fd_sc_hd__a22o_1 _12708_ (.A1(net12),
    .A2(_05848_),
    .B1(_05868_),
    .B2(net14),
    .X(_05869_));
 sky130_fd_sc_hd__mux4_1 _12709_ (.A0(_04760_),
    .A1(_04603_),
    .A2(_04637_),
    .A3(_04165_),
    .S0(net10),
    .S1(net11),
    .X(_05870_));
 sky130_fd_sc_hd__a32o_1 _12710_ (.A1(net13),
    .A2(net14),
    .A3(_05867_),
    .B1(_05869_),
    .B2(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__a22o_1 _12711_ (.A1(_05825_),
    .A2(_05853_),
    .B1(_05854_),
    .B2(net3965),
    .X(_05872_));
 sky130_fd_sc_hd__a22o_1 _12712_ (.A1(_04802_),
    .A2(_05844_),
    .B1(_05852_),
    .B2(net4002),
    .X(_05873_));
 sky130_fd_sc_hd__a221o_1 _12713_ (.A1(net3937),
    .A2(_05853_),
    .B1(_05854_),
    .B2(net3930),
    .C1(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(_05872_),
    .A1(_05874_),
    .S(net13),
    .X(_05875_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(_04162_),
    .A1(net3993),
    .S(net10),
    .X(_05876_));
 sky130_fd_sc_hd__mux4_1 _12716_ (.A0(_04159_),
    .A1(_04718_),
    .A2(_04726_),
    .A3(_04777_),
    .S0(net10),
    .S1(net11),
    .X(_05877_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(_05876_),
    .A1(_05877_),
    .S(net13),
    .X(_05878_));
 sky130_fd_sc_hd__a22o_1 _12718_ (.A1(net14),
    .A2(_05875_),
    .B1(_05878_),
    .B2(_05869_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_1 _12719_ (.A0(_05871_),
    .A1(_05879_),
    .S(net12),
    .X(_05880_));
 sky130_fd_sc_hd__a22o_1 _12720_ (.A1(net54),
    .A2(_05844_),
    .B1(_05852_),
    .B2(net55),
    .X(_05881_));
 sky130_fd_sc_hd__a21o_1 _12721_ (.A1(net57),
    .A2(_05854_),
    .B1(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__and2b_1 _12722_ (.A_N(net13),
    .B(net12),
    .X(_05883_));
 sky130_fd_sc_hd__and3_2 _12723_ (.A(clknet_1_1__leaf__04800_),
    .B(_05843_),
    .C(_05854_),
    .X(_05884_));
 sky130_fd_sc_hd__a31o_2 _12724_ (.A1(net50),
    .A2(_05843_),
    .A3(_05852_),
    .B1(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__a22o_1 _12725_ (.A1(net6555),
    .A2(_05843_),
    .B1(_05883_),
    .B2(net56),
    .X(_05886_));
 sky130_fd_sc_hd__a21o_1 _12726_ (.A1(_05853_),
    .A2(_05886_),
    .B1(_05845_),
    .X(_05887_));
 sky130_fd_sc_hd__a211o_2 _12727_ (.A1(_05882_),
    .A2(_05883_),
    .B1(_05885_),
    .C1(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__a22o_2 _12728_ (.A1(net15),
    .A2(_05880_),
    .B1(_05888_),
    .B2(_05842_),
    .X(_05889_));
 sky130_fd_sc_hd__or2_2 _12729_ (.A(_05865_),
    .B(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__o22a_2 _12730_ (.A1(net4066),
    .A2(_05846_),
    .B1(_05851_),
    .B2(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__mux2_2 _12731_ (.A0(\reg_gpout[1] ),
    .A1(clknet_1_1__leaf__05891_),
    .S(_05204_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _12732_ (.A(_05892_),
    .X(net59));
 sky130_fd_sc_hd__nor2_1 _12733_ (.A(net21),
    .B(net20),
    .Y(_05893_));
 sky130_fd_sc_hd__nor2_1 _12734_ (.A(net19),
    .B(net18),
    .Y(_05894_));
 sky130_fd_sc_hd__nor2_2 _12735_ (.A(net17),
    .B(net16),
    .Y(_05895_));
 sky130_fd_sc_hd__and2_1 _12736_ (.A(_05894_),
    .B(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__nand2_1 _12737_ (.A(_05893_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__mux4_1 _12738_ (.A0(net4045),
    .A1(net4066),
    .A2(net4083),
    .A3(net4078),
    .S0(net16),
    .S1(net19),
    .X(_05898_));
 sky130_fd_sc_hd__and2b_1 _12739_ (.A_N(net20),
    .B(net19),
    .X(_05899_));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(net4095),
    .A1(_05446_),
    .S(net16),
    .X(_05900_));
 sky130_fd_sc_hd__a22o_1 _12741_ (.A1(net20),
    .A2(_05898_),
    .B1(_05899_),
    .B2(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__and4b_1 _12742_ (.A_N(net21),
    .B(_05901_),
    .C(net17),
    .D(net18),
    .X(_05902_));
 sky130_fd_sc_hd__nor2b_2 _12743_ (.A(net17),
    .B_N(net16),
    .Y(_05903_));
 sky130_fd_sc_hd__and2_2 _12744_ (.A(net17),
    .B(net16),
    .X(_05904_));
 sky130_fd_sc_hd__nor2b_2 _12745_ (.A(net16),
    .B_N(net17),
    .Y(_05905_));
 sky130_fd_sc_hd__a22o_1 _12746_ (.A1(net52),
    .A2(_05904_),
    .B1(_05905_),
    .B2(net51),
    .X(_05906_));
 sky130_fd_sc_hd__a221oi_1 _12747_ (.A1(_05201_),
    .A2(_05895_),
    .B1(_05903_),
    .B2(net73),
    .C1(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_1 _12748_ (.A(net53),
    .B(_05895_),
    .Y(_05908_));
 sky130_fd_sc_hd__a22o_1 _12749_ (.A1(net40),
    .A2(_05903_),
    .B1(_05905_),
    .B2(net41),
    .X(_05909_));
 sky130_fd_sc_hd__a21oi_1 _12750_ (.A1(_05207_),
    .A2(_05904_),
    .B1(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__a31o_1 _12751_ (.A1(net19),
    .A2(_05908_),
    .A3(_05910_),
    .B1(net18),
    .X(_05911_));
 sky130_fd_sc_hd__o21ai_1 _12752_ (.A1(net19),
    .A2(_05907_),
    .B1(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__a21bo_1 _12753_ (.A1(net44),
    .A2(_05905_),
    .B1_N(_05894_),
    .X(_05913_));
 sky130_fd_sc_hd__a22o_1 _12754_ (.A1(net43),
    .A2(_05895_),
    .B1(_05903_),
    .B2(net46),
    .X(_05914_));
 sky130_fd_sc_hd__a211o_1 _12755_ (.A1(net4043),
    .A2(_05904_),
    .B1(_05913_),
    .C1(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__and4b_1 _12756_ (.A_N(net20),
    .B(_05912_),
    .C(_05915_),
    .D(net21),
    .X(_05916_));
 sky130_fd_sc_hd__a22o_1 _12757_ (.A1(net4021),
    .A2(_05895_),
    .B1(_05903_),
    .B2(_05299_),
    .X(_05917_));
 sky130_fd_sc_hd__a221o_1 _12758_ (.A1(net4060),
    .A2(_05904_),
    .B1(_05905_),
    .B2(_05816_),
    .C1(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__a21oi_1 _12759_ (.A1(net17),
    .A2(net18),
    .B1(net19),
    .Y(_05919_));
 sky130_fd_sc_hd__a22o_1 _12760_ (.A1(net18),
    .A2(_05899_),
    .B1(_05919_),
    .B2(net20),
    .X(_05920_));
 sky130_fd_sc_hd__mux4_1 _12761_ (.A0(_04760_),
    .A1(_04603_),
    .A2(_04637_),
    .A3(_04165_),
    .S0(net16),
    .S1(net17),
    .X(_05921_));
 sky130_fd_sc_hd__a32o_1 _12762_ (.A1(net19),
    .A2(net20),
    .A3(_05918_),
    .B1(_05920_),
    .B2(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__a22o_1 _12763_ (.A1(_05825_),
    .A2(_05904_),
    .B1(_05905_),
    .B2(net3965),
    .X(_05923_));
 sky130_fd_sc_hd__a22o_1 _12764_ (.A1(_04802_),
    .A2(_05895_),
    .B1(_05903_),
    .B2(net4002),
    .X(_05924_));
 sky130_fd_sc_hd__a221o_1 _12765_ (.A1(net3937),
    .A2(_05904_),
    .B1(_05905_),
    .B2(net3930),
    .C1(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(_05923_),
    .A1(_05925_),
    .S(net19),
    .X(_05926_));
 sky130_fd_sc_hd__mux2_1 _12767_ (.A0(_04162_),
    .A1(net3993),
    .S(net16),
    .X(_05927_));
 sky130_fd_sc_hd__mux4_1 _12768_ (.A0(_04159_),
    .A1(net4891),
    .A2(_04726_),
    .A3(_04777_),
    .S0(net16),
    .S1(net17),
    .X(_05928_));
 sky130_fd_sc_hd__mux2_1 _12769_ (.A0(_05927_),
    .A1(_05928_),
    .S(net19),
    .X(_05929_));
 sky130_fd_sc_hd__a22o_1 _12770_ (.A1(net20),
    .A2(_05926_),
    .B1(_05929_),
    .B2(_05920_),
    .X(_05930_));
 sky130_fd_sc_hd__mux2_1 _12771_ (.A0(_05922_),
    .A1(_05930_),
    .S(net18),
    .X(_05931_));
 sky130_fd_sc_hd__a22o_1 _12772_ (.A1(net54),
    .A2(_05895_),
    .B1(_05903_),
    .B2(net55),
    .X(_05932_));
 sky130_fd_sc_hd__a21o_1 _12773_ (.A1(net57),
    .A2(_05905_),
    .B1(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__and2b_1 _12774_ (.A_N(net19),
    .B(net18),
    .X(_05934_));
 sky130_fd_sc_hd__and3_2 _12775_ (.A(clknet_1_1__leaf__04800_),
    .B(_05894_),
    .C(_05905_),
    .X(_05935_));
 sky130_fd_sc_hd__a31o_2 _12776_ (.A1(net49),
    .A2(_05894_),
    .A3(_05903_),
    .B1(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__a22o_1 _12777_ (.A1(net6355),
    .A2(_05894_),
    .B1(_05934_),
    .B2(net56),
    .X(_05937_));
 sky130_fd_sc_hd__a21o_1 _12778_ (.A1(_05904_),
    .A2(_05937_),
    .B1(_05896_),
    .X(_05938_));
 sky130_fd_sc_hd__a211o_2 _12779_ (.A1(_05933_),
    .A2(_05934_),
    .B1(_05936_),
    .C1(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__a22o_2 _12780_ (.A1(net21),
    .A2(_05931_),
    .B1(_05939_),
    .B2(_05893_),
    .X(_05940_));
 sky130_fd_sc_hd__or2_2 _12781_ (.A(_05916_),
    .B(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__o22a_2 _12782_ (.A1(net4095),
    .A2(_05897_),
    .B1(_05902_),
    .B2(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__mux2_2 _12783_ (.A0(\reg_gpout[2] ),
    .A1(clknet_1_1__leaf__05942_),
    .S(net45),
    .X(_05943_));
 sky130_fd_sc_hd__buf_1 _12784_ (.A(_05943_),
    .X(net60));
 sky130_fd_sc_hd__nor2_1 _12785_ (.A(net26),
    .B(net27),
    .Y(_05944_));
 sky130_fd_sc_hd__nor2_1 _12786_ (.A(net25),
    .B(net24),
    .Y(_05945_));
 sky130_fd_sc_hd__nor2_2 _12787_ (.A(net23),
    .B(net22),
    .Y(_05946_));
 sky130_fd_sc_hd__and2_1 _12788_ (.A(_05945_),
    .B(_05946_),
    .X(_05947_));
 sky130_fd_sc_hd__nand2_1 _12789_ (.A(_05944_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__mux4_1 _12790_ (.A0(net4045),
    .A1(net4066),
    .A2(net4083),
    .A3(net4078),
    .S0(net22),
    .S1(net25),
    .X(_05949_));
 sky130_fd_sc_hd__inv_2 _12791_ (.A(net25),
    .Y(_05950_));
 sky130_fd_sc_hd__nor2_1 _12792_ (.A(_05950_),
    .B(net26),
    .Y(_05951_));
 sky130_fd_sc_hd__mux2_1 _12793_ (.A0(net4095),
    .A1(_05446_),
    .S(net22),
    .X(_05952_));
 sky130_fd_sc_hd__a22o_1 _12794_ (.A1(net26),
    .A2(_05949_),
    .B1(_05951_),
    .B2(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__and4b_1 _12795_ (.A_N(net27),
    .B(_05953_),
    .C(net23),
    .D(net24),
    .X(_05954_));
 sky130_fd_sc_hd__inv_2 _12796_ (.A(net23),
    .Y(_05955_));
 sky130_fd_sc_hd__and2_2 _12797_ (.A(_05955_),
    .B(net22),
    .X(_05956_));
 sky130_fd_sc_hd__and2_2 _12798_ (.A(net23),
    .B(net22),
    .X(_05957_));
 sky130_fd_sc_hd__nor2_2 _12799_ (.A(_05955_),
    .B(net22),
    .Y(_05958_));
 sky130_fd_sc_hd__a22o_1 _12800_ (.A1(net52),
    .A2(_05957_),
    .B1(_05958_),
    .B2(net51),
    .X(_05959_));
 sky130_fd_sc_hd__a221o_1 _12801_ (.A1(_05201_),
    .A2(_05946_),
    .B1(_05956_),
    .B2(net73),
    .C1(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(net53),
    .B(_05946_),
    .Y(_05961_));
 sky130_fd_sc_hd__a22o_1 _12803_ (.A1(net40),
    .A2(_05956_),
    .B1(_05958_),
    .B2(net41),
    .X(_05962_));
 sky130_fd_sc_hd__a21oi_1 _12804_ (.A1(_05207_),
    .A2(_05957_),
    .B1(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a31o_1 _12805_ (.A1(net25),
    .A2(_05961_),
    .A3(_05963_),
    .B1(net24),
    .X(_05964_));
 sky130_fd_sc_hd__a21boi_1 _12806_ (.A1(_05950_),
    .A2(_05960_),
    .B1_N(_05964_),
    .Y(_05965_));
 sky130_fd_sc_hd__a21bo_1 _12807_ (.A1(net44),
    .A2(_05958_),
    .B1_N(_05945_),
    .X(_05966_));
 sky130_fd_sc_hd__a22o_1 _12808_ (.A1(net43),
    .A2(_05946_),
    .B1(_05956_),
    .B2(net46),
    .X(_05967_));
 sky130_fd_sc_hd__a211o_1 _12809_ (.A1(net4043),
    .A2(_05957_),
    .B1(_05966_),
    .C1(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__and4bb_1 _12810_ (.A_N(net26),
    .B_N(_05965_),
    .C(_05968_),
    .D(net27),
    .X(_05969_));
 sky130_fd_sc_hd__a22o_1 _12811_ (.A1(net4021),
    .A2(_05946_),
    .B1(_05956_),
    .B2(_05299_),
    .X(_05970_));
 sky130_fd_sc_hd__a221o_1 _12812_ (.A1(net4060),
    .A2(_05957_),
    .B1(_05958_),
    .B2(_05194_),
    .C1(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__a21oi_1 _12813_ (.A1(net23),
    .A2(net24),
    .B1(net25),
    .Y(_05972_));
 sky130_fd_sc_hd__a22o_1 _12814_ (.A1(net24),
    .A2(_05951_),
    .B1(_05972_),
    .B2(net26),
    .X(_05973_));
 sky130_fd_sc_hd__mux4_1 _12815_ (.A0(_04760_),
    .A1(_04603_),
    .A2(_04637_),
    .A3(_04165_),
    .S0(net22),
    .S1(net23),
    .X(_05974_));
 sky130_fd_sc_hd__a32o_1 _12816_ (.A1(net25),
    .A2(net26),
    .A3(_05971_),
    .B1(_05973_),
    .B2(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__a22o_1 _12817_ (.A1(_05825_),
    .A2(_05957_),
    .B1(_05958_),
    .B2(net3964),
    .X(_05976_));
 sky130_fd_sc_hd__a22o_1 _12818_ (.A1(net4972),
    .A2(_05946_),
    .B1(_05956_),
    .B2(net4002),
    .X(_05977_));
 sky130_fd_sc_hd__a221o_1 _12819_ (.A1(net3937),
    .A2(_05957_),
    .B1(_05958_),
    .B2(net3930),
    .C1(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__mux2_1 _12820_ (.A0(_05976_),
    .A1(_05978_),
    .S(net25),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_1 _12821_ (.A0(_04162_),
    .A1(net3993),
    .S(net22),
    .X(_05980_));
 sky130_fd_sc_hd__mux4_1 _12822_ (.A0(_04159_),
    .A1(net4891),
    .A2(_04726_),
    .A3(_04777_),
    .S0(net22),
    .S1(net23),
    .X(_05981_));
 sky130_fd_sc_hd__mux2_1 _12823_ (.A0(_05980_),
    .A1(_05981_),
    .S(net25),
    .X(_05982_));
 sky130_fd_sc_hd__a22o_1 _12824_ (.A1(net26),
    .A2(_05979_),
    .B1(_05982_),
    .B2(_05973_),
    .X(_05983_));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(_05975_),
    .A1(_05983_),
    .S(net24),
    .X(_05984_));
 sky130_fd_sc_hd__a22o_1 _12826_ (.A1(net54),
    .A2(_05946_),
    .B1(_05956_),
    .B2(net55),
    .X(_05985_));
 sky130_fd_sc_hd__a21o_1 _12827_ (.A1(net57),
    .A2(_05958_),
    .B1(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__and2_1 _12828_ (.A(_05950_),
    .B(net24),
    .X(_05987_));
 sky130_fd_sc_hd__a22o_2 _12829_ (.A1(net48),
    .A2(_05956_),
    .B1(_05958_),
    .B2(clknet_1_1__leaf__04800_),
    .X(_05988_));
 sky130_fd_sc_hd__a22o_1 _12830_ (.A1(net6357),
    .A2(_05945_),
    .B1(_05987_),
    .B2(net56),
    .X(_05989_));
 sky130_fd_sc_hd__a221o_2 _12831_ (.A1(_05945_),
    .A2(_05988_),
    .B1(_05989_),
    .B2(_05957_),
    .C1(_05947_),
    .X(_05990_));
 sky130_fd_sc_hd__a21o_2 _12832_ (.A1(_05986_),
    .A2(_05987_),
    .B1(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__a22o_2 _12833_ (.A1(net27),
    .A2(_05984_),
    .B1(_05991_),
    .B2(_05944_),
    .X(_05992_));
 sky130_fd_sc_hd__or2_2 _12834_ (.A(_05969_),
    .B(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__o22a_2 _12835_ (.A1(_05446_),
    .A2(_05948_),
    .B1(_05954_),
    .B2(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__mux2_2 _12836_ (.A0(\reg_gpout[3] ),
    .A1(clknet_1_1__leaf__05994_),
    .S(net45),
    .X(_05995_));
 sky130_fd_sc_hd__buf_1 _12837_ (.A(_05995_),
    .X(net61));
 sky130_fd_sc_hd__nor2_1 _12838_ (.A(net32),
    .B(net33),
    .Y(_05996_));
 sky130_fd_sc_hd__nor2_1 _12839_ (.A(net31),
    .B(net30),
    .Y(_05997_));
 sky130_fd_sc_hd__nor2_2 _12840_ (.A(net29),
    .B(net28),
    .Y(_05998_));
 sky130_fd_sc_hd__and2_1 _12841_ (.A(_05997_),
    .B(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__nand2_1 _12842_ (.A(_05996_),
    .B(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__mux4_1 _12843_ (.A0(net4045),
    .A1(net4066),
    .A2(net4083),
    .A3(net4078),
    .S0(net28),
    .S1(net31),
    .X(_06001_));
 sky130_fd_sc_hd__inv_2 _12844_ (.A(net31),
    .Y(_06002_));
 sky130_fd_sc_hd__nor2_1 _12845_ (.A(_06002_),
    .B(net32),
    .Y(_06003_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(net4095),
    .A1(_05446_),
    .S(net28),
    .X(_06004_));
 sky130_fd_sc_hd__a22o_1 _12847_ (.A1(net32),
    .A2(_06001_),
    .B1(_06003_),
    .B2(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__and4b_1 _12848_ (.A_N(net33),
    .B(_06005_),
    .C(net29),
    .D(net30),
    .X(_06006_));
 sky130_fd_sc_hd__nor2b_2 _12849_ (.A(net29),
    .B_N(net28),
    .Y(_06007_));
 sky130_fd_sc_hd__nor2b_2 _12850_ (.A(net28),
    .B_N(net29),
    .Y(_06008_));
 sky130_fd_sc_hd__and3_1 _12851_ (.A(_05207_),
    .B(net29),
    .C(net28),
    .X(_06009_));
 sky130_fd_sc_hd__a221o_1 _12852_ (.A1(net40),
    .A2(_06007_),
    .B1(_06008_),
    .B2(net41),
    .C1(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__a211oi_1 _12853_ (.A1(net53),
    .A2(_05998_),
    .B1(_06010_),
    .C1(_06002_),
    .Y(_06011_));
 sky130_fd_sc_hd__and2_2 _12854_ (.A(net29),
    .B(net28),
    .X(_06012_));
 sky130_fd_sc_hd__a22o_1 _12855_ (.A1(net52),
    .A2(_06012_),
    .B1(_06008_),
    .B2(net51),
    .X(_06013_));
 sky130_fd_sc_hd__a221o_1 _12856_ (.A1(_05201_),
    .A2(_05998_),
    .B1(_06007_),
    .B2(net73),
    .C1(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__a2bb2o_1 _12857_ (.A1_N(net30),
    .A2_N(_06011_),
    .B1(_06014_),
    .B2(_06002_),
    .X(_06015_));
 sky130_fd_sc_hd__a21bo_1 _12858_ (.A1(net44),
    .A2(_06008_),
    .B1_N(_05997_),
    .X(_06016_));
 sky130_fd_sc_hd__a22o_1 _12859_ (.A1(net43),
    .A2(_05998_),
    .B1(_06007_),
    .B2(net46),
    .X(_06017_));
 sky130_fd_sc_hd__a211o_1 _12860_ (.A1(net4043),
    .A2(_06012_),
    .B1(_06016_),
    .C1(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__and4b_1 _12861_ (.A_N(net32),
    .B(net33),
    .C(_06015_),
    .D(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_1 _12862_ (.A1(net4021),
    .A2(_05998_),
    .B1(_06007_),
    .B2(_05299_),
    .X(_06020_));
 sky130_fd_sc_hd__a221o_1 _12863_ (.A1(net4060),
    .A2(_06012_),
    .B1(_06008_),
    .B2(_05194_),
    .C1(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__a21oi_1 _12864_ (.A1(net29),
    .A2(net30),
    .B1(net31),
    .Y(_06022_));
 sky130_fd_sc_hd__a22o_1 _12865_ (.A1(net30),
    .A2(_06003_),
    .B1(_06022_),
    .B2(net32),
    .X(_06023_));
 sky130_fd_sc_hd__mux4_1 _12866_ (.A0(_04760_),
    .A1(_04603_),
    .A2(_04637_),
    .A3(_04165_),
    .S0(net28),
    .S1(net29),
    .X(_06024_));
 sky130_fd_sc_hd__a32o_1 _12867_ (.A1(net31),
    .A2(net32),
    .A3(_06021_),
    .B1(_06023_),
    .B2(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__a22o_1 _12868_ (.A1(net6265),
    .A2(_06012_),
    .B1(_06008_),
    .B2(net3964),
    .X(_06026_));
 sky130_fd_sc_hd__a22o_1 _12869_ (.A1(net4972),
    .A2(_05998_),
    .B1(_06007_),
    .B2(net4002),
    .X(_06027_));
 sky130_fd_sc_hd__a221o_1 _12870_ (.A1(net3937),
    .A2(_06012_),
    .B1(_06008_),
    .B2(net3930),
    .C1(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(_06026_),
    .A1(_06028_),
    .S(net31),
    .X(_06029_));
 sky130_fd_sc_hd__mux2_1 _12872_ (.A0(_04161_),
    .A1(net3993),
    .S(net28),
    .X(_06030_));
 sky130_fd_sc_hd__mux4_1 _12873_ (.A0(net4049),
    .A1(net4891),
    .A2(_04726_),
    .A3(_04777_),
    .S0(net28),
    .S1(net29),
    .X(_06031_));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(_06030_),
    .A1(_06031_),
    .S(net31),
    .X(_06032_));
 sky130_fd_sc_hd__a22o_1 _12875_ (.A1(net32),
    .A2(_06029_),
    .B1(_06032_),
    .B2(_06023_),
    .X(_06033_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(_06025_),
    .A1(_06033_),
    .S(net30),
    .X(_06034_));
 sky130_fd_sc_hd__a22o_1 _12877_ (.A1(net54),
    .A2(_05998_),
    .B1(_06007_),
    .B2(net55),
    .X(_06035_));
 sky130_fd_sc_hd__a21o_1 _12878_ (.A1(net57),
    .A2(_06008_),
    .B1(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__and2b_1 _12879_ (.A_N(net31),
    .B(net30),
    .X(_06037_));
 sky130_fd_sc_hd__a22o_2 _12880_ (.A1(net3),
    .A2(_06007_),
    .B1(_06008_),
    .B2(clknet_leaf_67_i_clk),
    .X(_06038_));
 sky130_fd_sc_hd__a22o_1 _12881_ (.A1(net6341),
    .A2(_05997_),
    .B1(_06037_),
    .B2(net56),
    .X(_06039_));
 sky130_fd_sc_hd__a221o_2 _12882_ (.A1(_05997_),
    .A2(_06038_),
    .B1(_06039_),
    .B2(_06012_),
    .C1(_05999_),
    .X(_06040_));
 sky130_fd_sc_hd__a21o_2 _12883_ (.A1(_06036_),
    .A2(_06037_),
    .B1(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__a22o_2 _12884_ (.A1(net33),
    .A2(_06034_),
    .B1(_06041_),
    .B2(_05996_),
    .X(_06042_));
 sky130_fd_sc_hd__or2_2 _12885_ (.A(_06019_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__o22a_2 _12886_ (.A1(net4083),
    .A2(_06000_),
    .B1(_06006_),
    .B2(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__mux2_2 _12887_ (.A0(\reg_gpout[4] ),
    .A1(clknet_1_1__leaf__06044_),
    .S(net45),
    .X(_06045_));
 sky130_fd_sc_hd__buf_1 _12888_ (.A(_06045_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 _12889_ (.A(net34),
    .X(_06046_));
 sky130_fd_sc_hd__mux4_1 _12890_ (.A0(net4045),
    .A1(net4066),
    .A2(net4083),
    .A3(net4078),
    .S0(_06046_),
    .S1(net37),
    .X(_06047_));
 sky130_fd_sc_hd__inv_2 _12891_ (.A(net37),
    .Y(_06048_));
 sky130_fd_sc_hd__nor2_1 _12892_ (.A(_06048_),
    .B(net38),
    .Y(_06049_));
 sky130_fd_sc_hd__mux2_1 _12893_ (.A0(net4095),
    .A1(_05446_),
    .S(_06046_),
    .X(_06050_));
 sky130_fd_sc_hd__a22o_1 _12894_ (.A1(net38),
    .A2(_06047_),
    .B1(_06049_),
    .B2(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__buf_2 _12895_ (.A(net35),
    .X(_06052_));
 sky130_fd_sc_hd__and4b_1 _12896_ (.A_N(net39),
    .B(_06051_),
    .C(_06052_),
    .D(net36),
    .X(_06053_));
 sky130_fd_sc_hd__mux4_1 _12897_ (.A0(net54),
    .A1(net55),
    .A2(net57),
    .A3(net56),
    .S0(_06046_),
    .S1(_06052_),
    .X(_06054_));
 sky130_fd_sc_hd__a21oi_2 _12898_ (.A1(net141),
    .A2(_06052_),
    .B1(_06046_),
    .Y(_06055_));
 sky130_fd_sc_hd__and3_1 _12899_ (.A(_06052_),
    .B(_06046_),
    .C(net6347),
    .X(_06056_));
 sky130_fd_sc_hd__or2_1 _12900_ (.A(net37),
    .B(net36),
    .X(_06057_));
 sky130_fd_sc_hd__o21ba_2 _12901_ (.A1(_06055_),
    .A2(_06056_),
    .B1_N(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__a31o_2 _12902_ (.A1(_06048_),
    .A2(net36),
    .A3(_06054_),
    .B1(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__nor2_1 _12903_ (.A(net38),
    .B(net39),
    .Y(_06060_));
 sky130_fd_sc_hd__and3b_1 _12904_ (.A_N(_06046_),
    .B(_06052_),
    .C(net41),
    .X(_06061_));
 sky130_fd_sc_hd__a31o_1 _12905_ (.A1(_05207_),
    .A2(_06052_),
    .A3(_06046_),
    .B1(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__and4b_1 _12906_ (.A_N(net36),
    .B(net39),
    .C(_06049_),
    .D(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__a21o_2 _12907_ (.A1(_06059_),
    .A2(_06060_),
    .B1(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__nor2_1 _12908_ (.A(net35),
    .B(net34),
    .Y(_06065_));
 sky130_fd_sc_hd__and2b_1 _12909_ (.A_N(net35),
    .B(net34),
    .X(_06066_));
 sky130_fd_sc_hd__and3b_1 _12910_ (.A_N(net34),
    .B(net35),
    .C(net51),
    .X(_06067_));
 sky130_fd_sc_hd__a31o_1 _12911_ (.A1(net52),
    .A2(net35),
    .A3(net34),
    .B1(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__a221o_1 _12912_ (.A1(_05201_),
    .A2(_06065_),
    .B1(_06066_),
    .B2(net73),
    .C1(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__a21bo_1 _12913_ (.A1(_06048_),
    .A2(_06069_),
    .B1_N(net36),
    .X(_06070_));
 sky130_fd_sc_hd__nand2_1 _12914_ (.A(net44),
    .B(net35),
    .Y(_06071_));
 sky130_fd_sc_hd__a2bb2o_1 _12915_ (.A1_N(net34),
    .A2_N(_06071_),
    .B1(_06065_),
    .B2(net43),
    .X(_06072_));
 sky130_fd_sc_hd__a31o_1 _12916_ (.A1(net35),
    .A2(_06046_),
    .A3(net4043),
    .B1(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__a211o_1 _12917_ (.A1(net46),
    .A2(_06066_),
    .B1(_06073_),
    .C1(_06057_),
    .X(_06074_));
 sky130_fd_sc_hd__a221o_1 _12918_ (.A1(net53),
    .A2(_06065_),
    .B1(_06066_),
    .B2(net40),
    .C1(_06048_),
    .X(_06075_));
 sky130_fd_sc_hd__and3_1 _12919_ (.A(_06070_),
    .B(_06074_),
    .C(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__mux4_1 _12920_ (.A0(_04160_),
    .A1(_04718_),
    .A2(_04727_),
    .A3(_04777_),
    .S0(_06046_),
    .S1(_06052_),
    .X(_06077_));
 sky130_fd_sc_hd__a31o_1 _12921_ (.A1(net37),
    .A2(net36),
    .A3(_06077_),
    .B1(net38),
    .X(_06078_));
 sky130_fd_sc_hd__mux2_1 _12922_ (.A0(net3965),
    .A1(_05825_),
    .S(_06046_),
    .X(_06079_));
 sky130_fd_sc_hd__mux4_1 _12923_ (.A0(_04760_),
    .A1(_04603_),
    .A2(_04637_),
    .A3(_04165_),
    .S0(net34),
    .S1(net35),
    .X(_06080_));
 sky130_fd_sc_hd__a22o_1 _12924_ (.A1(_04162_),
    .A2(_06065_),
    .B1(_06066_),
    .B2(net3993),
    .X(_06081_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(_06080_),
    .A1(_06081_),
    .S(net36),
    .X(_06082_));
 sky130_fd_sc_hd__a31o_1 _12926_ (.A1(_06052_),
    .A2(net36),
    .A3(_06079_),
    .B1(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__mux4_1 _12927_ (.A0(net4021),
    .A1(_05299_),
    .A2(_04802_),
    .A3(net4002),
    .S0(net34),
    .S1(net36),
    .X(_06084_));
 sky130_fd_sc_hd__mux4_1 _12928_ (.A0(_05194_),
    .A1(net4060),
    .A2(net3930),
    .A3(net3937),
    .S0(net34),
    .S1(net36),
    .X(_06085_));
 sky130_fd_sc_hd__or2b_1 _12929_ (.A(_06085_),
    .B_N(_06052_),
    .X(_06086_));
 sky130_fd_sc_hd__o211a_1 _12930_ (.A1(_06052_),
    .A2(_06084_),
    .B1(_06086_),
    .C1(net37),
    .X(_06087_));
 sky130_fd_sc_hd__a21o_1 _12931_ (.A1(_06048_),
    .A2(_06083_),
    .B1(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(net38),
    .Y(_06089_));
 sky130_fd_sc_hd__o221a_1 _12933_ (.A1(_06076_),
    .A2(_06078_),
    .B1(_06088_),
    .B2(_06089_),
    .C1(net39),
    .X(_06090_));
 sky130_fd_sc_hd__or4bb_1 _12934_ (.A(net4078),
    .B(_06057_),
    .C_N(_06065_),
    .D_N(_06060_),
    .X(_06091_));
 sky130_fd_sc_hd__o31a_2 _12935_ (.A1(_06053_),
    .A2(_06064_),
    .A3(_06090_),
    .B1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__mux2_2 _12936_ (.A0(\reg_gpout[5] ),
    .A1(clknet_1_1__leaf__06092_),
    .S(net45),
    .X(_06093_));
 sky130_fd_sc_hd__buf_1 _12937_ (.A(_06093_),
    .X(net63));
 sky130_fd_sc_hd__or2_1 _12938_ (.A(net3876),
    .B(net3018),
    .X(_06094_));
 sky130_fd_sc_hd__nor2_1 _12939_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06095_));
 sky130_fd_sc_hd__and2_1 _12940_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06096_));
 sky130_fd_sc_hd__nor2_1 _12941_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_06097_));
 sky130_fd_sc_hd__nor2_1 _12942_ (.A(_06096_),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__xor2_2 _12943_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _12944_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06100_));
 sky130_fd_sc_hd__a31o_1 _12945_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_06099_),
    .B1(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__nand2_1 _12946_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06102_));
 sky130_fd_sc_hd__or2b_1 _12947_ (.A(_06096_),
    .B_N(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__a21oi_1 _12948_ (.A1(_06098_),
    .A2(_06101_),
    .B1(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_1 _12949_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_06105_));
 sky130_fd_sc_hd__or2_1 _12950_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_06106_));
 sky130_fd_sc_hd__and2_1 _12951_ (.A(_06105_),
    .B(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__inv_2 _12952_ (.A(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__nand2_1 _12953_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06109_));
 sky130_fd_sc_hd__or2_1 _12954_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_06110_));
 sky130_fd_sc_hd__xor2_2 _12955_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_06111_));
 sky130_fd_sc_hd__nand3_1 _12956_ (.A(_06109_),
    .B(_06110_),
    .C(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_1 _12957_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06113_));
 sky130_fd_sc_hd__nand2_1 _12958_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06114_));
 sky130_fd_sc_hd__or2b_1 _12959_ (.A(_06113_),
    .B_N(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__or2_1 _12960_ (.A(_06112_),
    .B(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__or4_4 _12961_ (.A(_06095_),
    .B(_06104_),
    .C(_06108_),
    .D(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__a21o_1 _12962_ (.A1(_06105_),
    .A2(_06114_),
    .B1(_06113_),
    .X(_06118_));
 sky130_fd_sc_hd__nand2_1 _12963_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06119_));
 sky130_fd_sc_hd__or2b_1 _12964_ (.A(_06119_),
    .B_N(_06110_),
    .X(_06120_));
 sky130_fd_sc_hd__o211a_1 _12965_ (.A1(_06112_),
    .A2(_06118_),
    .B1(_06120_),
    .C1(_06109_),
    .X(_06121_));
 sky130_fd_sc_hd__nand2_1 _12966_ (.A(net4600),
    .B(net3090),
    .Y(_06122_));
 sky130_fd_sc_hd__or2_1 _12967_ (.A(net4600),
    .B(net3090),
    .X(_06123_));
 sky130_fd_sc_hd__nand2_1 _12968_ (.A(_06122_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__a21oi_4 _12969_ (.A1(_06117_),
    .A2(_06121_),
    .B1(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(net3857),
    .B(net3135),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_1 _12971_ (.A(_06122_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__or2_1 _12972_ (.A(net3876),
    .B(net3085),
    .X(_06128_));
 sky130_fd_sc_hd__or2_2 _12973_ (.A(net3857),
    .B(net3135),
    .X(_06129_));
 sky130_fd_sc_hd__o211ai_4 _12974_ (.A1(_06125_),
    .A2(_06127_),
    .B1(_06128_),
    .C1(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__nand2_2 _12975_ (.A(net3876),
    .B(net3085),
    .Y(_06131_));
 sky130_fd_sc_hd__and2_1 _12976_ (.A(net3876),
    .B(net3018),
    .X(_06132_));
 sky130_fd_sc_hd__a31o_1 _12977_ (.A1(_06094_),
    .A2(_06130_),
    .A3(_06131_),
    .B1(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__or2b_1 _12978_ (.A(_06132_),
    .B_N(_06094_),
    .X(_06134_));
 sky130_fd_sc_hd__a21bo_1 _12979_ (.A1(_06130_),
    .A2(_06131_),
    .B1_N(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__inv_2 _12980_ (.A(_06131_),
    .Y(_06136_));
 sky130_fd_sc_hd__or3b_1 _12981_ (.A(_06134_),
    .B(_06136_),
    .C_N(_06130_),
    .X(_06137_));
 sky130_fd_sc_hd__nand2_1 _12982_ (.A(_06135_),
    .B(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__o2111a_1 _12983_ (.A1(_06125_),
    .A2(_06127_),
    .B1(_06131_),
    .C1(_06129_),
    .D1(_06128_),
    .X(_06139_));
 sky130_fd_sc_hd__a21o_1 _12984_ (.A1(_06117_),
    .A2(_06121_),
    .B1(_06124_),
    .X(_06140_));
 sky130_fd_sc_hd__nand2_1 _12985_ (.A(_06129_),
    .B(_06126_),
    .Y(_06141_));
 sky130_fd_sc_hd__nor2_1 _12986_ (.A(net3876),
    .B(net3085),
    .Y(_06142_));
 sky130_fd_sc_hd__and3_1 _12987_ (.A(net4600),
    .B(net3090),
    .C(_06129_),
    .X(_06143_));
 sky130_fd_sc_hd__a21oi_1 _12988_ (.A1(net3857),
    .A2(net3135),
    .B1(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__o221a_1 _12989_ (.A1(_06140_),
    .A2(_06141_),
    .B1(_06136_),
    .B2(_06142_),
    .C1(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__nor2_1 _12990_ (.A(_06139_),
    .B(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__nand2_1 _12991_ (.A(_06109_),
    .B(_06110_),
    .Y(_06147_));
 sky130_fd_sc_hd__nor2_1 _12992_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06148_));
 sky130_fd_sc_hd__o41a_1 _12993_ (.A1(_06095_),
    .A2(_06104_),
    .A3(_06108_),
    .A4(_06115_),
    .B1(_06118_),
    .X(_06149_));
 sky130_fd_sc_hd__o21a_1 _12994_ (.A1(_06148_),
    .A2(_06149_),
    .B1(_06119_),
    .X(_06150_));
 sky130_fd_sc_hd__xnor2_2 _12995_ (.A(_06147_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__xnor2_2 _12996_ (.A(_06111_),
    .B(_06149_),
    .Y(_06152_));
 sky130_fd_sc_hd__or2_1 _12997_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_06153_));
 sky130_fd_sc_hd__nand2_1 _12998_ (.A(_06153_),
    .B(_06102_),
    .Y(_06154_));
 sky130_fd_sc_hd__a21o_1 _12999_ (.A1(_06098_),
    .A2(_06101_),
    .B1(_06096_),
    .X(_06155_));
 sky130_fd_sc_hd__xnor2_2 _13000_ (.A(_06154_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__nand3_1 _13001_ (.A(_06124_),
    .B(_06117_),
    .C(_06121_),
    .Y(_06157_));
 sky130_fd_sc_hd__and2_1 _13002_ (.A(_06140_),
    .B(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__a21o_1 _13003_ (.A1(_06098_),
    .A2(_06101_),
    .B1(_06103_),
    .X(_06159_));
 sky130_fd_sc_hd__and3_1 _13004_ (.A(_06153_),
    .B(_06159_),
    .C(_06107_),
    .X(_06160_));
 sky130_fd_sc_hd__a21oi_1 _13005_ (.A1(_06153_),
    .A2(_06159_),
    .B1(_06107_),
    .Y(_06161_));
 sky130_fd_sc_hd__nor2_1 _13006_ (.A(_06160_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__xor2_1 _13007_ (.A(_06098_),
    .B(_06101_),
    .X(_06163_));
 sky130_fd_sc_hd__nand2_1 _13008_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_06164_));
 sky130_fd_sc_hd__xnor2_1 _13009_ (.A(_06164_),
    .B(_06099_),
    .Y(_06165_));
 sky130_fd_sc_hd__xor2_1 _13010_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_06166_));
 sky130_fd_sc_hd__or4_1 _13011_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_06165_),
    .D(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__or4_1 _13012_ (.A(_06158_),
    .B(_06162_),
    .C(_06163_),
    .D(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__nor2_1 _13013_ (.A(_06156_),
    .B(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__o31a_1 _13014_ (.A1(_06095_),
    .A2(_06104_),
    .A3(_06108_),
    .B1(_06105_),
    .X(_06170_));
 sky130_fd_sc_hd__xnor2_2 _13015_ (.A(_06115_),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__a21oi_1 _13016_ (.A1(_06122_),
    .A2(_06140_),
    .B1(_06141_),
    .Y(_06172_));
 sky130_fd_sc_hd__and3_1 _13017_ (.A(_06122_),
    .B(_06140_),
    .C(_06141_),
    .X(_06173_));
 sky130_fd_sc_hd__or2_1 _13018_ (.A(_06172_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__and4b_1 _13019_ (.A_N(_06152_),
    .B(_06169_),
    .C(_06171_),
    .D(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__and4bb_1 _13020_ (.A_N(_06138_),
    .B_N(_06146_),
    .C(_06151_),
    .D(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__or2_2 _13021_ (.A(_06133_),
    .B(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__buf_4 _13022_ (.A(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__clkbuf_4 _13023_ (.A(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__xor2_1 _13024_ (.A(net2388),
    .B(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__inv_2 _13025_ (.A(net3034),
    .Y(_06181_));
 sky130_fd_sc_hd__xnor2_1 _13026_ (.A(_06181_),
    .B(_06179_),
    .Y(_06182_));
 sky130_fd_sc_hd__clkbuf_4 _13027_ (.A(net4912),
    .X(_06183_));
 sky130_fd_sc_hd__and2_1 _13028_ (.A(net6185),
    .B(_06178_),
    .X(_06184_));
 sky130_fd_sc_hd__buf_2 _13029_ (.A(net4896),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_4 _13030_ (.A(net6185),
    .X(_06186_));
 sky130_fd_sc_hd__nor2_1 _13031_ (.A(_06186_),
    .B(_06178_),
    .Y(_06187_));
 sky130_fd_sc_hd__nor2_1 _13032_ (.A(net6186),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__and2_1 _13033_ (.A(_06185_),
    .B(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__inv_2 _13034_ (.A(net3804),
    .Y(_06190_));
 sky130_fd_sc_hd__xnor2_1 _13035_ (.A(_06190_),
    .B(_06178_),
    .Y(_06191_));
 sky130_fd_sc_hd__o21a_1 _13036_ (.A1(net6186),
    .A2(_06189_),
    .B1(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__a21o_1 _13037_ (.A1(net3804),
    .A2(_06178_),
    .B1(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__o21a_1 _13038_ (.A1(_06183_),
    .A2(_06179_),
    .B1(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__a21oi_1 _13039_ (.A1(_06183_),
    .A2(_06179_),
    .B1(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__inv_2 _13040_ (.A(net4821),
    .Y(_06196_));
 sky130_fd_sc_hd__xnor2_1 _13041_ (.A(_06196_),
    .B(_06179_),
    .Y(_06197_));
 sky130_fd_sc_hd__and2b_1 _13042_ (.A_N(_06195_),
    .B(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__o21a_1 _13043_ (.A1(net4821),
    .A2(net3034),
    .B1(_06179_),
    .X(_06199_));
 sky130_fd_sc_hd__a21o_1 _13044_ (.A1(_06182_),
    .A2(_06198_),
    .B1(net4822),
    .X(_06200_));
 sky130_fd_sc_hd__or2_1 _13045_ (.A(_06180_),
    .B(net4823),
    .X(_06201_));
 sky130_fd_sc_hd__nand2_1 _13046_ (.A(_06180_),
    .B(net4823),
    .Y(_06202_));
 sky130_fd_sc_hd__or2_1 _13047_ (.A(net3507),
    .B(net4910),
    .X(_06203_));
 sky130_fd_sc_hd__buf_4 _13048_ (.A(net4911),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_8 _13049_ (.A(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__buf_4 _13050_ (.A(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__nor2b_2 _13051_ (.A(net4909),
    .B_N(net6168),
    .Y(_06207_));
 sky130_fd_sc_hd__nand3b_4 _13052_ (.A_N(_04627_),
    .B(_06207_),
    .C(_04626_),
    .Y(_06208_));
 sky130_fd_sc_hd__buf_6 _13053_ (.A(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_8 _13054_ (.A(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_8 _13055_ (.A(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _13056_ (.A(net3983),
    .X(_06212_));
 sky130_fd_sc_hd__inv_2 _13057_ (.A(net3984),
    .Y(_06213_));
 sky130_fd_sc_hd__a22o_1 _13058_ (.A1(net2825),
    .A2(_06213_),
    .B1(net4874),
    .B2(net3620),
    .X(_06214_));
 sky130_fd_sc_hd__a21o_1 _13059_ (.A1(net3620),
    .A2(_04899_),
    .B1(net4874),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_4 _13060_ (.A(net6248),
    .X(_06216_));
 sky130_fd_sc_hd__buf_2 _13061_ (.A(net6251),
    .X(_06217_));
 sky130_fd_sc_hd__nor2_1 _13062_ (.A(net2774),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__inv_2 _13063_ (.A(net6251),
    .Y(_06219_));
 sky130_fd_sc_hd__nor2_1 _13064_ (.A(_04895_),
    .B(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__inv_2 _13065_ (.A(net6248),
    .Y(_06221_));
 sky130_fd_sc_hd__clkbuf_4 _13066_ (.A(net6216),
    .X(_06222_));
 sky130_fd_sc_hd__xnor2_1 _13067_ (.A(net4345),
    .B(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__o221a_1 _13068_ (.A1(net2895),
    .A2(_06221_),
    .B1(_06213_),
    .B2(net2825),
    .C1(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__o221a_1 _13069_ (.A1(_04894_),
    .A2(_06216_),
    .B1(_06218_),
    .B2(_06220_),
    .C1(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__inv_2 _13070_ (.A(net3853),
    .Y(_06226_));
 sky130_fd_sc_hd__inv_2 _13071_ (.A(net4896),
    .Y(_06227_));
 sky130_fd_sc_hd__a2bb2o_1 _13072_ (.A1_N(net3917),
    .A2_N(net4897),
    .B1(_06213_),
    .B2(net4090),
    .X(_06228_));
 sky130_fd_sc_hd__inv_2 _13073_ (.A(net4874),
    .Y(_06229_));
 sky130_fd_sc_hd__a22o_1 _13074_ (.A1(_04823_),
    .A2(net3983),
    .B1(_06181_),
    .B2(net3952),
    .X(_06230_));
 sky130_fd_sc_hd__a221o_1 _13075_ (.A1(net3853),
    .A2(_06229_),
    .B1(_06190_),
    .B2(net4387),
    .C1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__inv_2 _13076_ (.A(net3880),
    .Y(_06232_));
 sky130_fd_sc_hd__a2bb2o_1 _13077_ (.A1_N(net3952),
    .A2_N(_06181_),
    .B1(_06221_),
    .B2(net3995),
    .X(_06233_));
 sky130_fd_sc_hd__a221o_1 _13078_ (.A1(net3881),
    .A2(_06186_),
    .B1(_06196_),
    .B2(net3279),
    .C1(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__a2bb2o_1 _13079_ (.A1_N(net4387),
    .A2_N(_06190_),
    .B1(net4912),
    .B2(_04822_),
    .X(_06235_));
 sky130_fd_sc_hd__a221o_1 _13080_ (.A1(net3996),
    .A2(_06216_),
    .B1(net4821),
    .B2(_04827_),
    .C1(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__or3_1 _13081_ (.A(_06231_),
    .B(_06234_),
    .C(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__a211o_1 _13082_ (.A1(_06226_),
    .A2(net4874),
    .B1(_06228_),
    .C1(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__nand2_1 _13083_ (.A(net3921),
    .B(net6216),
    .Y(_06239_));
 sky130_fd_sc_hd__or2_1 _13084_ (.A(net3921),
    .B(\rbzero.map_rom.f1 ),
    .X(_06240_));
 sky130_fd_sc_hd__or4_1 _13085_ (.A(net2388),
    .B(net2907),
    .C(net1130),
    .D(net1064),
    .X(_06241_));
 sky130_fd_sc_hd__or4_1 _13086_ (.A(net2787),
    .B(net1249),
    .C(net977),
    .D(net2768),
    .X(_06242_));
 sky130_fd_sc_hd__a211o_1 _13087_ (.A1(_06239_),
    .A2(_06240_),
    .B1(_06241_),
    .C1(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__inv_2 _13088_ (.A(_06186_),
    .Y(_06244_));
 sky130_fd_sc_hd__inv_2 _13089_ (.A(net4912),
    .Y(_06245_));
 sky130_fd_sc_hd__a22o_1 _13090_ (.A1(net3917),
    .A2(net4897),
    .B1(net4913),
    .B2(net3893),
    .X(_06246_));
 sky130_fd_sc_hd__a221o_1 _13091_ (.A1(_04837_),
    .A2(_06217_),
    .B1(_06244_),
    .B2(net4675),
    .C1(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__inv_2 _13092_ (.A(net3265),
    .Y(_06248_));
 sky130_fd_sc_hd__a211o_1 _13093_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_06248_),
    .B1(net2611),
    .C1(net2807),
    .X(_06249_));
 sky130_fd_sc_hd__o22a_1 _13094_ (.A1(_04837_),
    .A2(_06217_),
    .B1(_06248_),
    .B2(\rbzero.debug_overlay.playerX[5] ),
    .X(_06250_));
 sky130_fd_sc_hd__or4b_1 _13095_ (.A(_06243_),
    .B(_06247_),
    .C(_06249_),
    .D_N(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__or4_1 _13096_ (.A(net3772),
    .B(net3718),
    .C(net3627),
    .D(net3222),
    .X(_06252_));
 sky130_fd_sc_hd__or4_1 _13097_ (.A(net4524),
    .B(net4581),
    .C(net4783),
    .D(net673),
    .X(_06253_));
 sky130_fd_sc_hd__or4_1 _13098_ (.A(net656),
    .B(net695),
    .C(net692),
    .D(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__or4_1 _13099_ (.A(net4779),
    .B(net3633),
    .C(_06252_),
    .D(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__inv_2 _13100_ (.A(net7770),
    .Y(_06256_));
 sky130_fd_sc_hd__o211a_1 _13101_ (.A1(_06238_),
    .A2(_06251_),
    .B1(_06255_),
    .C1(net4828),
    .X(_06257_));
 sky130_fd_sc_hd__and4b_1 _13102_ (.A_N(_06214_),
    .B(net3621),
    .C(_06225_),
    .D(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__xnor2_1 _13103_ (.A(net2791),
    .B(_06183_),
    .Y(_06259_));
 sky130_fd_sc_hd__o221a_1 _13104_ (.A1(_04886_),
    .A2(_06185_),
    .B1(_06196_),
    .B2(net2726),
    .C1(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__o221a_1 _13105_ (.A1(net2802),
    .A2(net4897),
    .B1(_06244_),
    .B2(net2879),
    .C1(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__or4_1 _13106_ (.A(_06186_),
    .B(net3804),
    .C(_06183_),
    .D(net4821),
    .X(_06262_));
 sky130_fd_sc_hd__nor2_1 _13107_ (.A(_06185_),
    .B(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__xor2_1 _13108_ (.A(net2789),
    .B(net3804),
    .X(_06264_));
 sky130_fd_sc_hd__a221o_1 _13109_ (.A1(net2879),
    .A2(_06244_),
    .B1(_06196_),
    .B2(net2726),
    .C1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__nor2_1 _13110_ (.A(_06263_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__and3_1 _13111_ (.A(_06257_),
    .B(net4898),
    .C(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__nor2_1 _13112_ (.A(net3622),
    .B(net4899),
    .Y(_06268_));
 sky130_fd_sc_hd__inv_2 _13113_ (.A(net4342),
    .Y(_06269_));
 sky130_fd_sc_hd__and2_1 _13114_ (.A(_06269_),
    .B(net4577),
    .X(_06270_));
 sky130_fd_sc_hd__inv_2 _13115_ (.A(net3494),
    .Y(_06271_));
 sky130_fd_sc_hd__inv_2 _13116_ (.A(net3851),
    .Y(_06272_));
 sky130_fd_sc_hd__a22o_1 _13117_ (.A1(_06271_),
    .A2(net3369),
    .B1(_06272_),
    .B2(net3852),
    .X(_06273_));
 sky130_fd_sc_hd__inv_2 _13118_ (.A(net3742),
    .Y(_06274_));
 sky130_fd_sc_hd__o22a_1 _13119_ (.A1(_06269_),
    .A2(net4577),
    .B1(net3780),
    .B2(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__inv_2 _13120_ (.A(net3284),
    .Y(_06276_));
 sky130_fd_sc_hd__inv_2 _13121_ (.A(net3373),
    .Y(_06277_));
 sky130_fd_sc_hd__o22a_1 _13122_ (.A1(net3462),
    .A2(_06276_),
    .B1(net3500),
    .B2(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__inv_2 _13123_ (.A(net3852),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_1 _13124_ (.A(_06271_),
    .B(net3369),
    .Y(_06280_));
 sky130_fd_sc_hd__inv_2 _13125_ (.A(net3240),
    .Y(_06281_));
 sky130_fd_sc_hd__nor2_1 _13126_ (.A(net3447),
    .B(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__inv_2 _13127_ (.A(net3503),
    .Y(_06283_));
 sky130_fd_sc_hd__a2bb2o_1 _13128_ (.A1_N(net3327),
    .A2_N(_06283_),
    .B1(net3447),
    .B2(_06281_),
    .X(_06284_));
 sky130_fd_sc_hd__inv_2 _13129_ (.A(net3566),
    .Y(_06285_));
 sky130_fd_sc_hd__nor2_1 _13130_ (.A(net3542),
    .B(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__inv_2 _13131_ (.A(net3493),
    .Y(_06287_));
 sky130_fd_sc_hd__nor2_1 _13132_ (.A(_06287_),
    .B(net3426),
    .Y(_06288_));
 sky130_fd_sc_hd__and2_1 _13133_ (.A(net3500),
    .B(_06277_),
    .X(_06289_));
 sky130_fd_sc_hd__and2_1 _13134_ (.A(net3780),
    .B(_06274_),
    .X(_06290_));
 sky130_fd_sc_hd__or4_1 _13135_ (.A(_06286_),
    .B(_06288_),
    .C(_06289_),
    .D(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__a22o_1 _13136_ (.A1(_06287_),
    .A2(net3426),
    .B1(net3542),
    .B2(_06285_),
    .X(_06292_));
 sky130_fd_sc_hd__and2_1 _13137_ (.A(net3462),
    .B(_06276_),
    .X(_06293_));
 sky130_fd_sc_hd__a211o_1 _13138_ (.A1(net3327),
    .A2(_06283_),
    .B1(_06292_),
    .C1(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__or4_1 _13139_ (.A(_06282_),
    .B(_06284_),
    .C(_06291_),
    .D(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__a2111oi_1 _13140_ (.A1(net3851),
    .A2(_06279_),
    .B1(_06270_),
    .C1(_06280_),
    .D1(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__and4b_1 _13141_ (.A_N(_06273_),
    .B(_06275_),
    .C(_06278_),
    .D(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__inv_2 _13142_ (.A(net3179),
    .Y(_06298_));
 sky130_fd_sc_hd__inv_2 _13143_ (.A(net3433),
    .Y(_06299_));
 sky130_fd_sc_hd__o22a_1 _13144_ (.A1(net3381),
    .A2(_06298_),
    .B1(net3555),
    .B2(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__inv_2 _13145_ (.A(net3501),
    .Y(_06301_));
 sky130_fd_sc_hd__and2_1 _13146_ (.A(net3381),
    .B(_06298_),
    .X(_06302_));
 sky130_fd_sc_hd__a221oi_1 _13147_ (.A1(net3555),
    .A2(_06299_),
    .B1(net3472),
    .B2(_06301_),
    .C1(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__and2_1 _13148_ (.A(_06300_),
    .B(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__inv_2 _13149_ (.A(net4433),
    .Y(_06305_));
 sky130_fd_sc_hd__a2bb2o_1 _13150_ (.A1_N(net3472),
    .A2_N(_06301_),
    .B1(net3321),
    .B2(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__o21ba_1 _13151_ (.A1(net4483),
    .A2(_06305_),
    .B1_N(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__inv_2 _13152_ (.A(net3047),
    .Y(_06308_));
 sky130_fd_sc_hd__inv_2 _13153_ (.A(net3417),
    .Y(_06309_));
 sky130_fd_sc_hd__o22a_1 _13154_ (.A1(_06308_),
    .A2(net3233),
    .B1(_06309_),
    .B2(net3221),
    .X(_06310_));
 sky130_fd_sc_hd__inv_2 _13155_ (.A(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__inv_2 _13156_ (.A(net3184),
    .Y(_06312_));
 sky130_fd_sc_hd__a2bb2o_1 _13157_ (.A1_N(_06312_),
    .A2_N(net3200),
    .B1(_06309_),
    .B2(net3221),
    .X(_06313_));
 sky130_fd_sc_hd__inv_2 _13158_ (.A(net3578),
    .Y(_06314_));
 sky130_fd_sc_hd__a22o_1 _13159_ (.A1(_06314_),
    .A2(net3174),
    .B1(_06308_),
    .B2(net3233),
    .X(_06315_));
 sky130_fd_sc_hd__inv_2 _13160_ (.A(net3054),
    .Y(_06316_));
 sky130_fd_sc_hd__a2bb2o_1 _13161_ (.A1_N(_06314_),
    .A2_N(net3174),
    .B1(_06316_),
    .B2(net3460),
    .X(_06317_));
 sky130_fd_sc_hd__or4_1 _13162_ (.A(_06311_),
    .B(_06313_),
    .C(_06315_),
    .D(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__inv_2 _13163_ (.A(net3155),
    .Y(_06319_));
 sky130_fd_sc_hd__inv_2 _13164_ (.A(net3432),
    .Y(_06320_));
 sky130_fd_sc_hd__a22o_1 _13165_ (.A1(_06319_),
    .A2(net3209),
    .B1(_06320_),
    .B2(net3554),
    .X(_06321_));
 sky130_fd_sc_hd__nor2_1 _13166_ (.A(_06319_),
    .B(net3209),
    .Y(_06322_));
 sky130_fd_sc_hd__a211o_1 _13167_ (.A1(_06312_),
    .A2(net3795),
    .B1(_06321_),
    .C1(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__inv_2 _13168_ (.A(net3474),
    .Y(_06324_));
 sky130_fd_sc_hd__o22a_1 _13169_ (.A1(_06320_),
    .A2(net3554),
    .B1(_06324_),
    .B2(net3314),
    .X(_06325_));
 sky130_fd_sc_hd__o2bb2a_1 _13170_ (.A1_N(_06324_),
    .A2_N(net3314),
    .B1(_06316_),
    .B2(net3460),
    .X(_06326_));
 sky130_fd_sc_hd__and4bb_1 _13171_ (.A_N(_06318_),
    .B_N(_06323_),
    .C(_06325_),
    .D(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__nor2_1 _13172_ (.A(_06280_),
    .B(_06286_),
    .Y(_06328_));
 sky130_fd_sc_hd__nor2_1 _13173_ (.A(_06282_),
    .B(_06284_),
    .Y(_06329_));
 sky130_fd_sc_hd__o22a_1 _13174_ (.A1(_06272_),
    .A2(net3852),
    .B1(_06282_),
    .B2(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__or2_1 _13175_ (.A(_06273_),
    .B(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__a21oi_1 _13176_ (.A1(_06328_),
    .A2(_06331_),
    .B1(_06292_),
    .Y(_06332_));
 sky130_fd_sc_hd__o31a_1 _13177_ (.A1(_06288_),
    .A2(_06289_),
    .A3(_06332_),
    .B1(_06278_),
    .X(_06333_));
 sky130_fd_sc_hd__nor2_1 _13178_ (.A(_06293_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__a21oi_1 _13179_ (.A1(_06310_),
    .A2(_06313_),
    .B1(_06315_),
    .Y(_06335_));
 sky130_fd_sc_hd__o21ai_1 _13180_ (.A1(_06317_),
    .A2(_06335_),
    .B1(_06326_),
    .Y(_06336_));
 sky130_fd_sc_hd__a21oi_1 _13181_ (.A1(_06325_),
    .A2(_06336_),
    .B1(_06321_),
    .Y(_06337_));
 sky130_fd_sc_hd__o2bb2a_1 _13182_ (.A1_N(_06327_),
    .A2_N(_06334_),
    .B1(_06337_),
    .B2(_06322_),
    .X(_06338_));
 sky130_fd_sc_hd__nand3b_1 _13183_ (.A_N(_06338_),
    .B(_06307_),
    .C(_06304_),
    .Y(_06339_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(_06304_),
    .B(_06306_),
    .Y(_06340_));
 sky130_fd_sc_hd__o211a_1 _13185_ (.A1(_06300_),
    .A2(_06302_),
    .B1(_06339_),
    .C1(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__o21a_1 _13186_ (.A1(_06290_),
    .A2(_06341_),
    .B1(_06275_),
    .X(_06342_));
 sky130_fd_sc_hd__a41o_1 _13187_ (.A1(_06297_),
    .A2(_06304_),
    .A3(_06307_),
    .A4(_06327_),
    .B1(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__or2_2 _13188_ (.A(_06270_),
    .B(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__a22o_1 _13189_ (.A1(_04863_),
    .A2(_06222_),
    .B1(net4913),
    .B2(net2536),
    .X(_06345_));
 sky130_fd_sc_hd__a221o_1 _13190_ (.A1(net2677),
    .A2(_06219_),
    .B1(_06216_),
    .B2(_04860_),
    .C1(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__o22a_1 _13191_ (.A1(net2864),
    .A2(_06190_),
    .B1(net4913),
    .B2(net2536),
    .X(_06347_));
 sky130_fd_sc_hd__o221a_1 _13192_ (.A1(net2905),
    .A2(_06244_),
    .B1(net4821),
    .B2(_04876_),
    .C1(net4914),
    .X(_06348_));
 sky130_fd_sc_hd__o22a_1 _13193_ (.A1(net2677),
    .A2(_06219_),
    .B1(_06196_),
    .B2(net2823),
    .X(_06349_));
 sky130_fd_sc_hd__inv_2 _13194_ (.A(net2925),
    .Y(_06350_));
 sky130_fd_sc_hd__o22a_1 _13195_ (.A1(_04868_),
    .A2(net3984),
    .B1(_06185_),
    .B2(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__a2bb2o_1 _13196_ (.A1_N(net2839),
    .A2_N(_06229_),
    .B1(_06190_),
    .B2(net2864),
    .X(_06352_));
 sky130_fd_sc_hd__a221o_1 _13197_ (.A1(_04868_),
    .A2(net3984),
    .B1(_06185_),
    .B2(_06350_),
    .C1(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__inv_2 _13198_ (.A(_06222_),
    .Y(_06354_));
 sky130_fd_sc_hd__a22o_1 _13199_ (.A1(net2839),
    .A2(_06229_),
    .B1(_06244_),
    .B2(net2905),
    .X(_06355_));
 sky130_fd_sc_hd__a221o_1 _13200_ (.A1(net2705),
    .A2(_06221_),
    .B1(_06354_),
    .B2(net2043),
    .C1(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__nor2_1 _13201_ (.A(_06353_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__and3_1 _13202_ (.A(_06349_),
    .B(_06351_),
    .C(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__nand3b_1 _13203_ (.A_N(_06346_),
    .B(net4915),
    .C(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__a22o_1 _13204_ (.A1(_06216_),
    .A2(_06185_),
    .B1(_06190_),
    .B2(_06219_),
    .X(_06360_));
 sky130_fd_sc_hd__xnor2_1 _13205_ (.A(net3984),
    .B(_06183_),
    .Y(_06361_));
 sky130_fd_sc_hd__a22o_1 _13206_ (.A1(_06222_),
    .A2(_06186_),
    .B1(net3804),
    .B2(_06217_),
    .X(_06362_));
 sky130_fd_sc_hd__a221o_1 _13207_ (.A1(_06221_),
    .A2(net4897),
    .B1(_06244_),
    .B2(_06354_),
    .C1(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__or4_1 _13208_ (.A(_06217_),
    .B(net3984),
    .C(_06185_),
    .D(net3804),
    .X(_06364_));
 sky130_fd_sc_hd__and4_1 _13209_ (.A(_06222_),
    .B(_06186_),
    .C(_06183_),
    .D(_06196_),
    .X(_06365_));
 sky130_fd_sc_hd__or4b_1 _13210_ (.A(_06216_),
    .B(net4874),
    .C(_06364_),
    .D_N(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__o31a_1 _13211_ (.A1(_06360_),
    .A2(_06361_),
    .A3(_06363_),
    .B1(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__and4_1 _13212_ (.A(_06186_),
    .B(net3804),
    .C(_06183_),
    .D(net4821),
    .X(_06368_));
 sky130_fd_sc_hd__and3_1 _13213_ (.A(net3984),
    .B(_06222_),
    .C(net4874),
    .X(_06369_));
 sky130_fd_sc_hd__xnor2_1 _13214_ (.A(net4896),
    .B(_06186_),
    .Y(_06370_));
 sky130_fd_sc_hd__a22o_1 _13215_ (.A1(_06219_),
    .A2(net4897),
    .B1(_06370_),
    .B2(_06216_),
    .X(_06371_));
 sky130_fd_sc_hd__or4_1 _13216_ (.A(_06217_),
    .B(_06216_),
    .C(net3984),
    .D(net4874),
    .X(_06372_));
 sky130_fd_sc_hd__a21o_1 _13217_ (.A1(_06213_),
    .A2(_06190_),
    .B1(_06183_),
    .X(_06373_));
 sky130_fd_sc_hd__a22o_1 _13218_ (.A1(_06219_),
    .A2(net4897),
    .B1(net3804),
    .B2(net3984),
    .X(_06374_));
 sky130_fd_sc_hd__a22o_1 _13219_ (.A1(\rbzero.map_rom.f4 ),
    .A2(net4896),
    .B1(_06186_),
    .B2(_06216_),
    .X(_06375_));
 sky130_fd_sc_hd__a2111o_1 _13220_ (.A1(_06221_),
    .A2(_06244_),
    .B1(_06373_),
    .C1(_06374_),
    .D1(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__a21oi_1 _13221_ (.A1(_06372_),
    .A2(_06376_),
    .B1(_06222_),
    .Y(_06377_));
 sky130_fd_sc_hd__a31o_1 _13222_ (.A1(net3984),
    .A2(net3804),
    .A3(_06371_),
    .B1(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__inv_2 _13223_ (.A(_06364_),
    .Y(_06379_));
 sky130_fd_sc_hd__a311o_1 _13224_ (.A1(_06217_),
    .A2(_06216_),
    .A3(_06369_),
    .B1(_06378_),
    .C1(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__a211oi_1 _13225_ (.A1(_06185_),
    .A2(_06368_),
    .B1(_06380_),
    .C1(_06263_),
    .Y(_06381_));
 sky130_fd_sc_hd__inv_2 _13226_ (.A(_06257_),
    .Y(_06382_));
 sky130_fd_sc_hd__a31o_1 _13227_ (.A1(net4916),
    .A2(_06367_),
    .A3(_06381_),
    .B1(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__nand2_1 _13228_ (.A(net4917),
    .B(net4900),
    .Y(_06384_));
 sky130_fd_sc_hd__or2_1 _13229_ (.A(_06203_),
    .B(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__buf_2 _13230_ (.A(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__or2_1 _13231_ (.A(_06344_),
    .B(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__o21ai_1 _13232_ (.A1(net4911),
    .A2(net4900),
    .B1(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__inv_2 _13233_ (.A(net4917),
    .Y(_06389_));
 sky130_fd_sc_hd__nor2_1 _13234_ (.A(net3507),
    .B(net4910),
    .Y(_06390_));
 sky130_fd_sc_hd__a31o_1 _13235_ (.A1(net4918),
    .A2(net3508),
    .A3(net4900),
    .B1(_04621_),
    .X(_06391_));
 sky130_fd_sc_hd__a211o_2 _13236_ (.A1(_06204_),
    .A2(_06211_),
    .B1(_06388_),
    .C1(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__nor2_2 _13237_ (.A(_06206_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__clkbuf_4 _13238_ (.A(_06392_),
    .X(_06394_));
 sky130_fd_sc_hd__a32o_1 _13239_ (.A1(net4824),
    .A2(_06202_),
    .A3(_06393_),
    .B1(_06394_),
    .B2(net2388),
    .X(_00386_));
 sky130_fd_sc_hd__xor2_1 _13240_ (.A(net5706),
    .B(_06179_),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_4 _13241_ (.A(_06179_),
    .X(_06396_));
 sky130_fd_sc_hd__a21bo_1 _13242_ (.A1(net2388),
    .A2(_06396_),
    .B1_N(_06202_),
    .X(_06397_));
 sky130_fd_sc_hd__xor2_1 _13243_ (.A(_06395_),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a22o_1 _13244_ (.A1(net5706),
    .A2(_06394_),
    .B1(_06393_),
    .B2(_06398_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _13245_ (.A(net4887),
    .B(_06179_),
    .X(_06399_));
 sky130_fd_sc_hd__nor2_1 _13246_ (.A(net4887),
    .B(_06396_),
    .Y(_06400_));
 sky130_fd_sc_hd__nor2_1 _13247_ (.A(_06399_),
    .B(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__and4_1 _13248_ (.A(_06180_),
    .B(_06182_),
    .C(_06198_),
    .D(_06395_),
    .X(_06402_));
 sky130_fd_sc_hd__o21a_1 _13249_ (.A1(net2768),
    .A2(net2388),
    .B1(_06179_),
    .X(_06403_));
 sky130_fd_sc_hd__or3_1 _13250_ (.A(net4822),
    .B(_06402_),
    .C(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__xor2_1 _13251_ (.A(_06401_),
    .B(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__a22o_1 _13252_ (.A1(net4887),
    .A2(_06394_),
    .B1(_06393_),
    .B2(_06405_),
    .X(_00388_));
 sky130_fd_sc_hd__xnor2_1 _13253_ (.A(net5491),
    .B(_06396_),
    .Y(_06406_));
 sky130_fd_sc_hd__a21o_1 _13254_ (.A1(_06401_),
    .A2(_06404_),
    .B1(_06399_),
    .X(_06407_));
 sky130_fd_sc_hd__xnor2_1 _13255_ (.A(_06406_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__a22o_1 _13256_ (.A1(net5491),
    .A2(_06394_),
    .B1(_06393_),
    .B2(_06408_),
    .X(_00389_));
 sky130_fd_sc_hd__o21a_1 _13257_ (.A1(net5491),
    .A2(_06396_),
    .B1(_06407_),
    .X(_06409_));
 sky130_fd_sc_hd__a21oi_1 _13258_ (.A1(net5491),
    .A2(_06396_),
    .B1(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_1 _13259_ (.A(net5510),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__or2_1 _13260_ (.A(_06396_),
    .B(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__nand2_1 _13261_ (.A(_06396_),
    .B(_06411_),
    .Y(_06413_));
 sky130_fd_sc_hd__a32o_1 _13262_ (.A1(_06393_),
    .A2(_06412_),
    .A3(_06413_),
    .B1(_06394_),
    .B2(net5510),
    .X(_00390_));
 sky130_fd_sc_hd__inv_2 _13263_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06414_));
 sky130_fd_sc_hd__mux2_2 _13264_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_06165_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06415_));
 sky130_fd_sc_hd__nand2_1 _13265_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_06416_));
 sky130_fd_sc_hd__xor2_4 _13266_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_06417_));
 sky130_fd_sc_hd__xnor2_2 _13267_ (.A(_06416_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__and2_1 _13268_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .B(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__mux2_4 _13269_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06420_));
 sky130_fd_sc_hd__mux2_4 _13270_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_06420_),
    .S(_06414_),
    .X(_06421_));
 sky130_fd_sc_hd__mux2_4 _13271_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06422_));
 sky130_fd_sc_hd__mux2_4 _13272_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_06422_),
    .S(_06414_),
    .X(_06423_));
 sky130_fd_sc_hd__or2_4 _13273_ (.A(_06421_),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__mux2_1 _13274_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_06166_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06425_));
 sky130_fd_sc_hd__or2_1 _13275_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_06426_));
 sky130_fd_sc_hd__and2_1 _13276_ (.A(_06416_),
    .B(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__mux2_4 _13277_ (.A0(_06425_),
    .A1(_06427_),
    .S(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06428_));
 sky130_fd_sc_hd__a2111oi_4 _13278_ (.A1(_06414_),
    .A2(_06415_),
    .B1(_06419_),
    .C1(_06424_),
    .D1(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__clkbuf_4 _13279_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06430_));
 sky130_fd_sc_hd__buf_2 _13280_ (.A(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__o21ai_1 _13281_ (.A1(_06172_),
    .A2(_06173_),
    .B1(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__clkbuf_4 _13282_ (.A(_06414_),
    .X(_06433_));
 sky130_fd_sc_hd__o21a_1 _13283_ (.A1(net6259),
    .A2(_06430_),
    .B1(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__or2_2 _13284_ (.A(net4561),
    .B(net7146),
    .X(_06435_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(net4561),
    .B(net7146),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _13286_ (.A(_06435_),
    .B(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__nor2_1 _13287_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(net3796),
    .Y(_06438_));
 sky130_fd_sc_hd__and2_1 _13288_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_06439_));
 sky130_fd_sc_hd__a31oi_4 _13289_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A3(_06417_),
    .B1(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_1 _13290_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06441_));
 sky130_fd_sc_hd__nand2_1 _13291_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06442_));
 sky130_fd_sc_hd__o21a_2 _13292_ (.A1(_06440_),
    .A2(_06441_),
    .B1(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__nand2_1 _13293_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(net3796),
    .Y(_06444_));
 sky130_fd_sc_hd__o21ai_4 _13294_ (.A1(_06438_),
    .A2(_06443_),
    .B1(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__and2_1 _13295_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06446_));
 sky130_fd_sc_hd__nor2_1 _13296_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_06447_));
 sky130_fd_sc_hd__nor2_2 _13297_ (.A(_06446_),
    .B(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__nand2_1 _13298_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_06449_));
 sky130_fd_sc_hd__or2_1 _13299_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06450_));
 sky130_fd_sc_hd__and3_1 _13300_ (.A(_06448_),
    .B(_06449_),
    .C(_06450_),
    .X(_06451_));
 sky130_fd_sc_hd__nand2_1 _13301_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_06452_));
 sky130_fd_sc_hd__inv_2 _13302_ (.A(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__nor2_1 _13303_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_06454_));
 sky130_fd_sc_hd__nor2_2 _13304_ (.A(_06453_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__and2_1 _13305_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06456_));
 sky130_fd_sc_hd__nor2_1 _13306_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_06457_));
 sky130_fd_sc_hd__nor2_4 _13307_ (.A(_06456_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__and3_1 _13308_ (.A(_06451_),
    .B(_06455_),
    .C(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__nand2_1 _13309_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_06460_));
 sky130_fd_sc_hd__a21o_1 _13310_ (.A1(_06452_),
    .A2(_06460_),
    .B1(_06454_),
    .X(_06461_));
 sky130_fd_sc_hd__inv_2 _13311_ (.A(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__and2_1 _13312_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06463_));
 sky130_fd_sc_hd__a221o_1 _13313_ (.A1(_06446_),
    .A2(_06450_),
    .B1(_06451_),
    .B2(_06462_),
    .C1(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__a21o_1 _13314_ (.A1(_06445_),
    .A2(_06459_),
    .B1(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__and2_1 _13315_ (.A(net3786),
    .B(net3043),
    .X(_06466_));
 sky130_fd_sc_hd__nor2_1 _13316_ (.A(net3786),
    .B(net3043),
    .Y(_06467_));
 sky130_fd_sc_hd__nor2_1 _13317_ (.A(_06466_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__a21o_1 _13318_ (.A1(_06465_),
    .A2(_06468_),
    .B1(_06466_),
    .X(_06469_));
 sky130_fd_sc_hd__xnor2_2 _13319_ (.A(_06437_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__a22o_1 _13320_ (.A1(_06432_),
    .A2(_06434_),
    .B1(_06470_),
    .B2(net4947),
    .X(_06471_));
 sky130_fd_sc_hd__nand2_2 _13321_ (.A(net4406),
    .B(net6304),
    .Y(_06472_));
 sky130_fd_sc_hd__or2_1 _13322_ (.A(net4406),
    .B(net4787),
    .X(_06473_));
 sky130_fd_sc_hd__a221o_1 _13323_ (.A1(net4561),
    .A2(net7146),
    .B1(_06465_),
    .B2(_06468_),
    .C1(_06466_),
    .X(_06474_));
 sky130_fd_sc_hd__and2_1 _13324_ (.A(net4406),
    .B(net4787),
    .X(_06475_));
 sky130_fd_sc_hd__nor2_1 _13325_ (.A(net4406),
    .B(net6304),
    .Y(_06476_));
 sky130_fd_sc_hd__a311o_1 _13326_ (.A1(_06473_),
    .A2(_06435_),
    .A3(_06474_),
    .B1(_06475_),
    .C1(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__a21oi_2 _13327_ (.A1(_06472_),
    .A2(_06477_),
    .B1(_06433_),
    .Y(_06478_));
 sky130_fd_sc_hd__a311oi_4 _13328_ (.A1(_06094_),
    .A2(_06130_),
    .A3(_06131_),
    .B1(_06132_),
    .C1(net7582),
    .Y(_06479_));
 sky130_fd_sc_hd__nor2_1 _13329_ (.A(net7770),
    .B(_06430_),
    .Y(_06480_));
 sky130_fd_sc_hd__nor3_4 _13330_ (.A(_04635_),
    .B(_06479_),
    .C(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__xnor2_2 _13331_ (.A(_06465_),
    .B(_06468_),
    .Y(_06482_));
 sky130_fd_sc_hd__o21a_1 _13332_ (.A1(net6281),
    .A2(_06430_),
    .B1(_06414_),
    .X(_06483_));
 sky130_fd_sc_hd__a21o_1 _13333_ (.A1(_06140_),
    .A2(_06157_),
    .B1(net7582),
    .X(_06484_));
 sky130_fd_sc_hd__a2bb2o_2 _13334_ (.A1_N(_06433_),
    .A2_N(_06482_),
    .B1(_06483_),
    .B2(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(_06449_),
    .B(_06450_),
    .Y(_06486_));
 sky130_fd_sc_hd__a31oi_4 _13336_ (.A1(_06455_),
    .A2(_06445_),
    .A3(_06458_),
    .B1(_06462_),
    .Y(_06487_));
 sky130_fd_sc_hd__o21bai_1 _13337_ (.A1(_06447_),
    .A2(_06487_),
    .B1_N(_06446_),
    .Y(_06488_));
 sky130_fd_sc_hd__xnor2_2 _13338_ (.A(_06486_),
    .B(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__nor2_1 _13339_ (.A(net6278),
    .B(_06430_),
    .Y(_06490_));
 sky130_fd_sc_hd__a211oi_1 _13340_ (.A1(_06430_),
    .A2(_06151_),
    .B1(_06490_),
    .C1(_04635_),
    .Y(_06491_));
 sky130_fd_sc_hd__xor2_4 _13341_ (.A(_06448_),
    .B(_06487_),
    .X(_06492_));
 sky130_fd_sc_hd__o21a_1 _13342_ (.A1(net6253),
    .A2(_06430_),
    .B1(_06414_),
    .X(_06493_));
 sky130_fd_sc_hd__o21ai_2 _13343_ (.A1(net7582),
    .A2(_06152_),
    .B1(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__o21ai_4 _13344_ (.A1(_06433_),
    .A2(_06492_),
    .B1(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__a21oi_2 _13345_ (.A1(_06445_),
    .A2(_06458_),
    .B1(_06456_),
    .Y(_06496_));
 sky130_fd_sc_hd__xnor2_4 _13346_ (.A(_06455_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__nor2_1 _13347_ (.A(net645),
    .B(_06430_),
    .Y(_06498_));
 sky130_fd_sc_hd__a211oi_2 _13348_ (.A1(_06430_),
    .A2(_06171_),
    .B1(_06498_),
    .C1(_04635_),
    .Y(_06499_));
 sky130_fd_sc_hd__xnor2_4 _13349_ (.A(_06445_),
    .B(_06458_),
    .Y(_06500_));
 sky130_fd_sc_hd__a21oi_1 _13350_ (.A1(net3262),
    .A2(net7582),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06501_));
 sky130_fd_sc_hd__o31a_1 _13351_ (.A1(net7582),
    .A2(_06160_),
    .A3(_06161_),
    .B1(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__a21oi_4 _13352_ (.A1(_04635_),
    .A2(_06500_),
    .B1(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__or2_1 _13353_ (.A(net3356),
    .B(_06430_),
    .X(_06504_));
 sky130_fd_sc_hd__o21ai_4 _13354_ (.A1(net7582),
    .A2(_06156_),
    .B1(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__and2b_1 _13355_ (.A_N(_06438_),
    .B(_06444_),
    .X(_06506_));
 sky130_fd_sc_hd__xnor2_2 _13356_ (.A(_06443_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__nand2_2 _13357_ (.A(_04635_),
    .B(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__and2b_1 _13358_ (.A_N(_06441_),
    .B(_06442_),
    .X(_06509_));
 sky130_fd_sc_hd__xnor2_2 _13359_ (.A(_06440_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__or2_1 _13360_ (.A(_06414_),
    .B(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__and2_1 _13361_ (.A(net3206),
    .B(net7582),
    .X(_06512_));
 sky130_fd_sc_hd__a211o_1 _13362_ (.A1(\rbzero.wall_tracer.rcp_sel[2] ),
    .A2(_06163_),
    .B1(_06512_),
    .C1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06513_));
 sky130_fd_sc_hd__a21boi_4 _13363_ (.A1(_06511_),
    .A2(_06513_),
    .B1_N(_06429_),
    .Y(_06514_));
 sky130_fd_sc_hd__o211ai_4 _13364_ (.A1(_04635_),
    .A2(_06505_),
    .B1(_06508_),
    .C1(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__a2111o_1 _13365_ (.A1(_04635_),
    .A2(_06497_),
    .B1(_06499_),
    .C1(_06503_),
    .D1(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__a2111o_4 _13366_ (.A1(_04635_),
    .A2(_06489_),
    .B1(_06491_),
    .C1(_06495_),
    .D1(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__o22a_1 _13367_ (.A1(_06478_),
    .A2(net82),
    .B1(_06485_),
    .B2(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__xor2_2 _13368_ (.A(_06471_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__nor2_1 _13369_ (.A(net4406),
    .B(net4787),
    .Y(_06520_));
 sky130_fd_sc_hd__nor2_1 _13370_ (.A(_06520_),
    .B(_06475_),
    .Y(_06521_));
 sky130_fd_sc_hd__inv_2 _13371_ (.A(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__nand3_1 _13372_ (.A(_06435_),
    .B(_06474_),
    .C(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__a21o_1 _13373_ (.A1(_06435_),
    .A2(_06474_),
    .B1(_06522_),
    .X(_06524_));
 sky130_fd_sc_hd__a21oi_1 _13374_ (.A1(net7552),
    .A2(net7582),
    .B1(_04635_),
    .Y(_06525_));
 sky130_fd_sc_hd__o31a_1 _13375_ (.A1(net7582),
    .A2(_06139_),
    .A3(_06145_),
    .B1(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__a31o_2 _13376_ (.A1(net4947),
    .A2(_06523_),
    .A3(_06524_),
    .B1(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__a221o_1 _13377_ (.A1(_06432_),
    .A2(_06434_),
    .B1(_06470_),
    .B2(net4947),
    .C1(_06485_),
    .X(_06528_));
 sky130_fd_sc_hd__o22a_1 _13378_ (.A1(_06478_),
    .A2(net82),
    .B1(_06517_),
    .B2(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__xor2_2 _13379_ (.A(_06527_),
    .B(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__or2b_4 _13380_ (.A(_06519_),
    .B_N(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__a31o_1 _13381_ (.A1(_06473_),
    .A2(_06435_),
    .A3(_06474_),
    .B1(_06475_),
    .X(_06532_));
 sky130_fd_sc_hd__inv_2 _13382_ (.A(_06472_),
    .Y(_06533_));
 sky130_fd_sc_hd__nor2_1 _13383_ (.A(_06533_),
    .B(_06476_),
    .Y(_06534_));
 sky130_fd_sc_hd__xnor2_2 _13384_ (.A(_06532_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__nor2_1 _13385_ (.A(net7476),
    .B(_06431_),
    .Y(_06536_));
 sky130_fd_sc_hd__a311o_1 _13386_ (.A1(_06431_),
    .A2(_06135_),
    .A3(_06137_),
    .B1(_06536_),
    .C1(net4947),
    .X(_06537_));
 sky130_fd_sc_hd__o21a_1 _13387_ (.A1(_06433_),
    .A2(_06535_),
    .B1(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__nor2_2 _13388_ (.A(_06517_),
    .B(_06528_),
    .Y(_06539_));
 sky130_fd_sc_hd__clkbuf_8 _13389_ (.A(_06478_),
    .X(_06540_));
 sky130_fd_sc_hd__nor2_4 _13390_ (.A(_06540_),
    .B(_06481_),
    .Y(_06541_));
 sky130_fd_sc_hd__a21oi_1 _13391_ (.A1(_06527_),
    .A2(_06539_),
    .B1(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__xnor2_2 _13392_ (.A(_06538_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__or2_4 _13393_ (.A(_06531_),
    .B(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__nor2_4 _13394_ (.A(net4947),
    .B(_06479_),
    .Y(_06545_));
 sky130_fd_sc_hd__or2_1 _13395_ (.A(net6098),
    .B(_06431_),
    .X(_06546_));
 sky130_fd_sc_hd__a21oi_4 _13396_ (.A1(_06545_),
    .A2(_06546_),
    .B1(_06540_),
    .Y(_06547_));
 sky130_fd_sc_hd__or2_1 _13397_ (.A(net6123),
    .B(_06431_),
    .X(_06548_));
 sky130_fd_sc_hd__a21oi_4 _13398_ (.A1(_06545_),
    .A2(_06548_),
    .B1(_06540_),
    .Y(_06549_));
 sky130_fd_sc_hd__o211a_1 _13399_ (.A1(_06433_),
    .A2(_06535_),
    .B1(_06527_),
    .C1(_06537_),
    .X(_06550_));
 sky130_fd_sc_hd__a31o_1 _13400_ (.A1(_06549_),
    .A2(_06539_),
    .A3(_06550_),
    .B1(_06541_),
    .X(_06551_));
 sky130_fd_sc_hd__xor2_4 _13401_ (.A(_06547_),
    .B(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__a21oi_2 _13402_ (.A1(_06539_),
    .A2(_06550_),
    .B1(_06541_),
    .Y(_06553_));
 sky130_fd_sc_hd__xnor2_2 _13403_ (.A(_06549_),
    .B(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__o21ai_2 _13404_ (.A1(_06540_),
    .A2(net82),
    .B1(_06517_),
    .Y(_06555_));
 sky130_fd_sc_hd__xnor2_2 _13405_ (.A(_06485_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__or4_4 _13406_ (.A(_06544_),
    .B(_06552_),
    .C(_06554_),
    .D(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__or2_1 _13407_ (.A(net6150),
    .B(_06431_),
    .X(_06558_));
 sky130_fd_sc_hd__a21o_1 _13408_ (.A1(_06545_),
    .A2(_06558_),
    .B1(_06540_),
    .X(_06559_));
 sky130_fd_sc_hd__a21o_2 _13409_ (.A1(_06472_),
    .A2(_06477_),
    .B1(_06433_),
    .X(_06560_));
 sky130_fd_sc_hd__a41o_2 _13410_ (.A1(_06547_),
    .A2(_06549_),
    .A3(_06539_),
    .A4(_06550_),
    .B1(_06541_),
    .X(_06561_));
 sky130_fd_sc_hd__o21ai_1 _13411_ (.A1(net6148),
    .A2(_06431_),
    .B1(_06545_),
    .Y(_06562_));
 sky130_fd_sc_hd__a31o_1 _13412_ (.A1(_06560_),
    .A2(_06561_),
    .A3(_06562_),
    .B1(_06541_),
    .X(_06563_));
 sky130_fd_sc_hd__xor2_1 _13413_ (.A(_06559_),
    .B(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__buf_2 _13414_ (.A(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__nand2_1 _13415_ (.A(_06560_),
    .B(_06562_),
    .Y(_06566_));
 sky130_fd_sc_hd__xor2_1 _13416_ (.A(_06561_),
    .B(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__nor2_1 _13417_ (.A(net7440),
    .B(_06431_),
    .Y(_06568_));
 sky130_fd_sc_hd__o21a_1 _13418_ (.A1(_06479_),
    .A2(_06568_),
    .B1(_06433_),
    .X(_06569_));
 sky130_fd_sc_hd__nand2_1 _13419_ (.A(_06472_),
    .B(_06477_),
    .Y(_06570_));
 sky130_fd_sc_hd__o21ba_1 _13420_ (.A1(_06433_),
    .A2(_06570_),
    .B1_N(_06569_),
    .X(_06571_));
 sky130_fd_sc_hd__and4_1 _13421_ (.A(_06547_),
    .B(_06549_),
    .C(_06539_),
    .D(_06550_),
    .X(_06572_));
 sky130_fd_sc_hd__and2b_1 _13422_ (.A_N(_06559_),
    .B(_06562_),
    .X(_06573_));
 sky130_fd_sc_hd__or2_1 _13423_ (.A(net6146),
    .B(_06431_),
    .X(_06574_));
 sky130_fd_sc_hd__a21o_1 _13424_ (.A1(_06545_),
    .A2(_06574_),
    .B1(_06540_),
    .X(_06575_));
 sky130_fd_sc_hd__inv_2 _13425_ (.A(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__o21ai_1 _13426_ (.A1(net7442),
    .A2(_06431_),
    .B1(_06545_),
    .Y(_06577_));
 sky130_fd_sc_hd__a41o_1 _13427_ (.A1(_06572_),
    .A2(_06573_),
    .A3(_06576_),
    .A4(_06577_),
    .B1(_06541_),
    .X(_06578_));
 sky130_fd_sc_hd__mux2_1 _13428_ (.A0(_06569_),
    .A1(_06571_),
    .S(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__and4_1 _13429_ (.A(_06572_),
    .B(_06573_),
    .C(_06576_),
    .D(_06577_),
    .X(_06580_));
 sky130_fd_sc_hd__nand3_1 _13430_ (.A(_06481_),
    .B(_06568_),
    .C(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand2_1 _13431_ (.A(_06560_),
    .B(_06577_),
    .Y(_06582_));
 sky130_fd_sc_hd__a31o_1 _13432_ (.A1(_06572_),
    .A2(_06573_),
    .A3(_06576_),
    .B1(_06541_),
    .X(_06583_));
 sky130_fd_sc_hd__xor2_2 _13433_ (.A(_06582_),
    .B(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__o21a_1 _13434_ (.A1(_06541_),
    .A2(_06573_),
    .B1(_06561_),
    .X(_06585_));
 sky130_fd_sc_hd__xnor2_2 _13435_ (.A(_06576_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__and4b_2 _13436_ (.A_N(_06579_),
    .B(_06581_),
    .C(_06584_),
    .D(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__and4b_2 _13437_ (.A_N(_06557_),
    .B(_06565_),
    .C(_06567_),
    .D(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__buf_4 _13438_ (.A(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__o21ai_2 _13439_ (.A1(_06540_),
    .A2(net82),
    .B1(_06516_),
    .Y(_06590_));
 sky130_fd_sc_hd__xnor2_4 _13440_ (.A(_06495_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__a21o_1 _13441_ (.A1(net4947),
    .A2(_06489_),
    .B1(_06491_),
    .X(_06592_));
 sky130_fd_sc_hd__or3_2 _13442_ (.A(net4947),
    .B(_06479_),
    .C(_06480_),
    .X(_06593_));
 sky130_fd_sc_hd__a2bb2o_2 _13443_ (.A1_N(_06516_),
    .A2_N(_06495_),
    .B1(_06560_),
    .B2(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__xnor2_4 _13444_ (.A(_06592_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__or2_1 _13445_ (.A(_06591_),
    .B(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__inv_2 _13446_ (.A(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__a21o_1 _13447_ (.A1(net4947),
    .A2(_06497_),
    .B1(_06499_),
    .X(_06598_));
 sky130_fd_sc_hd__a2bb2o_2 _13448_ (.A1_N(_06515_),
    .A2_N(_06503_),
    .B1(_06560_),
    .B2(_06593_),
    .X(_06599_));
 sky130_fd_sc_hd__xnor2_4 _13449_ (.A(_06598_),
    .B(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__o21ai_4 _13450_ (.A1(net4947),
    .A2(_06505_),
    .B1(_06508_),
    .Y(_06601_));
 sky130_fd_sc_hd__a21o_1 _13451_ (.A1(_06560_),
    .A2(_06593_),
    .B1(_06514_),
    .X(_06602_));
 sky130_fd_sc_hd__xnor2_2 _13452_ (.A(_06601_),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__nand2_2 _13453_ (.A(_06511_),
    .B(_06513_),
    .Y(_06604_));
 sky130_fd_sc_hd__a21o_1 _13454_ (.A1(_06560_),
    .A2(_06593_),
    .B1(_06429_),
    .X(_06605_));
 sky130_fd_sc_hd__xnor2_4 _13455_ (.A(_06604_),
    .B(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__o21ai_4 _13456_ (.A1(_06540_),
    .A2(net82),
    .B1(_06515_),
    .Y(_06607_));
 sky130_fd_sc_hd__xor2_2 _13457_ (.A(_06503_),
    .B(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__or4bb_2 _13458_ (.A(_06600_),
    .B(_06603_),
    .C_N(_06606_),
    .D_N(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__inv_2 _13459_ (.A(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__nand4_4 _13460_ (.A(net84),
    .B(_06589_),
    .C(_06597_),
    .D(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__xnor2_2 _13461_ (.A(_06561_),
    .B(_06566_),
    .Y(_06612_));
 sky130_fd_sc_hd__or4bb_4 _13462_ (.A(_06612_),
    .B(_06557_),
    .C_N(_06564_),
    .D_N(_06587_),
    .X(_06613_));
 sky130_fd_sc_hd__inv_2 _13463_ (.A(_06421_),
    .Y(_06614_));
 sky130_fd_sc_hd__or2_2 _13464_ (.A(_06614_),
    .B(_06541_),
    .X(_06615_));
 sky130_fd_sc_hd__xnor2_4 _13465_ (.A(_06423_),
    .B(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__a21o_2 _13466_ (.A1(_06433_),
    .A2(_06415_),
    .B1(_06419_),
    .X(_06617_));
 sky130_fd_sc_hd__o22a_2 _13467_ (.A1(_06424_),
    .A2(_06428_),
    .B1(_06540_),
    .B2(net82),
    .X(_06618_));
 sky130_fd_sc_hd__xnor2_4 _13468_ (.A(_06617_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__o21a_2 _13469_ (.A1(_06540_),
    .A2(net82),
    .B1(_06424_),
    .X(_06620_));
 sky130_fd_sc_hd__xnor2_2 _13470_ (.A(_06428_),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand2_1 _13471_ (.A(_06619_),
    .B(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__or3_1 _13472_ (.A(_06614_),
    .B(_06616_),
    .C(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__or4_4 _13473_ (.A(_06613_),
    .B(_06596_),
    .C(_06609_),
    .D(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__and2_2 _13474_ (.A(net3538),
    .B(net3237),
    .X(_06625_));
 sky130_fd_sc_hd__nand2_4 _13475_ (.A(net7757),
    .B(net3237),
    .Y(_06626_));
 sky130_fd_sc_hd__xnor2_2 _13476_ (.A(_06503_),
    .B(_06607_),
    .Y(_06627_));
 sky130_fd_sc_hd__and4b_2 _13477_ (.A_N(_06600_),
    .B(_06597_),
    .C(_06588_),
    .D(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__nor2_1 _13478_ (.A(_06612_),
    .B(_06552_),
    .Y(_06629_));
 sky130_fd_sc_hd__and4_1 _13479_ (.A(_06565_),
    .B(_06587_),
    .C(_06554_),
    .D(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__inv_2 _13480_ (.A(_06543_),
    .Y(_06631_));
 sky130_fd_sc_hd__xor2_2 _13481_ (.A(_06549_),
    .B(_06553_),
    .X(_06632_));
 sky130_fd_sc_hd__and3_1 _13482_ (.A(_06631_),
    .B(_06632_),
    .C(_06629_),
    .X(_06633_));
 sky130_fd_sc_hd__nor2_1 _13483_ (.A(_06591_),
    .B(_06609_),
    .Y(_06634_));
 sky130_fd_sc_hd__or2_1 _13484_ (.A(_06556_),
    .B(_06595_),
    .X(_06635_));
 sky130_fd_sc_hd__nor2_1 _13485_ (.A(_06531_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__and4b_1 _13486_ (.A_N(_06622_),
    .B(_06634_),
    .C(_06636_),
    .D(_06616_),
    .X(_06637_));
 sky130_fd_sc_hd__inv_2 _13487_ (.A(_06591_),
    .Y(_06638_));
 sky130_fd_sc_hd__nor4_1 _13488_ (.A(_06531_),
    .B(_06543_),
    .C(_06554_),
    .D(_06635_),
    .Y(_06639_));
 sky130_fd_sc_hd__and3_1 _13489_ (.A(_06638_),
    .B(_06600_),
    .C(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__or2_1 _13490_ (.A(_06612_),
    .B(_06552_),
    .X(_06641_));
 sky130_fd_sc_hd__a211oi_1 _13491_ (.A1(_06633_),
    .A2(_06637_),
    .B1(_06640_),
    .C1(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__a21boi_1 _13492_ (.A1(_06565_),
    .A2(_06642_),
    .B1_N(_06587_),
    .Y(_06643_));
 sky130_fd_sc_hd__nor2_1 _13493_ (.A(_06638_),
    .B(_06595_),
    .Y(_06644_));
 sky130_fd_sc_hd__xor2_1 _13494_ (.A(_06485_),
    .B(_06555_),
    .X(_06645_));
 sky130_fd_sc_hd__and3b_1 _13495_ (.A_N(_06531_),
    .B(_06645_),
    .C(_06595_),
    .X(_06646_));
 sky130_fd_sc_hd__and4_1 _13496_ (.A(_06565_),
    .B(_06587_),
    .C(_06633_),
    .D(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__a21oi_1 _13497_ (.A1(_06589_),
    .A2(_06644_),
    .B1(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__or4b_2 _13498_ (.A(_06628_),
    .B(_06630_),
    .C(_06643_),
    .D_N(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__and4_1 _13499_ (.A(_06565_),
    .B(_06587_),
    .C(_06632_),
    .D(_06629_),
    .X(_06650_));
 sky130_fd_sc_hd__and2_1 _13500_ (.A(_06544_),
    .B(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__and3_1 _13501_ (.A(_06565_),
    .B(_06587_),
    .C(_06629_),
    .X(_06652_));
 sky130_fd_sc_hd__or2_1 _13502_ (.A(_06544_),
    .B(_06645_),
    .X(_06653_));
 sky130_fd_sc_hd__inv_2 _13503_ (.A(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__a22o_1 _13504_ (.A1(_06652_),
    .A2(_06640_),
    .B1(_06650_),
    .B2(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__or4b_2 _13505_ (.A(_06628_),
    .B(_06651_),
    .C(_06655_),
    .D_N(_06648_),
    .X(_06656_));
 sky130_fd_sc_hd__or3_4 _13506_ (.A(_06626_),
    .B(_06649_),
    .C(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__o21ai_2 _13507_ (.A1(_06626_),
    .A2(_06649_),
    .B1(_06656_),
    .Y(_06658_));
 sky130_fd_sc_hd__nand2_2 _13508_ (.A(_06657_),
    .B(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__clkbuf_2 _13509_ (.A(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__nor2_2 _13510_ (.A(_06626_),
    .B(_06649_),
    .Y(_06661_));
 sky130_fd_sc_hd__buf_2 _13511_ (.A(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_2 _13512_ (.A(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__buf_2 _13513_ (.A(net7843),
    .X(_06664_));
 sky130_fd_sc_hd__and3_1 _13514_ (.A(_06588_),
    .B(_06597_),
    .C(_06610_),
    .X(_06665_));
 sky130_fd_sc_hd__xor2_4 _13515_ (.A(_06428_),
    .B(_06620_),
    .X(_06666_));
 sky130_fd_sc_hd__a31o_4 _13516_ (.A1(_06665_),
    .A2(_06619_),
    .A3(_06666_),
    .B1(_06628_),
    .X(_06667_));
 sky130_fd_sc_hd__and4_4 _13517_ (.A(net84),
    .B(_06588_),
    .C(_06597_),
    .D(_06610_),
    .X(_06668_));
 sky130_fd_sc_hd__inv_2 _13518_ (.A(_06619_),
    .Y(_06669_));
 sky130_fd_sc_hd__and4_1 _13519_ (.A(_06519_),
    .B(_06530_),
    .C(_06631_),
    .D(_06632_),
    .X(_06670_));
 sky130_fd_sc_hd__a311o_1 _13520_ (.A1(_06669_),
    .A2(_06634_),
    .A3(_06639_),
    .B1(_06670_),
    .C1(_06552_),
    .X(_06671_));
 sky130_fd_sc_hd__nand2_1 _13521_ (.A(_06584_),
    .B(_06586_),
    .Y(_06672_));
 sky130_fd_sc_hd__and3b_1 _13522_ (.A_N(_06579_),
    .B(_06581_),
    .C(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__a41o_1 _13523_ (.A1(_06567_),
    .A2(_06565_),
    .A3(_06587_),
    .A4(_06671_),
    .B1(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__or4_2 _13524_ (.A(_06668_),
    .B(_06630_),
    .C(_06655_),
    .D(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__nor2_4 _13525_ (.A(_06667_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__clkbuf_4 _13526_ (.A(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__clkbuf_4 _13527_ (.A(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__and4bb_1 _13528_ (.A_N(_06579_),
    .B_N(_06586_),
    .C(_06581_),
    .D(_06584_),
    .X(_06679_));
 sky130_fd_sc_hd__a311o_1 _13529_ (.A1(_06612_),
    .A2(_06565_),
    .A3(_06587_),
    .B1(_06679_),
    .C1(_06579_),
    .X(_06680_));
 sky130_fd_sc_hd__a211o_1 _13530_ (.A1(_06588_),
    .A2(_06644_),
    .B1(_06630_),
    .C1(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__nor2_1 _13531_ (.A(_06530_),
    .B(_06543_),
    .Y(_06682_));
 sky130_fd_sc_hd__o21ai_2 _13532_ (.A1(_06654_),
    .A2(_06682_),
    .B1(_06650_),
    .Y(_06683_));
 sky130_fd_sc_hd__or4_1 _13533_ (.A(_06606_),
    .B(_06627_),
    .C(_06600_),
    .D(_06603_),
    .X(_06684_));
 sky130_fd_sc_hd__or3_4 _13534_ (.A(_06613_),
    .B(_06596_),
    .C(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__nand4b_4 _13535_ (.A_N(_06681_),
    .B(_06683_),
    .C(_06624_),
    .D(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__nor2_8 _13536_ (.A(_06667_),
    .B(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__clkbuf_4 _13537_ (.A(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__buf_1 _13538_ (.A(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__clkbuf_4 _13539_ (.A(net7908),
    .X(_06690_));
 sky130_fd_sc_hd__or2_1 _13540_ (.A(_06667_),
    .B(_06675_),
    .X(_06691_));
 sky130_fd_sc_hd__clkbuf_4 _13541_ (.A(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__a31oi_4 _13542_ (.A1(_06665_),
    .A2(_06619_),
    .A3(_06666_),
    .B1(_06628_),
    .Y(_06693_));
 sky130_fd_sc_hd__and4b_2 _13543_ (.A_N(_06681_),
    .B(_06683_),
    .C(_06624_),
    .D(_06685_),
    .X(_06694_));
 sky130_fd_sc_hd__nand2_4 _13544_ (.A(_06694_),
    .B(_06693_),
    .Y(_06695_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(_06556_),
    .A1(_06595_),
    .S(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__buf_2 _13546_ (.A(_06693_),
    .X(_06697_));
 sky130_fd_sc_hd__buf_4 _13547_ (.A(_06694_),
    .X(_06698_));
 sky130_fd_sc_hd__a21oi_1 _13548_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06519_),
    .Y(_06699_));
 sky130_fd_sc_hd__a211oi_1 _13549_ (.A1(net538),
    .A2(_06687_),
    .B1(_06699_),
    .C1(_06692_),
    .Y(_06700_));
 sky130_fd_sc_hd__a21oi_1 _13550_ (.A1(_06692_),
    .A2(_06696_),
    .B1(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand2_1 _13551_ (.A(_06663_),
    .B(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__mux2_1 _13552_ (.A0(_06612_),
    .A1(_06552_),
    .S(_06695_),
    .X(_06703_));
 sky130_fd_sc_hd__mux2_1 _13553_ (.A0(_06543_),
    .A1(_06554_),
    .S(_06687_),
    .X(_06704_));
 sky130_fd_sc_hd__mux2_1 _13554_ (.A0(_06703_),
    .A1(_06704_),
    .S(_06692_),
    .X(_06705_));
 sky130_fd_sc_hd__or2_1 _13555_ (.A(_06663_),
    .B(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__clkbuf_4 _13556_ (.A(_06692_),
    .X(_06707_));
 sky130_fd_sc_hd__mux2_1 _13557_ (.A0(_06565_),
    .A1(_06586_),
    .S(_06689_),
    .X(_06708_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(_06584_),
    .B(_06678_),
    .Y(_06709_));
 sky130_fd_sc_hd__a21boi_1 _13559_ (.A1(_06707_),
    .A2(_06708_),
    .B1_N(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__a31o_1 _13560_ (.A1(_06657_),
    .A2(_06702_),
    .A3(_06706_),
    .B1(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__nand2_1 _13561_ (.A(_06650_),
    .B(_06654_),
    .Y(_06712_));
 sky130_fd_sc_hd__a21o_2 _13562_ (.A1(_06675_),
    .A2(_06686_),
    .B1(_06667_),
    .X(_06713_));
 sky130_fd_sc_hd__a22o_2 _13563_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06713_),
    .B2(_06661_),
    .X(_06714_));
 sky130_fd_sc_hd__nand2_2 _13564_ (.A(net7431),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__nand2_2 _13565_ (.A(_06589_),
    .B(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__xnor2_4 _13566_ (.A(_06676_),
    .B(_06687_),
    .Y(_06717_));
 sky130_fd_sc_hd__a21oi_1 _13567_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06600_),
    .Y(_06718_));
 sky130_fd_sc_hd__a21oi_1 _13568_ (.A1(_06608_),
    .A2(_06688_),
    .B1(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__nor2_1 _13569_ (.A(_06717_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__xnor2_2 _13570_ (.A(_06707_),
    .B(_06688_),
    .Y(_06721_));
 sky130_fd_sc_hd__buf_2 _13571_ (.A(_06695_),
    .X(_06722_));
 sky130_fd_sc_hd__mux2_1 _13572_ (.A0(_06591_),
    .A1(_06595_),
    .S(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__xnor2_2 _13573_ (.A(_06661_),
    .B(_06713_),
    .Y(_06724_));
 sky130_fd_sc_hd__clkbuf_2 _13574_ (.A(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__o21ai_1 _13575_ (.A1(_06721_),
    .A2(_06723_),
    .B1(_06725_),
    .Y(_06726_));
 sky130_fd_sc_hd__xor2_2 _13576_ (.A(_06601_),
    .B(_06602_),
    .X(_06727_));
 sky130_fd_sc_hd__mux4_2 _13577_ (.A0(_06606_),
    .A1(_06619_),
    .A2(_06621_),
    .A3(_06727_),
    .S0(_06722_),
    .S1(_06692_),
    .X(_06728_));
 sky130_fd_sc_hd__o22a_1 _13578_ (.A1(_06720_),
    .A2(_06726_),
    .B1(_06728_),
    .B2(_06725_),
    .X(_06729_));
 sky130_fd_sc_hd__a21o_1 _13579_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06616_),
    .X(_06730_));
 sky130_fd_sc_hd__o21a_1 _13580_ (.A1(_06421_),
    .A2(_06695_),
    .B1(_06730_),
    .X(_06731_));
 sky130_fd_sc_hd__and3_1 _13581_ (.A(_06724_),
    .B(_06717_),
    .C(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__buf_4 _13582_ (.A(_06613_),
    .X(_06733_));
 sky130_fd_sc_hd__nor2_2 _13583_ (.A(net7433),
    .B(_06715_),
    .Y(_06734_));
 sky130_fd_sc_hd__a2bb2o_1 _13584_ (.A1_N(_06716_),
    .A2_N(_06729_),
    .B1(_06732_),
    .B2(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__nor2_4 _13585_ (.A(_06711_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__buf_4 _13586_ (.A(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__inv_2 _13587_ (.A(_06552_),
    .Y(_06738_));
 sky130_fd_sc_hd__mux2_4 _13588_ (.A0(_06738_),
    .A1(_06632_),
    .S(_06695_),
    .X(_06739_));
 sky130_fd_sc_hd__mux2_1 _13589_ (.A0(_06530_),
    .A1(_06631_),
    .S(_06687_),
    .X(_06740_));
 sky130_fd_sc_hd__mux2_2 _13590_ (.A0(_06739_),
    .A1(_06740_),
    .S(_06692_),
    .X(_06741_));
 sky130_fd_sc_hd__or2_1 _13591_ (.A(_06626_),
    .B(_06649_),
    .X(_06742_));
 sky130_fd_sc_hd__buf_2 _13592_ (.A(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__or3_1 _13593_ (.A(_06519_),
    .B(_06667_),
    .C(_06686_),
    .X(_06744_));
 sky130_fd_sc_hd__a21o_1 _13594_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06556_),
    .X(_06745_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(_06744_),
    .A2(_06745_),
    .B1(_06692_),
    .Y(_06746_));
 sky130_fd_sc_hd__a21o_1 _13596_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06591_),
    .X(_06747_));
 sky130_fd_sc_hd__or3_1 _13597_ (.A(_06595_),
    .B(_06667_),
    .C(_06686_),
    .X(_06748_));
 sky130_fd_sc_hd__a21oi_1 _13598_ (.A1(_06747_),
    .A2(_06748_),
    .B1(_06676_),
    .Y(_06749_));
 sky130_fd_sc_hd__or3_1 _13599_ (.A(_06743_),
    .B(_06746_),
    .C(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__o21a_1 _13600_ (.A1(_06662_),
    .A2(_06741_),
    .B1(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__nor2_1 _13601_ (.A(_06743_),
    .B(_06656_),
    .Y(_06752_));
 sky130_fd_sc_hd__a21oi_2 _13602_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06603_),
    .Y(_06753_));
 sky130_fd_sc_hd__a211o_1 _13603_ (.A1(_06608_),
    .A2(_06687_),
    .B1(_06753_),
    .C1(_06676_),
    .X(_06754_));
 sky130_fd_sc_hd__a211o_1 _13604_ (.A1(_06638_),
    .A2(_06687_),
    .B1(_06718_),
    .C1(_06691_),
    .X(_06755_));
 sky130_fd_sc_hd__a21o_1 _13605_ (.A1(_06754_),
    .A2(_06755_),
    .B1(_06661_),
    .X(_06756_));
 sky130_fd_sc_hd__or3_1 _13606_ (.A(_06666_),
    .B(_06628_),
    .C(_06686_),
    .X(_06757_));
 sky130_fd_sc_hd__a21oi_1 _13607_ (.A1(_06730_),
    .A2(_06757_),
    .B1(_06676_),
    .Y(_06758_));
 sky130_fd_sc_hd__and3_1 _13608_ (.A(_06606_),
    .B(_06693_),
    .C(_06694_),
    .X(_06759_));
 sky130_fd_sc_hd__a21oi_1 _13609_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06669_),
    .Y(_06760_));
 sky130_fd_sc_hd__o21a_1 _13610_ (.A1(_06759_),
    .A2(_06760_),
    .B1(_06676_),
    .X(_06761_));
 sky130_fd_sc_hd__and2_1 _13611_ (.A(_06657_),
    .B(_06658_),
    .X(_06762_));
 sky130_fd_sc_hd__o31a_1 _13612_ (.A1(_06743_),
    .A2(_06758_),
    .A3(_06761_),
    .B1(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__a221o_1 _13613_ (.A1(_06752_),
    .A2(_06701_),
    .B1(_06756_),
    .B2(_06763_),
    .C1(_06589_),
    .X(_06764_));
 sky130_fd_sc_hd__a21oi_4 _13614_ (.A1(net7431),
    .A2(_06714_),
    .B1(net7433),
    .Y(_06765_));
 sky130_fd_sc_hd__nand2_1 _13615_ (.A(_06732_),
    .B(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__a21oi_1 _13616_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06614_),
    .Y(_06767_));
 sky130_fd_sc_hd__a211o_1 _13617_ (.A1(_06616_),
    .A2(_06688_),
    .B1(_06767_),
    .C1(_06677_),
    .X(_06768_));
 sky130_fd_sc_hd__and3_1 _13618_ (.A(_06669_),
    .B(_06693_),
    .C(_06694_),
    .X(_06769_));
 sky130_fd_sc_hd__a21oi_1 _13619_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06621_),
    .Y(_06770_));
 sky130_fd_sc_hd__or3_1 _13620_ (.A(_06691_),
    .B(_06769_),
    .C(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a21o_1 _13621_ (.A1(_06768_),
    .A2(_06771_),
    .B1(_06743_),
    .X(_06772_));
 sky130_fd_sc_hd__or3_1 _13622_ (.A(_06600_),
    .B(_06667_),
    .C(_06686_),
    .X(_06773_));
 sky130_fd_sc_hd__a21o_1 _13623_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06627_),
    .X(_06774_));
 sky130_fd_sc_hd__and3_1 _13624_ (.A(_06676_),
    .B(_06773_),
    .C(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__a21o_1 _13625_ (.A1(_06693_),
    .A2(_06694_),
    .B1(_06606_),
    .X(_06776_));
 sky130_fd_sc_hd__or3_1 _13626_ (.A(_06727_),
    .B(_06667_),
    .C(_06686_),
    .X(_06777_));
 sky130_fd_sc_hd__a21oi_1 _13627_ (.A1(_06776_),
    .A2(_06777_),
    .B1(_06677_),
    .Y(_06778_));
 sky130_fd_sc_hd__or3_1 _13628_ (.A(_06662_),
    .B(_06775_),
    .C(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__a21oi_2 _13629_ (.A1(_06772_),
    .A2(_06779_),
    .B1(_06659_),
    .Y(_06780_));
 sky130_fd_sc_hd__a221o_2 _13630_ (.A1(_06660_),
    .A2(_06751_),
    .B1(_06764_),
    .B2(_06766_),
    .C1(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__nand2_1 _13631_ (.A(_06747_),
    .B(_06748_),
    .Y(_06782_));
 sky130_fd_sc_hd__a21oi_1 _13632_ (.A1(_06773_),
    .A2(_06774_),
    .B1(_06677_),
    .Y(_06783_));
 sky130_fd_sc_hd__a21o_1 _13633_ (.A1(_06677_),
    .A2(_06782_),
    .B1(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__and3_1 _13634_ (.A(_06676_),
    .B(_06776_),
    .C(_06777_),
    .X(_06785_));
 sky130_fd_sc_hd__or3_1 _13635_ (.A(_06676_),
    .B(_06769_),
    .C(_06770_),
    .X(_06786_));
 sky130_fd_sc_hd__or3b_1 _13636_ (.A(_06743_),
    .B(_06785_),
    .C_N(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__clkbuf_2 _13637_ (.A(_06762_),
    .X(_06788_));
 sky130_fd_sc_hd__o211a_1 _13638_ (.A1(_06662_),
    .A2(_06784_),
    .B1(_06787_),
    .C1(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__nand2_1 _13639_ (.A(_06744_),
    .B(_06745_),
    .Y(_06790_));
 sky130_fd_sc_hd__mux2_1 _13640_ (.A0(_06790_),
    .A1(_06740_),
    .S(_06677_),
    .X(_06791_));
 sky130_fd_sc_hd__a21o_1 _13641_ (.A1(_06662_),
    .A2(_06791_),
    .B1(_06589_),
    .X(_06792_));
 sky130_fd_sc_hd__a21o_1 _13642_ (.A1(_06616_),
    .A2(_06688_),
    .B1(_06770_),
    .X(_06793_));
 sky130_fd_sc_hd__a22o_1 _13643_ (.A1(_06677_),
    .A2(_06767_),
    .B1(_06793_),
    .B2(_06717_),
    .X(_06794_));
 sky130_fd_sc_hd__nand2_1 _13644_ (.A(_06725_),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__o22a_4 _13645_ (.A1(_06789_),
    .A2(_06792_),
    .B1(_06795_),
    .B2(_06716_),
    .X(_06796_));
 sky130_fd_sc_hd__o21ai_1 _13646_ (.A1(_06775_),
    .A2(_06778_),
    .B1(_06662_),
    .Y(_06797_));
 sky130_fd_sc_hd__o31a_1 _13647_ (.A1(_06662_),
    .A2(_06746_),
    .A3(_06749_),
    .B1(_06762_),
    .X(_06798_));
 sky130_fd_sc_hd__a22o_1 _13648_ (.A1(_06752_),
    .A2(_06741_),
    .B1(_06797_),
    .B2(_06798_),
    .X(_06799_));
 sky130_fd_sc_hd__xnor2_2 _13649_ (.A(_06742_),
    .B(_06713_),
    .Y(_06800_));
 sky130_fd_sc_hd__inv_2 _13650_ (.A(_06616_),
    .Y(_06801_));
 sky130_fd_sc_hd__mux4_1 _13651_ (.A0(_06606_),
    .A1(_06801_),
    .A2(_06621_),
    .A3(_06619_),
    .S0(_06687_),
    .S1(_06677_),
    .X(_06802_));
 sky130_fd_sc_hd__nor2_1 _13652_ (.A(_06800_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__and3_1 _13653_ (.A(_06743_),
    .B(_06707_),
    .C(_06767_),
    .X(_06804_));
 sky130_fd_sc_hd__o21a_1 _13654_ (.A1(_06803_),
    .A2(_06804_),
    .B1(_06765_),
    .X(_06805_));
 sky130_fd_sc_hd__o21ba_1 _13655_ (.A1(_06589_),
    .A2(_06799_),
    .B1_N(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__a21oi_1 _13656_ (.A1(_06638_),
    .A2(_06687_),
    .B1(_06718_),
    .Y(_06807_));
 sky130_fd_sc_hd__mux2_1 _13657_ (.A0(_06696_),
    .A1(_06807_),
    .S(_06692_),
    .X(_06808_));
 sky130_fd_sc_hd__a211o_1 _13658_ (.A1(_06608_),
    .A2(_06688_),
    .B1(_06753_),
    .C1(_06692_),
    .X(_06809_));
 sky130_fd_sc_hd__or3_1 _13659_ (.A(_06676_),
    .B(_06759_),
    .C(_06760_),
    .X(_06810_));
 sky130_fd_sc_hd__a21oi_1 _13660_ (.A1(_06809_),
    .A2(_06810_),
    .B1(_06743_),
    .Y(_06811_));
 sky130_fd_sc_hd__a211o_1 _13661_ (.A1(_06743_),
    .A2(_06808_),
    .B1(_06811_),
    .C1(_06659_),
    .X(_06812_));
 sky130_fd_sc_hd__a21oi_1 _13662_ (.A1(net539),
    .A2(_06688_),
    .B1(_06699_),
    .Y(_06813_));
 sky130_fd_sc_hd__mux2_1 _13663_ (.A0(_06813_),
    .A1(_06704_),
    .S(_06677_),
    .X(_06814_));
 sky130_fd_sc_hd__or2_1 _13664_ (.A(_06657_),
    .B(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__o21a_1 _13665_ (.A1(_06669_),
    .A2(_06687_),
    .B1(_06757_),
    .X(_06816_));
 sky130_fd_sc_hd__mux2_1 _13666_ (.A0(_06731_),
    .A1(_06816_),
    .S(_06717_),
    .X(_06817_));
 sky130_fd_sc_hd__and3_1 _13667_ (.A(_06724_),
    .B(_06765_),
    .C(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__a31oi_4 _13668_ (.A1(_06733_),
    .A2(_06812_),
    .A3(_06815_),
    .B1(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__a211oi_1 _13669_ (.A1(_06707_),
    .A2(_06696_),
    .B1(_06700_),
    .C1(_06662_),
    .Y(_06820_));
 sky130_fd_sc_hd__and3_1 _13670_ (.A(_06662_),
    .B(_06754_),
    .C(_06755_),
    .X(_06821_));
 sky130_fd_sc_hd__o21ai_1 _13671_ (.A1(_06820_),
    .A2(_06821_),
    .B1(_06788_),
    .Y(_06822_));
 sky130_fd_sc_hd__o21a_1 _13672_ (.A1(_06657_),
    .A2(_06705_),
    .B1(_06733_),
    .X(_06823_));
 sky130_fd_sc_hd__nand2_1 _13673_ (.A(_06717_),
    .B(_06731_),
    .Y(_06824_));
 sky130_fd_sc_hd__mux2_1 _13674_ (.A0(_06824_),
    .A1(_06728_),
    .S(_06724_),
    .X(_06825_));
 sky130_fd_sc_hd__o2bb2a_4 _13675_ (.A1_N(_06822_),
    .A2_N(_06823_),
    .B1(_06716_),
    .B2(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__a2111o_1 _13676_ (.A1(_06781_),
    .A2(_06796_),
    .B1(_06806_),
    .C1(net562),
    .D1(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__mux4_1 _13677_ (.A0(_06606_),
    .A1(_06608_),
    .A2(_06727_),
    .A3(_06619_),
    .S0(_06692_),
    .S1(_06688_),
    .X(_06828_));
 sky130_fd_sc_hd__nor2_1 _13678_ (.A(_06725_),
    .B(_06794_),
    .Y(_06829_));
 sky130_fd_sc_hd__a211o_1 _13679_ (.A1(_06725_),
    .A2(_06828_),
    .B1(_06829_),
    .C1(_06716_),
    .X(_06830_));
 sky130_fd_sc_hd__nand2_1 _13680_ (.A(_06662_),
    .B(_06784_),
    .Y(_06831_));
 sky130_fd_sc_hd__or3b_2 _13681_ (.A(_06659_),
    .B(_06791_),
    .C_N(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__mux2_1 _13682_ (.A0(_06567_),
    .A1(_06565_),
    .S(_06688_),
    .X(_06833_));
 sky130_fd_sc_hd__mux2_1 _13683_ (.A0(_06739_),
    .A1(_06833_),
    .S(_06678_),
    .X(_06834_));
 sky130_fd_sc_hd__or2_1 _13684_ (.A(_06743_),
    .B(_06834_),
    .X(_06835_));
 sky130_fd_sc_hd__and3_1 _13685_ (.A(_06830_),
    .B(_06832_),
    .C(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__buf_4 _13686_ (.A(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__clkbuf_2 _13687_ (.A(_06743_),
    .X(_06838_));
 sky130_fd_sc_hd__mux2_1 _13688_ (.A0(_06808_),
    .A1(_06814_),
    .S(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__nor2_1 _13689_ (.A(_06759_),
    .B(_06753_),
    .Y(_06840_));
 sky130_fd_sc_hd__mux4_1 _13690_ (.A0(_06731_),
    .A1(_06840_),
    .A2(_06816_),
    .A3(_06719_),
    .S0(_06724_),
    .S1(_06717_),
    .X(_06841_));
 sky130_fd_sc_hd__nor2_1 _13691_ (.A(_06707_),
    .B(_06708_),
    .Y(_06842_));
 sky130_fd_sc_hd__a221o_1 _13692_ (.A1(_06707_),
    .A2(_06703_),
    .B1(_06765_),
    .B2(_06841_),
    .C1(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__a21o_4 _13693_ (.A1(_06788_),
    .A2(_06839_),
    .B1(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__a21bo_1 _13694_ (.A1(net3132),
    .A2(_06837_),
    .B1_N(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__buf_6 _13695_ (.A(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__nor2_1 _13696_ (.A(_06660_),
    .B(_06751_),
    .Y(_06847_));
 sky130_fd_sc_hd__mux2_1 _13697_ (.A0(_06584_),
    .A1(_06586_),
    .S(_06722_),
    .X(_06848_));
 sky130_fd_sc_hd__mux2_1 _13698_ (.A0(_06833_),
    .A1(_06848_),
    .S(_06678_),
    .X(_06849_));
 sky130_fd_sc_hd__nand2_1 _13699_ (.A(_06733_),
    .B(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__and3_1 _13700_ (.A(_06421_),
    .B(_06663_),
    .C(_06713_),
    .X(_06851_));
 sky130_fd_sc_hd__mux4_1 _13701_ (.A0(_06591_),
    .A1(_06627_),
    .A2(_06603_),
    .A3(_06600_),
    .S0(_06677_),
    .S1(_06688_),
    .X(_06852_));
 sky130_fd_sc_hd__nand2_1 _13702_ (.A(_06800_),
    .B(_06802_),
    .Y(_06853_));
 sky130_fd_sc_hd__o21a_1 _13703_ (.A1(_06800_),
    .A2(_06852_),
    .B1(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__mux2_1 _13704_ (.A0(_06851_),
    .A1(_06854_),
    .S(_06715_),
    .X(_06855_));
 sky130_fd_sc_hd__o22ai_2 _13705_ (.A1(_06847_),
    .A2(_06850_),
    .B1(_06855_),
    .B2(_06733_),
    .Y(_06856_));
 sky130_fd_sc_hd__nor2_8 _13706_ (.A(_06846_),
    .B(net79),
    .Y(_06857_));
 sky130_fd_sc_hd__xnor2_4 _13707_ (.A(_06737_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__clkbuf_4 _13708_ (.A(net573),
    .X(_06859_));
 sky130_fd_sc_hd__a21o_4 _13709_ (.A1(_06660_),
    .A2(_06751_),
    .B1(net582),
    .X(_06860_));
 sky130_fd_sc_hd__clkbuf_4 _13710_ (.A(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__clkbuf_4 _13711_ (.A(_06861_),
    .X(_06862_));
 sky130_fd_sc_hd__and2_1 _13712_ (.A(_06764_),
    .B(_06766_),
    .X(_06863_));
 sky130_fd_sc_hd__buf_4 _13713_ (.A(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__buf_4 _13714_ (.A(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__inv_2 _13715_ (.A(_06737_),
    .Y(_06866_));
 sky130_fd_sc_hd__a21o_2 _13716_ (.A1(_06866_),
    .A2(_06857_),
    .B1(_06668_),
    .X(_06867_));
 sky130_fd_sc_hd__or4_4 _13717_ (.A(_06862_),
    .B(_06865_),
    .C(_06858_),
    .D(_06867_),
    .X(_06868_));
 sky130_fd_sc_hd__clkbuf_4 _13718_ (.A(_06796_),
    .X(_06869_));
 sky130_fd_sc_hd__nor2_1 _13719_ (.A(_06869_),
    .B(_06858_),
    .Y(_06870_));
 sky130_fd_sc_hd__nor2_1 _13720_ (.A(_06865_),
    .B(_06867_),
    .Y(_06871_));
 sky130_fd_sc_hd__xnor2_2 _13721_ (.A(_06870_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__nor2_1 _13722_ (.A(_06868_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_1 _13723_ (.A(_06870_),
    .B(_06871_),
    .Y(_06874_));
 sky130_fd_sc_hd__or2_1 _13724_ (.A(_06869_),
    .B(_06867_),
    .X(_06875_));
 sky130_fd_sc_hd__buf_2 _13725_ (.A(net553),
    .X(_06876_));
 sky130_fd_sc_hd__nor2_1 _13726_ (.A(_06876_),
    .B(_06858_),
    .Y(_06877_));
 sky130_fd_sc_hd__xnor2_1 _13727_ (.A(_06875_),
    .B(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__xnor2_1 _13728_ (.A(_06874_),
    .B(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__buf_2 _13729_ (.A(_06844_),
    .X(_06880_));
 sky130_fd_sc_hd__nand3_4 _13730_ (.A(_06830_),
    .B(_06832_),
    .C(_06835_),
    .Y(_06881_));
 sky130_fd_sc_hd__a21o_2 _13731_ (.A1(net584),
    .A2(_06796_),
    .B1(_06819_),
    .X(_06882_));
 sky130_fd_sc_hd__nand3_1 _13732_ (.A(net580),
    .B(_06819_),
    .C(_06796_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_1 _13733_ (.A(net578),
    .B(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__clkbuf_8 _13734_ (.A(_06806_),
    .X(_06885_));
 sky130_fd_sc_hd__xnor2_4 _13735_ (.A(net579),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand4_4 _13736_ (.A(_06880_),
    .B(_06881_),
    .C(_06884_),
    .D(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__a211o_2 _13737_ (.A1(_06781_),
    .A2(_06796_),
    .B1(_06806_),
    .C1(net563),
    .X(_06888_));
 sky130_fd_sc_hd__nor2_2 _13738_ (.A(_06826_),
    .B(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__a22o_1 _13739_ (.A1(_06844_),
    .A2(_06884_),
    .B1(_06886_),
    .B2(_06881_),
    .X(_06890_));
 sky130_fd_sc_hd__nand3_2 _13740_ (.A(_06889_),
    .B(_06887_),
    .C(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__and2_1 _13741_ (.A(_06887_),
    .B(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__xor2_2 _13742_ (.A(_06846_),
    .B(net79),
    .X(_06893_));
 sky130_fd_sc_hd__nor2_1 _13743_ (.A(_06876_),
    .B(net572),
    .Y(_06894_));
 sky130_fd_sc_hd__clkbuf_4 _13744_ (.A(_06826_),
    .X(_06895_));
 sky130_fd_sc_hd__xnor2_4 _13745_ (.A(net540),
    .B(_06837_),
    .Y(_06896_));
 sky130_fd_sc_hd__nor2_1 _13746_ (.A(_06895_),
    .B(net547),
    .Y(_06897_));
 sky130_fd_sc_hd__or3b_4 _13747_ (.A(_06844_),
    .B(_06881_),
    .C_N(_06827_),
    .X(_06898_));
 sky130_fd_sc_hd__a21oi_2 _13748_ (.A1(net3370),
    .A2(_06898_),
    .B1(_06885_),
    .Y(_06899_));
 sky130_fd_sc_hd__xnor2_2 _13749_ (.A(_06897_),
    .B(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__xnor2_2 _13750_ (.A(_06894_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__and2b_1 _13751_ (.A_N(_06892_),
    .B(net576),
    .X(_06902_));
 sky130_fd_sc_hd__nor2_2 _13752_ (.A(_06885_),
    .B(net546),
    .Y(_06903_));
 sky130_fd_sc_hd__a21oi_2 _13753_ (.A1(_06846_),
    .A2(_06898_),
    .B1(net554),
    .Y(_06904_));
 sky130_fd_sc_hd__or2_4 _13754_ (.A(_06869_),
    .B(_06893_),
    .X(_06905_));
 sky130_fd_sc_hd__xnor2_2 _13755_ (.A(_06903_),
    .B(_06904_),
    .Y(_06906_));
 sky130_fd_sc_hd__nor2_1 _13756_ (.A(_06905_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__a21o_1 _13757_ (.A1(_06903_),
    .A2(_06904_),
    .B1(_06907_),
    .X(_06908_));
 sky130_fd_sc_hd__xnor2_2 _13758_ (.A(_06892_),
    .B(_06901_),
    .Y(_06909_));
 sky130_fd_sc_hd__and2_1 _13759_ (.A(_06908_),
    .B(net575),
    .X(_06910_));
 sky130_fd_sc_hd__or3_1 _13760_ (.A(_06879_),
    .B(_06902_),
    .C(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__o21a_1 _13761_ (.A1(_06902_),
    .A2(_06910_),
    .B1(_06879_),
    .X(_06912_));
 sky130_fd_sc_hd__a21o_1 _13762_ (.A1(_06873_),
    .A2(_06911_),
    .B1(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__xor2_1 _13763_ (.A(_06860_),
    .B(_06864_),
    .X(_06914_));
 sky130_fd_sc_hd__or3_4 _13764_ (.A(_06736_),
    .B(_06860_),
    .C(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__xnor2_2 _13765_ (.A(net561),
    .B(_06796_),
    .Y(_06916_));
 sky130_fd_sc_hd__nor2_1 _13766_ (.A(net79),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__buf_4 _13767_ (.A(_06914_),
    .X(_06918_));
 sky130_fd_sc_hd__o21ai_2 _13768_ (.A1(_06736_),
    .A2(_06918_),
    .B1(_06861_),
    .Y(_06919_));
 sky130_fd_sc_hd__nand3_4 _13769_ (.A(_06915_),
    .B(_06917_),
    .C(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__or4_2 _13770_ (.A(_06668_),
    .B(_06736_),
    .C(_06918_),
    .D(_06916_),
    .X(_06921_));
 sky130_fd_sc_hd__buf_6 _13771_ (.A(_06916_),
    .X(_06922_));
 sky130_fd_sc_hd__xnor2_4 _13772_ (.A(_06860_),
    .B(_06864_),
    .Y(_06923_));
 sky130_fd_sc_hd__a2bb2o_1 _13773_ (.A1_N(_06736_),
    .A2_N(_06922_),
    .B1(_06923_),
    .B2(_06611_),
    .X(_06924_));
 sky130_fd_sc_hd__nand2_1 _13774_ (.A(_06921_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__a21o_1 _13775_ (.A1(_06915_),
    .A2(_06920_),
    .B1(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__nand3_1 _13776_ (.A(_06925_),
    .B(_06915_),
    .C(_06920_),
    .Y(_06927_));
 sky130_fd_sc_hd__and2_1 _13777_ (.A(_06926_),
    .B(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__xor2_2 _13778_ (.A(_06826_),
    .B(_06888_),
    .X(_06929_));
 sky130_fd_sc_hd__or2_1 _13779_ (.A(_06837_),
    .B(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__buf_2 _13780_ (.A(net79),
    .X(_06931_));
 sky130_fd_sc_hd__and4b_1 _13781_ (.A_N(_06931_),
    .B(_06884_),
    .C(_06886_),
    .D(_06880_),
    .X(_06932_));
 sky130_fd_sc_hd__and2_4 _13782_ (.A(_06882_),
    .B(_06883_),
    .X(_06933_));
 sky130_fd_sc_hd__o2bb2a_1 _13783_ (.A1_N(_06880_),
    .A2_N(_06886_),
    .B1(_06933_),
    .B2(_06931_),
    .X(_06934_));
 sky130_fd_sc_hd__nor2_1 _13784_ (.A(_06932_),
    .B(_06934_),
    .Y(_06935_));
 sky130_fd_sc_hd__xnor2_2 _13785_ (.A(_06930_),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__xor2_2 _13786_ (.A(_06928_),
    .B(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__a21o_1 _13787_ (.A1(_06915_),
    .A2(_06919_),
    .B1(_06917_),
    .X(_06938_));
 sky130_fd_sc_hd__and2b_1 _13788_ (.A_N(_06844_),
    .B(_06916_),
    .X(_06939_));
 sky130_fd_sc_hd__o22ai_2 _13789_ (.A1(_06736_),
    .A2(_06861_),
    .B1(net79),
    .B2(_06918_),
    .Y(_06940_));
 sky130_fd_sc_hd__or4_4 _13790_ (.A(_06736_),
    .B(_06860_),
    .C(net79),
    .D(_06914_),
    .X(_06941_));
 sky130_fd_sc_hd__a21bo_1 _13791_ (.A1(_06939_),
    .A2(_06940_),
    .B1_N(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__nand3_1 _13792_ (.A(_06920_),
    .B(_06938_),
    .C(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__a21o_1 _13793_ (.A1(_06920_),
    .A2(_06938_),
    .B1(_06942_),
    .X(_06944_));
 sky130_fd_sc_hd__a21o_1 _13794_ (.A1(_06887_),
    .A2(_06890_),
    .B1(_06889_),
    .X(_06945_));
 sky130_fd_sc_hd__and4_1 _13795_ (.A(_06891_),
    .B(_06943_),
    .C(_06944_),
    .D(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__a31oi_4 _13796_ (.A1(_06920_),
    .A2(_06938_),
    .A3(net565),
    .B1(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__xnor2_2 _13797_ (.A(_06937_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__xor2_2 _13798_ (.A(_06908_),
    .B(_06909_),
    .X(_06949_));
 sky130_fd_sc_hd__or2b_1 _13799_ (.A(_06947_),
    .B_N(_06937_),
    .X(_06950_));
 sky130_fd_sc_hd__a21bo_1 _13800_ (.A1(_06948_),
    .A2(_06949_),
    .B1_N(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__or2b_1 _13801_ (.A(_06922_),
    .B_N(_06921_),
    .X(_06952_));
 sky130_fd_sc_hd__inv_2 _13802_ (.A(_06929_),
    .Y(_06953_));
 sky130_fd_sc_hd__nand2_1 _13803_ (.A(_06880_),
    .B(_06953_),
    .Y(_06954_));
 sky130_fd_sc_hd__xor2_4 _13804_ (.A(_06882_),
    .B(_06885_),
    .X(_06955_));
 sky130_fd_sc_hd__or2_1 _13805_ (.A(_06931_),
    .B(_06955_),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_4 _13806_ (.A(_06933_),
    .X(_06957_));
 sky130_fd_sc_hd__nor2_1 _13807_ (.A(_06737_),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__xnor2_2 _13808_ (.A(_06956_),
    .B(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__xnor2_2 _13809_ (.A(_06954_),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__xnor2_1 _13810_ (.A(_06952_),
    .B(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__a21bo_1 _13811_ (.A1(_06928_),
    .A2(_06936_),
    .B1_N(_06926_),
    .X(_06962_));
 sky130_fd_sc_hd__and2_1 _13812_ (.A(_06961_),
    .B(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__nor2_1 _13813_ (.A(_06961_),
    .B(_06962_),
    .Y(_06964_));
 sky130_fd_sc_hd__or2_1 _13814_ (.A(_06963_),
    .B(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__buf_6 _13815_ (.A(_06893_),
    .X(_06966_));
 sky130_fd_sc_hd__or3_1 _13816_ (.A(_06876_),
    .B(net529),
    .C(net577),
    .X(_06967_));
 sky130_fd_sc_hd__a21bo_1 _13817_ (.A1(_06897_),
    .A2(_06899_),
    .B1_N(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__a31o_1 _13818_ (.A1(_06881_),
    .A2(_06953_),
    .A3(_06935_),
    .B1(_06932_),
    .X(_06969_));
 sky130_fd_sc_hd__buf_2 _13819_ (.A(_06885_),
    .X(_06970_));
 sky130_fd_sc_hd__or2_1 _13820_ (.A(_06970_),
    .B(net529),
    .X(_06971_));
 sky130_fd_sc_hd__and2_4 _13821_ (.A(_06846_),
    .B(_06898_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_6 _13822_ (.A(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__nor2_1 _13823_ (.A(_06895_),
    .B(_06973_),
    .Y(_06974_));
 sky130_fd_sc_hd__nor2_1 _13824_ (.A(_06889_),
    .B(_06837_),
    .Y(_06975_));
 sky130_fd_sc_hd__xor2_2 _13825_ (.A(_06974_),
    .B(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__xnor2_2 _13826_ (.A(_06971_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__xnor2_2 _13827_ (.A(_06969_),
    .B(_06977_),
    .Y(_06978_));
 sky130_fd_sc_hd__xor2_2 _13828_ (.A(_06968_),
    .B(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__xnor2_2 _13829_ (.A(_06965_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__xor2_2 _13830_ (.A(_06951_),
    .B(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__and2b_1 _13831_ (.A_N(_06912_),
    .B(_06911_),
    .X(_06982_));
 sky130_fd_sc_hd__xnor2_2 _13832_ (.A(_06873_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__or2b_1 _13833_ (.A(_06980_),
    .B_N(_06951_),
    .X(_06984_));
 sky130_fd_sc_hd__o21ai_2 _13834_ (.A1(_06981_),
    .A2(_06983_),
    .B1(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__nor2_1 _13835_ (.A(_06965_),
    .B(_06979_),
    .Y(_06986_));
 sky130_fd_sc_hd__nand2_1 _13836_ (.A(_06866_),
    .B(_06886_),
    .Y(_06987_));
 sky130_fd_sc_hd__o21ai_1 _13837_ (.A1(_06668_),
    .A2(_06957_),
    .B1(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__o21a_1 _13838_ (.A1(_06957_),
    .A2(_06987_),
    .B1(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__clkbuf_4 _13839_ (.A(_06929_),
    .X(_06990_));
 sky130_fd_sc_hd__nor2_1 _13840_ (.A(_06931_),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__xnor2_1 _13841_ (.A(_06989_),
    .B(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__inv_2 _13842_ (.A(_06960_),
    .Y(_06993_));
 sky130_fd_sc_hd__o21a_1 _13843_ (.A1(_06922_),
    .A2(_06993_),
    .B1(_06921_),
    .X(_06994_));
 sky130_fd_sc_hd__xor2_1 _13844_ (.A(_06992_),
    .B(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__and2b_1 _13845_ (.A_N(_06971_),
    .B(_06976_),
    .X(_06996_));
 sky130_fd_sc_hd__a21oi_1 _13846_ (.A1(_06974_),
    .A2(_06975_),
    .B1(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__and2b_1 _13847_ (.A_N(_06956_),
    .B(_06958_),
    .X(_06998_));
 sky130_fd_sc_hd__and3_1 _13848_ (.A(_06880_),
    .B(_06953_),
    .C(_06959_),
    .X(_06999_));
 sky130_fd_sc_hd__inv_2 _13849_ (.A(net530),
    .Y(_07000_));
 sky130_fd_sc_hd__o2bb2a_1 _13850_ (.A1_N(_06880_),
    .A2_N(_06889_),
    .B1(net529),
    .B2(_06895_),
    .X(_07001_));
 sky130_fd_sc_hd__a31oi_2 _13851_ (.A1(_06880_),
    .A2(_06889_),
    .A3(_07000_),
    .B1(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__o21a_1 _13852_ (.A1(_06998_),
    .A2(_06999_),
    .B1(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__nor3_1 _13853_ (.A(_06998_),
    .B(_06999_),
    .C(_07002_),
    .Y(_07004_));
 sky130_fd_sc_hd__nor2_1 _13854_ (.A(_07003_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__xnor2_1 _13855_ (.A(_06997_),
    .B(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__xor2_1 _13856_ (.A(_06995_),
    .B(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__o21a_1 _13857_ (.A1(_06963_),
    .A2(_06986_),
    .B1(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__nor3_1 _13858_ (.A(_06963_),
    .B(_06986_),
    .C(_07007_),
    .Y(_07009_));
 sky130_fd_sc_hd__or2_1 _13859_ (.A(_07008_),
    .B(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__or2b_1 _13860_ (.A(_06874_),
    .B_N(_06878_),
    .X(_07011_));
 sky130_fd_sc_hd__and2b_1 _13861_ (.A_N(_06978_),
    .B(_06968_),
    .X(_07012_));
 sky130_fd_sc_hd__a21o_1 _13862_ (.A1(_06969_),
    .A2(_06977_),
    .B1(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__or3_1 _13863_ (.A(_06876_),
    .B(_06859_),
    .C(_06875_),
    .X(_07014_));
 sky130_fd_sc_hd__or2_1 _13864_ (.A(_06876_),
    .B(_06867_),
    .X(_07015_));
 sky130_fd_sc_hd__or3_1 _13865_ (.A(_06970_),
    .B(_06858_),
    .C(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__o21ai_1 _13866_ (.A1(_06970_),
    .A2(_06859_),
    .B1(_07015_),
    .Y(_07017_));
 sky130_fd_sc_hd__and2_1 _13867_ (.A(_07016_),
    .B(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__xnor2_1 _13868_ (.A(_07014_),
    .B(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__xnor2_1 _13869_ (.A(_07013_),
    .B(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__xnor2_1 _13870_ (.A(_07011_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__xor2_1 _13871_ (.A(_07010_),
    .B(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__xnor2_1 _13872_ (.A(_06985_),
    .B(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__xnor2_1 _13873_ (.A(_06913_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__xnor2_4 _13874_ (.A(_06905_),
    .B(_06906_),
    .Y(_07025_));
 sky130_fd_sc_hd__or4_4 _13875_ (.A(_06826_),
    .B(_06837_),
    .C(_06933_),
    .D(_06955_),
    .X(_07026_));
 sky130_fd_sc_hd__or2_1 _13876_ (.A(_06885_),
    .B(_06929_),
    .X(_07027_));
 sky130_fd_sc_hd__o22ai_1 _13877_ (.A1(_06837_),
    .A2(_06957_),
    .B1(_06955_),
    .B2(_06895_),
    .Y(_07028_));
 sky130_fd_sc_hd__nand3b_1 _13878_ (.A_N(_07027_),
    .B(_07026_),
    .C(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__nand2_1 _13879_ (.A(_07026_),
    .B(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__and2b_1 _13880_ (.A_N(_07025_),
    .B(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__nor2_2 _13881_ (.A(_06864_),
    .B(_06966_),
    .Y(_07032_));
 sky130_fd_sc_hd__or2_1 _13882_ (.A(net554),
    .B(_06896_),
    .X(_07033_));
 sky130_fd_sc_hd__a21oi_1 _13883_ (.A1(net3408),
    .A2(_06898_),
    .B1(_06796_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_2 _13884_ (.A(_07033_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__or3_4 _13885_ (.A(_06869_),
    .B(_06973_),
    .C(_07033_),
    .X(_07036_));
 sky130_fd_sc_hd__a21bo_4 _13886_ (.A1(_07032_),
    .A2(net570),
    .B1_N(_07036_),
    .X(_07037_));
 sky130_fd_sc_hd__xnor2_2 _13887_ (.A(_07030_),
    .B(_07025_),
    .Y(_07038_));
 sky130_fd_sc_hd__and2_4 _13888_ (.A(_07037_),
    .B(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__xor2_2 _13889_ (.A(_06868_),
    .B(_06872_),
    .X(_07040_));
 sky130_fd_sc_hd__o21ai_4 _13890_ (.A1(_07031_),
    .A2(_07039_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__inv_2 _13891_ (.A(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__a22o_1 _13892_ (.A1(_06943_),
    .A2(_06944_),
    .B1(net585),
    .B2(_06891_),
    .X(_07043_));
 sky130_fd_sc_hd__or2b_4 _13893_ (.A(_06946_),
    .B_N(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__nand3_1 _13894_ (.A(_06941_),
    .B(_06939_),
    .C(_06940_),
    .Y(_07045_));
 sky130_fd_sc_hd__a21o_1 _13895_ (.A1(_06941_),
    .A2(_06940_),
    .B1(_06939_),
    .X(_07046_));
 sky130_fd_sc_hd__nor2_1 _13896_ (.A(_06837_),
    .B(_06922_),
    .Y(_07047_));
 sky130_fd_sc_hd__a2bb2o_1 _13897_ (.A1_N(_06861_),
    .A2_N(net79),
    .B1(_06923_),
    .B2(_06844_),
    .X(_07048_));
 sky130_fd_sc_hd__or4b_1 _13898_ (.A(_06861_),
    .B(net79),
    .C(_06864_),
    .D_N(_06844_),
    .X(_07049_));
 sky130_fd_sc_hd__a21bo_1 _13899_ (.A1(_07047_),
    .A2(_07048_),
    .B1_N(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__and3_1 _13900_ (.A(_07045_),
    .B(_07046_),
    .C(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__a21oi_1 _13901_ (.A1(_07045_),
    .A2(_07046_),
    .B1(_07050_),
    .Y(_07052_));
 sky130_fd_sc_hd__nor2_1 _13902_ (.A(_07051_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__a21bo_1 _13903_ (.A1(_07026_),
    .A2(_07028_),
    .B1_N(_07027_),
    .X(_07054_));
 sky130_fd_sc_hd__and2_4 _13904_ (.A(_07029_),
    .B(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__a21o_1 _13905_ (.A1(_07053_),
    .A2(_07055_),
    .B1(_07051_),
    .X(_07056_));
 sky130_fd_sc_hd__xnor2_2 _13906_ (.A(_07044_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__xor2_2 _13907_ (.A(_07037_),
    .B(_07038_),
    .X(_07058_));
 sky130_fd_sc_hd__and2b_1 _13908_ (.A_N(_07044_),
    .B(_07056_),
    .X(_07059_));
 sky130_fd_sc_hd__a21oi_2 _13909_ (.A1(_07057_),
    .A2(net1998),
    .B1(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__xnor2_2 _13910_ (.A(_06948_),
    .B(_06949_),
    .Y(_07061_));
 sky130_fd_sc_hd__xnor2_2 _13911_ (.A(_07060_),
    .B(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__or3_1 _13912_ (.A(_07031_),
    .B(_07039_),
    .C(_07040_),
    .X(_07063_));
 sky130_fd_sc_hd__and2_4 _13913_ (.A(_07041_),
    .B(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__or2b_1 _13914_ (.A(net566),
    .B_N(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__o21a_1 _13915_ (.A1(_07060_),
    .A2(_07061_),
    .B1(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__xor2_2 _13916_ (.A(_06981_),
    .B(_06983_),
    .X(_07067_));
 sky130_fd_sc_hd__xnor2_2 _13917_ (.A(_07066_),
    .B(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__and2b_1 _13918_ (.A_N(_07066_),
    .B(_07067_),
    .X(_07069_));
 sky130_fd_sc_hd__a21oi_1 _13919_ (.A1(_07042_),
    .A2(_07068_),
    .B1(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__xor2_1 _13920_ (.A(_07024_),
    .B(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__xnor2_2 _13921_ (.A(_07032_),
    .B(_07035_),
    .Y(_07072_));
 sky130_fd_sc_hd__xnor2_2 _13922_ (.A(net556),
    .B(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__nor2_1 _13923_ (.A(_06865_),
    .B(net564),
    .Y(_07074_));
 sky130_fd_sc_hd__nor2_1 _13924_ (.A(_06796_),
    .B(_06896_),
    .Y(_07075_));
 sky130_fd_sc_hd__nor2_8 _13925_ (.A(_06966_),
    .B(_06862_),
    .Y(_07076_));
 sky130_fd_sc_hd__a21o_1 _13926_ (.A1(_06846_),
    .A2(_06898_),
    .B1(_06864_),
    .X(_07077_));
 sky130_fd_sc_hd__xnor2_2 _13927_ (.A(_07077_),
    .B(_07075_),
    .Y(_07078_));
 sky130_fd_sc_hd__a22o_1 _13928_ (.A1(_07074_),
    .A2(_07075_),
    .B1(net571),
    .B2(net574),
    .X(_07079_));
 sky130_fd_sc_hd__or2b_1 _13929_ (.A(_07073_),
    .B_N(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__o21ai_2 _13930_ (.A1(net557),
    .A2(_07072_),
    .B1(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__xnor2_2 _13931_ (.A(_06866_),
    .B(net567),
    .Y(_07082_));
 sky130_fd_sc_hd__inv_2 _13932_ (.A(_06865_),
    .Y(_07083_));
 sky130_fd_sc_hd__a2bb2o_1 _13933_ (.A1_N(_06862_),
    .A2_N(_06867_),
    .B1(_07082_),
    .B2(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__and3_1 _13934_ (.A(net3405),
    .B(_07081_),
    .C(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__xor2_2 _13935_ (.A(_07053_),
    .B(_07055_),
    .X(_07086_));
 sky130_fd_sc_hd__nand3_1 _13936_ (.A(_07049_),
    .B(_07047_),
    .C(_07048_),
    .Y(_07087_));
 sky130_fd_sc_hd__a21o_1 _13937_ (.A1(_07049_),
    .A2(_07048_),
    .B1(_07047_),
    .X(_07088_));
 sky130_fd_sc_hd__nor2_1 _13938_ (.A(_06826_),
    .B(_06922_),
    .Y(_07089_));
 sky130_fd_sc_hd__inv_2 _13939_ (.A(_06861_),
    .Y(_07090_));
 sky130_fd_sc_hd__a22o_1 _13940_ (.A1(_06844_),
    .A2(_07090_),
    .B1(_06881_),
    .B2(_06923_),
    .X(_07091_));
 sky130_fd_sc_hd__nand4_2 _13941_ (.A(_06844_),
    .B(_07090_),
    .C(_06881_),
    .D(_06923_),
    .Y(_07092_));
 sky130_fd_sc_hd__a21bo_1 _13942_ (.A1(_07089_),
    .A2(_07091_),
    .B1_N(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__and3_1 _13943_ (.A(_07087_),
    .B(_07088_),
    .C(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__a21oi_1 _13944_ (.A1(_07087_),
    .A2(_07088_),
    .B1(_07093_),
    .Y(_07095_));
 sky130_fd_sc_hd__nor2_1 _13945_ (.A(_07094_),
    .B(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__o2bb2a_1 _13946_ (.A1_N(_06895_),
    .A2_N(_06876_),
    .B1(_06884_),
    .B2(_06953_),
    .X(_07097_));
 sky130_fd_sc_hd__a21oi_2 _13947_ (.A1(_07096_),
    .A2(_07097_),
    .B1(_07094_),
    .Y(_07098_));
 sky130_fd_sc_hd__xnor2_2 _13948_ (.A(_07086_),
    .B(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__xnor2_2 _13949_ (.A(_07079_),
    .B(_07073_),
    .Y(_07100_));
 sky130_fd_sc_hd__and2b_1 _13950_ (.A_N(_07098_),
    .B(_07086_),
    .X(_07101_));
 sky130_fd_sc_hd__a21oi_2 _13951_ (.A1(_07099_),
    .A2(_07100_),
    .B1(_07101_),
    .Y(_07102_));
 sky130_fd_sc_hd__xor2_2 _13952_ (.A(_07057_),
    .B(_07058_),
    .X(_07103_));
 sky130_fd_sc_hd__xnor2_2 _13953_ (.A(_07102_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__nand2_1 _13954_ (.A(net3405),
    .B(_07084_),
    .Y(_07105_));
 sky130_fd_sc_hd__xnor2_2 _13955_ (.A(_07081_),
    .B(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__and2b_1 _13956_ (.A_N(_07102_),
    .B(net535),
    .X(_07107_));
 sky130_fd_sc_hd__a21o_1 _13957_ (.A1(net555),
    .A2(net583),
    .B1(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__xnor2_2 _13958_ (.A(_07062_),
    .B(_07064_),
    .Y(_07109_));
 sky130_fd_sc_hd__xor2_2 _13959_ (.A(_07108_),
    .B(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__xnor2_2 _13960_ (.A(_07085_),
    .B(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__xnor2_2 _13961_ (.A(_07076_),
    .B(_07078_),
    .Y(_07112_));
 sky130_fd_sc_hd__nor2_1 _13962_ (.A(_06888_),
    .B(net548),
    .Y(_07113_));
 sky130_fd_sc_hd__xor2_1 _13963_ (.A(_06888_),
    .B(_07112_),
    .X(_07114_));
 sky130_fd_sc_hd__nor2_1 _13964_ (.A(_06865_),
    .B(net541),
    .Y(_07115_));
 sky130_fd_sc_hd__nor2_1 _13965_ (.A(_06862_),
    .B(net564),
    .Y(_07116_));
 sky130_fd_sc_hd__and3_1 _13966_ (.A(_07114_),
    .B(_07115_),
    .C(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__nor2_1 _13967_ (.A(_06862_),
    .B(net573),
    .Y(_07118_));
 sky130_fd_sc_hd__o21a_1 _13968_ (.A1(_07113_),
    .A2(_07117_),
    .B1(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__xnor2_1 _13969_ (.A(_07096_),
    .B(_07097_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand3_1 _13970_ (.A(_07092_),
    .B(_07089_),
    .C(_07091_),
    .Y(_07121_));
 sky130_fd_sc_hd__a21o_1 _13971_ (.A1(_07092_),
    .A2(_07091_),
    .B1(_07089_),
    .X(_07122_));
 sky130_fd_sc_hd__nor2_1 _13972_ (.A(_06885_),
    .B(_06922_),
    .Y(_07123_));
 sky130_fd_sc_hd__o22ai_1 _13973_ (.A1(_06861_),
    .A2(_06837_),
    .B1(_06918_),
    .B2(_06895_),
    .Y(_07124_));
 sky130_fd_sc_hd__and4b_1 _13974_ (.A_N(_06826_),
    .B(_07090_),
    .C(_06881_),
    .D(_06923_),
    .X(_07125_));
 sky130_fd_sc_hd__a21o_1 _13975_ (.A1(_07123_),
    .A2(_07124_),
    .B1(_07125_),
    .X(_07126_));
 sky130_fd_sc_hd__nand3_1 _13976_ (.A(_07121_),
    .B(_07122_),
    .C(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21o_1 _13977_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07126_),
    .X(_07128_));
 sky130_fd_sc_hd__or2_1 _13978_ (.A(_06876_),
    .B(_06970_),
    .X(_07129_));
 sky130_fd_sc_hd__nand2_1 _13979_ (.A(_06876_),
    .B(_06970_),
    .Y(_07130_));
 sky130_fd_sc_hd__nor2_1 _13980_ (.A(_06869_),
    .B(_06990_),
    .Y(_07131_));
 sky130_fd_sc_hd__a41o_1 _13981_ (.A1(_06781_),
    .A2(_06869_),
    .A3(_07129_),
    .A4(_07130_),
    .B1(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand3_1 _13982_ (.A(_07127_),
    .B(_07128_),
    .C(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_1 _13983_ (.A(_07127_),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__xnor2_1 _13984_ (.A(_07120_),
    .B(_07134_),
    .Y(_07135_));
 sky130_fd_sc_hd__nand2_1 _13985_ (.A(_07115_),
    .B(_07116_),
    .Y(_07136_));
 sky130_fd_sc_hd__xnor2_2 _13986_ (.A(net536),
    .B(_07136_),
    .Y(_07137_));
 sky130_fd_sc_hd__and2b_1 _13987_ (.A_N(_07120_),
    .B(_07134_),
    .X(_07138_));
 sky130_fd_sc_hd__a21oi_2 _13988_ (.A1(_07135_),
    .A2(_07137_),
    .B1(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__xnor2_2 _13989_ (.A(_07099_),
    .B(_07100_),
    .Y(_07140_));
 sky130_fd_sc_hd__xor2_1 _13990_ (.A(_07139_),
    .B(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__or3_4 _13991_ (.A(_07113_),
    .B(_07117_),
    .C(_07118_),
    .X(_07142_));
 sky130_fd_sc_hd__and2b_1 _13992_ (.A_N(_07119_),
    .B(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__nor2_1 _13993_ (.A(_07139_),
    .B(_07140_),
    .Y(_07144_));
 sky130_fd_sc_hd__a21oi_2 _13994_ (.A1(_07141_),
    .A2(_07143_),
    .B1(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__xor2_2 _13995_ (.A(_07104_),
    .B(_07106_),
    .X(_07146_));
 sky130_fd_sc_hd__xnor2_2 _13996_ (.A(_07145_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__or2b_1 _13997_ (.A(net3163),
    .B_N(_07146_),
    .X(_07148_));
 sky130_fd_sc_hd__a21boi_2 _13998_ (.A1(_07119_),
    .A2(_07147_),
    .B1_N(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_1 _13999_ (.A(_07111_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__xnor2_2 _14000_ (.A(_07041_),
    .B(_07068_),
    .Y(_07151_));
 sky130_fd_sc_hd__and2_1 _14001_ (.A(_07085_),
    .B(net75),
    .X(_07152_));
 sky130_fd_sc_hd__a21oi_2 _14002_ (.A1(_07108_),
    .A2(net550),
    .B1(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__xnor2_2 _14003_ (.A(_07151_),
    .B(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__nand2_1 _14004_ (.A(_07150_),
    .B(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__xor2_1 _14005_ (.A(_07119_),
    .B(_07147_),
    .X(_07156_));
 sky130_fd_sc_hd__xnor2_1 _14006_ (.A(_07115_),
    .B(_07116_),
    .Y(_07157_));
 sky130_fd_sc_hd__nor2_1 _14007_ (.A(_06865_),
    .B(_06990_),
    .Y(_07158_));
 sky130_fd_sc_hd__nor2_1 _14008_ (.A(_06781_),
    .B(_06876_),
    .Y(_07159_));
 sky130_fd_sc_hd__mux2_1 _14009_ (.A0(_06970_),
    .A1(_07159_),
    .S(_06869_),
    .X(_07160_));
 sky130_fd_sc_hd__or3_1 _14010_ (.A(_06876_),
    .B(_06869_),
    .C(_06970_),
    .X(_07161_));
 sky130_fd_sc_hd__a21bo_1 _14011_ (.A1(_07158_),
    .A2(_07160_),
    .B1_N(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__nand2b_1 _14012_ (.A_N(_07157_),
    .B(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__or2b_1 _14013_ (.A(_07162_),
    .B_N(_07157_),
    .X(_07164_));
 sky130_fd_sc_hd__nand2_1 _14014_ (.A(_07163_),
    .B(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__a21o_1 _14015_ (.A1(_07127_),
    .A2(_07128_),
    .B1(_07132_),
    .X(_07166_));
 sky130_fd_sc_hd__or2b_1 _14016_ (.A(_07125_),
    .B_N(_07124_),
    .X(_07167_));
 sky130_fd_sc_hd__xnor2_1 _14017_ (.A(_07123_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__nor2_1 _14018_ (.A(net552),
    .B(_06922_),
    .Y(_07169_));
 sky130_fd_sc_hd__o22ai_2 _14019_ (.A1(_06895_),
    .A2(_06861_),
    .B1(_06885_),
    .B2(_06918_),
    .Y(_07170_));
 sky130_fd_sc_hd__or4_1 _14020_ (.A(_06826_),
    .B(_06861_),
    .C(_06864_),
    .D(_06885_),
    .X(_07171_));
 sky130_fd_sc_hd__a21bo_1 _14021_ (.A1(_07169_),
    .A2(_07170_),
    .B1_N(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__xnor2_1 _14022_ (.A(_07158_),
    .B(_07160_),
    .Y(_07173_));
 sky130_fd_sc_hd__xnor2_1 _14023_ (.A(_07168_),
    .B(_07172_),
    .Y(_07174_));
 sky130_fd_sc_hd__nor2_1 _14024_ (.A(_07173_),
    .B(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__a21o_1 _14025_ (.A1(_07168_),
    .A2(_07172_),
    .B1(_07175_),
    .X(_07176_));
 sky130_fd_sc_hd__a21oi_1 _14026_ (.A1(_07133_),
    .A2(_07166_),
    .B1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__and3_1 _14027_ (.A(_07133_),
    .B(_07166_),
    .C(_07176_),
    .X(_07178_));
 sky130_fd_sc_hd__o21bai_1 _14028_ (.A1(_07165_),
    .A2(_07177_),
    .B1_N(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__xor2_1 _14029_ (.A(_07135_),
    .B(net551),
    .X(_07180_));
 sky130_fd_sc_hd__nor2_1 _14030_ (.A(_07179_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__and2_1 _14031_ (.A(_07179_),
    .B(_07180_),
    .X(_07182_));
 sky130_fd_sc_hd__o21ba_1 _14032_ (.A1(_07163_),
    .A2(_07181_),
    .B1_N(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__xor2_1 _14033_ (.A(net537),
    .B(_07143_),
    .X(_07184_));
 sky130_fd_sc_hd__and2b_1 _14034_ (.A_N(_07183_),
    .B(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__xor2_1 _14035_ (.A(_07111_),
    .B(_07149_),
    .X(_07186_));
 sky130_fd_sc_hd__and3_1 _14036_ (.A(net528),
    .B(_07185_),
    .C(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__nand2_1 _14037_ (.A(net528),
    .B(_07185_),
    .Y(_07188_));
 sky130_fd_sc_hd__xnor2_1 _14038_ (.A(_07188_),
    .B(_07186_),
    .Y(_07189_));
 sky130_fd_sc_hd__and2b_1 _14039_ (.A_N(_07184_),
    .B(_07183_),
    .X(_07190_));
 sky130_fd_sc_hd__or3b_4 _14040_ (.A(_07185_),
    .B(_07190_),
    .C_N(_07156_),
    .X(_07191_));
 sky130_fd_sc_hd__nor2_1 _14041_ (.A(_06862_),
    .B(net542),
    .Y(_07192_));
 sky130_fd_sc_hd__or2_1 _14042_ (.A(_06819_),
    .B(_06869_),
    .X(_07193_));
 sky130_fd_sc_hd__or3_1 _14043_ (.A(_06864_),
    .B(_07193_),
    .C(_06970_),
    .X(_07194_));
 sky130_fd_sc_hd__o21ai_1 _14044_ (.A1(_06865_),
    .A2(_06955_),
    .B1(_07193_),
    .Y(_07195_));
 sky130_fd_sc_hd__nand2_1 _14045_ (.A(_07194_),
    .B(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__o31ai_1 _14046_ (.A1(_06862_),
    .A2(_06990_),
    .A3(_07196_),
    .B1(_07194_),
    .Y(_07197_));
 sky130_fd_sc_hd__and2_1 _14047_ (.A(_07192_),
    .B(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__and3_1 _14048_ (.A(_07171_),
    .B(_07169_),
    .C(_07170_),
    .X(_07199_));
 sky130_fd_sc_hd__a21oi_1 _14049_ (.A1(_07171_),
    .A2(_07170_),
    .B1(_07169_),
    .Y(_07200_));
 sky130_fd_sc_hd__or2_1 _14050_ (.A(_07199_),
    .B(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__or2_1 _14051_ (.A(_06861_),
    .B(_06885_),
    .X(_07202_));
 sky130_fd_sc_hd__or2_1 _14052_ (.A(net552),
    .B(_06918_),
    .X(_07203_));
 sky130_fd_sc_hd__nand2_1 _14053_ (.A(_07202_),
    .B(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_06862_),
    .B(_06864_),
    .Y(_07205_));
 sky130_fd_sc_hd__nor2_1 _14055_ (.A(_07205_),
    .B(_06869_),
    .Y(_07206_));
 sky130_fd_sc_hd__nor2_1 _14056_ (.A(_07202_),
    .B(_07203_),
    .Y(_07207_));
 sky130_fd_sc_hd__a21oi_1 _14057_ (.A1(_07204_),
    .A2(_07206_),
    .B1(_07207_),
    .Y(_07208_));
 sky130_fd_sc_hd__nor2_1 _14058_ (.A(_07201_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__nor2_1 _14059_ (.A(_06862_),
    .B(_06990_),
    .Y(_07210_));
 sky130_fd_sc_hd__xnor2_1 _14060_ (.A(_07196_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__and2_1 _14061_ (.A(_07201_),
    .B(_07208_),
    .X(_07212_));
 sky130_fd_sc_hd__nor2_1 _14062_ (.A(_07209_),
    .B(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__and2_1 _14063_ (.A(_07211_),
    .B(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__and2_1 _14064_ (.A(_07173_),
    .B(_07174_),
    .X(_07215_));
 sky130_fd_sc_hd__nor2_1 _14065_ (.A(_07175_),
    .B(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__o21a_1 _14066_ (.A1(_07209_),
    .A2(_07214_),
    .B1(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__xnor2_1 _14067_ (.A(_07192_),
    .B(_07197_),
    .Y(_07218_));
 sky130_fd_sc_hd__nor3_1 _14068_ (.A(_07216_),
    .B(_07209_),
    .C(_07214_),
    .Y(_07219_));
 sky130_fd_sc_hd__or2_1 _14069_ (.A(_07217_),
    .B(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__nor2_1 _14070_ (.A(_07218_),
    .B(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__nor2_1 _14071_ (.A(_07178_),
    .B(_07177_),
    .Y(_07222_));
 sky130_fd_sc_hd__xnor2_1 _14072_ (.A(_07165_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__o21a_1 _14073_ (.A1(_07217_),
    .A2(_07221_),
    .B1(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__or3_1 _14074_ (.A(_07223_),
    .B(_07217_),
    .C(_07221_),
    .X(_07225_));
 sky130_fd_sc_hd__and2b_1 _14075_ (.A_N(_07224_),
    .B(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__a21o_1 _14076_ (.A1(_07198_),
    .A2(_07226_),
    .B1(_07224_),
    .X(_07227_));
 sky130_fd_sc_hd__nor2_1 _14077_ (.A(_07182_),
    .B(_07181_),
    .Y(_07228_));
 sky130_fd_sc_hd__xnor2_1 _14078_ (.A(_07163_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__and3b_1 _14079_ (.A_N(_07191_),
    .B(_07227_),
    .C(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__xnor2_2 _14080_ (.A(_07189_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__buf_2 _14081_ (.A(_06862_),
    .X(_07232_));
 sky130_fd_sc_hd__nor2_1 _14082_ (.A(_07211_),
    .B(_07213_),
    .Y(_07233_));
 sky130_fd_sc_hd__or2_1 _14083_ (.A(_07214_),
    .B(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__o22a_1 _14084_ (.A1(_06865_),
    .A2(_06957_),
    .B1(_06955_),
    .B2(_07232_),
    .X(_07235_));
 sky130_fd_sc_hd__or2_1 _14085_ (.A(_07207_),
    .B(_07235_),
    .X(_07236_));
 sky130_fd_sc_hd__o21a_1 _14086_ (.A1(_07204_),
    .A2(_07206_),
    .B1(_07208_),
    .X(_07237_));
 sky130_fd_sc_hd__nor2_1 _14087_ (.A(_07159_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__or3_1 _14088_ (.A(_07234_),
    .B(_07236_),
    .C(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__o21ai_1 _14089_ (.A1(_07236_),
    .A2(_07238_),
    .B1(_07234_),
    .Y(_07240_));
 sky130_fd_sc_hd__and2_1 _14090_ (.A(_07239_),
    .B(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__a2bb2o_1 _14091_ (.A1_N(_07207_),
    .A2_N(_07241_),
    .B1(_06865_),
    .B2(_07193_),
    .X(_07242_));
 sky130_fd_sc_hd__nand2_1 _14092_ (.A(_07218_),
    .B(_07220_),
    .Y(_07243_));
 sky130_fd_sc_hd__or2b_1 _14093_ (.A(_07221_),
    .B_N(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__o21a_1 _14094_ (.A1(_07232_),
    .A2(_07242_),
    .B1(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__nand2_1 _14095_ (.A(_07159_),
    .B(_06970_),
    .Y(_07246_));
 sky130_fd_sc_hd__a2bb2o_1 _14096_ (.A1_N(_07198_),
    .A2_N(_07226_),
    .B1(_07246_),
    .B2(_07239_),
    .X(_07247_));
 sky130_fd_sc_hd__nor2_1 _14097_ (.A(_07227_),
    .B(_07229_),
    .Y(_07248_));
 sky130_fd_sc_hd__or4_4 _14098_ (.A(_07191_),
    .B(_07245_),
    .C(_07247_),
    .D(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__and2_1 _14099_ (.A(_07189_),
    .B(_07230_),
    .X(_07250_));
 sky130_fd_sc_hd__o21bai_4 _14100_ (.A1(_07231_),
    .A2(_07249_),
    .B1_N(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__or2_4 _14101_ (.A(_07150_),
    .B(_07187_),
    .X(_07252_));
 sky130_fd_sc_hd__xor2_2 _14102_ (.A(_07154_),
    .B(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__a22o_4 _14103_ (.A1(_07154_),
    .A2(_07187_),
    .B1(_07251_),
    .B2(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__or2b_1 _14104_ (.A(_07153_),
    .B_N(_07151_),
    .X(_07255_));
 sky130_fd_sc_hd__nand2_1 _14105_ (.A(_07255_),
    .B(_07155_),
    .Y(_07256_));
 sky130_fd_sc_hd__xnor2_1 _14106_ (.A(_07071_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__a2bb2o_4 _14107_ (.A1_N(_07071_),
    .A2_N(_07155_),
    .B1(_07254_),
    .B2(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__or2_1 _14108_ (.A(_07011_),
    .B(_07020_),
    .X(_07259_));
 sky130_fd_sc_hd__a21bo_1 _14109_ (.A1(_07013_),
    .A2(_07019_),
    .B1_N(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__nor2_1 _14110_ (.A(_07010_),
    .B(_07021_),
    .Y(_07261_));
 sky130_fd_sc_hd__or2_1 _14111_ (.A(_06992_),
    .B(_06994_),
    .X(_07262_));
 sky130_fd_sc_hd__nand2_1 _14112_ (.A(_06995_),
    .B(_07006_),
    .Y(_07263_));
 sky130_fd_sc_hd__nor2_1 _14113_ (.A(_06668_),
    .B(_06955_),
    .Y(_07264_));
 sky130_fd_sc_hd__nor2_1 _14114_ (.A(_06737_),
    .B(_06990_),
    .Y(_07265_));
 sky130_fd_sc_hd__xor2_1 _14115_ (.A(_07264_),
    .B(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__a2bb2o_1 _14116_ (.A1_N(_06957_),
    .A2_N(_06987_),
    .B1(_06988_),
    .B2(_06991_),
    .X(_07267_));
 sky130_fd_sc_hd__inv_2 _14117_ (.A(net542),
    .Y(_07268_));
 sky130_fd_sc_hd__o22a_1 _14118_ (.A1(_06881_),
    .A2(net531),
    .B1(_07268_),
    .B2(_06931_),
    .X(_07269_));
 sky130_fd_sc_hd__xor2_1 _14119_ (.A(_07267_),
    .B(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__a21oi_1 _14120_ (.A1(_06889_),
    .A2(_06931_),
    .B1(_06846_),
    .Y(_07271_));
 sky130_fd_sc_hd__xor2_1 _14121_ (.A(_07270_),
    .B(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_07266_),
    .B(_07272_),
    .Y(_07273_));
 sky130_fd_sc_hd__a21o_1 _14123_ (.A1(_07262_),
    .A2(_07263_),
    .B1(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__nand3_1 _14124_ (.A(_07262_),
    .B(_07263_),
    .C(_07273_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand2_1 _14125_ (.A(_07274_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__or2b_1 _14126_ (.A(_07014_),
    .B_N(_07018_),
    .X(_07277_));
 sky130_fd_sc_hd__and2b_1 _14127_ (.A_N(_06997_),
    .B(_07005_),
    .X(_07278_));
 sky130_fd_sc_hd__or2_1 _14128_ (.A(_07003_),
    .B(_07278_),
    .X(_07279_));
 sky130_fd_sc_hd__or2_1 _14129_ (.A(_06970_),
    .B(_06867_),
    .X(_07280_));
 sky130_fd_sc_hd__or3_1 _14130_ (.A(_06895_),
    .B(_06858_),
    .C(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__o21ai_1 _14131_ (.A1(_06895_),
    .A2(_06858_),
    .B1(_07280_),
    .Y(_07282_));
 sky130_fd_sc_hd__and2_1 _14132_ (.A(_07281_),
    .B(_07282_),
    .X(_07283_));
 sky130_fd_sc_hd__xnor2_1 _14133_ (.A(_07016_),
    .B(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__xnor2_1 _14134_ (.A(_07279_),
    .B(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__xnor2_1 _14135_ (.A(_07277_),
    .B(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__xor2_1 _14136_ (.A(_07276_),
    .B(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__o21ai_2 _14137_ (.A1(_07008_),
    .A2(_07261_),
    .B1(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__or3_1 _14138_ (.A(_07008_),
    .B(_07261_),
    .C(_07287_),
    .X(_07289_));
 sky130_fd_sc_hd__and2_1 _14139_ (.A(_07288_),
    .B(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__xnor2_1 _14140_ (.A(_07260_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__or2b_1 _14141_ (.A(_07023_),
    .B_N(_06913_),
    .X(_07292_));
 sky130_fd_sc_hd__a21boi_1 _14142_ (.A1(_06985_),
    .A2(_07022_),
    .B1_N(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__nor2_2 _14143_ (.A(_07291_),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__and2_1 _14144_ (.A(_07291_),
    .B(_07293_),
    .X(_07295_));
 sky130_fd_sc_hd__nor2_4 _14145_ (.A(_07294_),
    .B(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__and2b_1 _14146_ (.A_N(_07070_),
    .B(_07024_),
    .X(_07297_));
 sky130_fd_sc_hd__nor2_1 _14147_ (.A(_07071_),
    .B(_07255_),
    .Y(_07298_));
 sky130_fd_sc_hd__nor2_1 _14148_ (.A(_07297_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__xnor2_2 _14149_ (.A(_07296_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__xnor2_2 _14150_ (.A(_07258_),
    .B(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__xor2_1 _14151_ (.A(_07254_),
    .B(_07257_),
    .X(_07302_));
 sky130_fd_sc_hd__xnor2_1 _14152_ (.A(_07251_),
    .B(_07253_),
    .Y(_07303_));
 sky130_fd_sc_hd__xnor2_4 _14153_ (.A(net559),
    .B(net560),
    .Y(_07304_));
 sky130_fd_sc_hd__nor2_1 _14154_ (.A(_07303_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_07302_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__nand2_1 _14156_ (.A(_07301_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__nand2_1 _14157_ (.A(_07260_),
    .B(_07290_),
    .Y(_07308_));
 sky130_fd_sc_hd__or2_1 _14158_ (.A(_07276_),
    .B(_07286_),
    .X(_07309_));
 sky130_fd_sc_hd__nand2_1 _14159_ (.A(_07266_),
    .B(_07272_),
    .Y(_07310_));
 sky130_fd_sc_hd__buf_2 _14160_ (.A(_06668_),
    .X(_07311_));
 sky130_fd_sc_hd__or2_1 _14161_ (.A(_07311_),
    .B(_06990_),
    .X(_07312_));
 sky130_fd_sc_hd__nand2_1 _14162_ (.A(_07264_),
    .B(_07265_),
    .Y(_07313_));
 sky130_fd_sc_hd__nand2_1 _14163_ (.A(_06880_),
    .B(_07000_),
    .Y(_07314_));
 sky130_fd_sc_hd__and4bb_1 _14164_ (.A_N(_06931_),
    .B_N(_06973_),
    .C(_07268_),
    .D(_06866_),
    .X(_07315_));
 sky130_fd_sc_hd__o22a_1 _14165_ (.A1(_06737_),
    .A2(net545),
    .B1(_06973_),
    .B2(_06931_),
    .X(_07316_));
 sky130_fd_sc_hd__nor2_1 _14166_ (.A(_07315_),
    .B(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__xnor2_1 _14167_ (.A(_07314_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__xnor2_1 _14168_ (.A(_07313_),
    .B(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__xnor2_1 _14169_ (.A(net568),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__xnor2_1 _14170_ (.A(_07312_),
    .B(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nor2_1 _14171_ (.A(_07310_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__and2_1 _14172_ (.A(_07310_),
    .B(_07321_),
    .X(_07323_));
 sky130_fd_sc_hd__or2_1 _14173_ (.A(_07322_),
    .B(_07323_),
    .X(_07324_));
 sky130_fd_sc_hd__and2b_1 _14174_ (.A_N(_07016_),
    .B(_07283_),
    .X(_07325_));
 sky130_fd_sc_hd__and2_1 _14175_ (.A(_07267_),
    .B(_07269_),
    .X(_07326_));
 sky130_fd_sc_hd__and2_1 _14176_ (.A(_07270_),
    .B(_07271_),
    .X(_07327_));
 sky130_fd_sc_hd__or2_1 _14177_ (.A(_06895_),
    .B(_06867_),
    .X(_07328_));
 sky130_fd_sc_hd__nand2_1 _14178_ (.A(_06881_),
    .B(_07082_),
    .Y(_07329_));
 sky130_fd_sc_hd__xor2_1 _14179_ (.A(_07328_),
    .B(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__xnor2_1 _14180_ (.A(_07281_),
    .B(_07330_),
    .Y(_07331_));
 sky130_fd_sc_hd__o21a_1 _14181_ (.A1(_07326_),
    .A2(_07327_),
    .B1(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__nor3_1 _14182_ (.A(_07326_),
    .B(_07327_),
    .C(_07331_),
    .Y(_07333_));
 sky130_fd_sc_hd__nor2_1 _14183_ (.A(_07332_),
    .B(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__xnor2_1 _14184_ (.A(_07325_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__xnor2_1 _14185_ (.A(_07324_),
    .B(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__a21o_1 _14186_ (.A1(_07274_),
    .A2(_07309_),
    .B1(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__nand3_1 _14187_ (.A(_07274_),
    .B(_07309_),
    .C(_07336_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_1 _14188_ (.A(_07337_),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__nand2_1 _14189_ (.A(_07279_),
    .B(_07284_),
    .Y(_07340_));
 sky130_fd_sc_hd__o21a_1 _14190_ (.A1(_07277_),
    .A2(_07285_),
    .B1(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__xnor2_1 _14191_ (.A(_07339_),
    .B(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__a21oi_2 _14192_ (.A1(_07288_),
    .A2(_07308_),
    .B1(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__and3_1 _14193_ (.A(_07288_),
    .B(_07308_),
    .C(_07342_),
    .X(_07344_));
 sky130_fd_sc_hd__or2_1 _14194_ (.A(_07343_),
    .B(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__inv_2 _14195_ (.A(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__a21oi_1 _14196_ (.A1(_07297_),
    .A2(_07296_),
    .B1(_07294_),
    .Y(_07347_));
 sky130_fd_sc_hd__xnor2_1 _14197_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__a22o_1 _14198_ (.A1(_07296_),
    .A2(_07298_),
    .B1(_07300_),
    .B2(_07258_),
    .X(_07349_));
 sky130_fd_sc_hd__xor2_1 _14199_ (.A(_07348_),
    .B(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__or2_4 _14200_ (.A(_07307_),
    .B(_07350_),
    .X(_07351_));
 sky130_fd_sc_hd__nand2_1 _14201_ (.A(_07307_),
    .B(_07350_),
    .Y(_07352_));
 sky130_fd_sc_hd__nand2_2 _14202_ (.A(_07351_),
    .B(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__buf_2 _14203_ (.A(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__or2_1 _14204_ (.A(_06859_),
    .B(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__clkbuf_4 _14205_ (.A(_06867_),
    .X(_07356_));
 sky130_fd_sc_hd__or2_1 _14206_ (.A(_07301_),
    .B(_07306_),
    .X(_07357_));
 sky130_fd_sc_hd__nand2_2 _14207_ (.A(_07307_),
    .B(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__clkbuf_4 _14208_ (.A(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__nor2_1 _14209_ (.A(_07356_),
    .B(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__and2b_1 _14210_ (.A_N(_07355_),
    .B(_07360_),
    .X(_07361_));
 sky130_fd_sc_hd__a32o_2 _14211_ (.A1(_07297_),
    .A2(_07296_),
    .A3(_07346_),
    .B1(_07348_),
    .B2(_07349_),
    .X(_07362_));
 sky130_fd_sc_hd__or2_1 _14212_ (.A(_07339_),
    .B(_07341_),
    .X(_07363_));
 sky130_fd_sc_hd__nor2_1 _14213_ (.A(_07324_),
    .B(_07335_),
    .Y(_07364_));
 sky130_fd_sc_hd__nor2_1 _14214_ (.A(_07312_),
    .B(_07320_),
    .Y(_07365_));
 sky130_fd_sc_hd__clkbuf_4 _14215_ (.A(_06973_),
    .X(_07366_));
 sky130_fd_sc_hd__buf_2 _14216_ (.A(net544),
    .X(_07367_));
 sky130_fd_sc_hd__o21ai_1 _14217_ (.A1(_06737_),
    .A2(_07366_),
    .B1(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__or3_1 _14218_ (.A(_06737_),
    .B(net543),
    .C(_07366_),
    .X(_07369_));
 sky130_fd_sc_hd__and2_1 _14219_ (.A(_07368_),
    .B(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__nand2_1 _14220_ (.A(_07365_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__or2_1 _14221_ (.A(_07365_),
    .B(_07370_),
    .X(_07372_));
 sky130_fd_sc_hd__nand2_1 _14222_ (.A(_07371_),
    .B(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__or2b_1 _14223_ (.A(_07281_),
    .B_N(_07330_),
    .X(_07374_));
 sky130_fd_sc_hd__a32o_1 _14224_ (.A1(_07264_),
    .A2(_07265_),
    .A3(_07318_),
    .B1(_07319_),
    .B2(net568),
    .X(_07375_));
 sky130_fd_sc_hd__or2_1 _14225_ (.A(_07328_),
    .B(_07329_),
    .X(_07376_));
 sky130_fd_sc_hd__or2_1 _14226_ (.A(_06837_),
    .B(_06867_),
    .X(_07377_));
 sky130_fd_sc_hd__nand2_1 _14227_ (.A(_06880_),
    .B(_07082_),
    .Y(_07378_));
 sky130_fd_sc_hd__xor2_1 _14228_ (.A(_07377_),
    .B(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__xnor2_1 _14229_ (.A(_07376_),
    .B(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__nand2_1 _14230_ (.A(_07375_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__or2_1 _14231_ (.A(_07375_),
    .B(_07380_),
    .X(_07382_));
 sky130_fd_sc_hd__nand2_1 _14232_ (.A(_07381_),
    .B(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__xor2_1 _14233_ (.A(_07374_),
    .B(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__xnor2_1 _14234_ (.A(_07373_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__o21ai_1 _14235_ (.A1(_07322_),
    .A2(_07364_),
    .B1(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__or3_1 _14236_ (.A(_07322_),
    .B(_07364_),
    .C(_07385_),
    .X(_07387_));
 sky130_fd_sc_hd__nand2_1 _14237_ (.A(_07386_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__a21oi_2 _14238_ (.A1(_07325_),
    .A2(_07334_),
    .B1(_07332_),
    .Y(_07389_));
 sky130_fd_sc_hd__xnor2_2 _14239_ (.A(_07388_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__a21oi_4 _14240_ (.A1(_07337_),
    .A2(_07363_),
    .B1(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__and3_1 _14241_ (.A(_07337_),
    .B(_07363_),
    .C(_07390_),
    .X(_07392_));
 sky130_fd_sc_hd__nor2_1 _14242_ (.A(_07391_),
    .B(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__xor2_1 _14243_ (.A(_07343_),
    .B(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__nand3_1 _14244_ (.A(_07294_),
    .B(_07346_),
    .C(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__a21o_1 _14245_ (.A1(_07294_),
    .A2(_07346_),
    .B1(_07394_),
    .X(_07396_));
 sky130_fd_sc_hd__and2_2 _14246_ (.A(_07395_),
    .B(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__xor2_4 _14247_ (.A(_07362_),
    .B(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__xnor2_2 _14248_ (.A(_07351_),
    .B(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__clkbuf_4 _14249_ (.A(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__or2_1 _14250_ (.A(_06859_),
    .B(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__nor2_1 _14251_ (.A(_07356_),
    .B(_07354_),
    .Y(_07402_));
 sky130_fd_sc_hd__xnor2_1 _14252_ (.A(_07401_),
    .B(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__or3_1 _14253_ (.A(_07356_),
    .B(_07354_),
    .C(_07401_),
    .X(_07404_));
 sky130_fd_sc_hd__nor2_8 _14254_ (.A(_07351_),
    .B(_07398_),
    .Y(_07405_));
 sky130_fd_sc_hd__a21boi_4 _14255_ (.A1(_07362_),
    .A2(_07397_),
    .B1_N(_07395_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand2_2 _14256_ (.A(_07343_),
    .B(_07393_),
    .Y(_07407_));
 sky130_fd_sc_hd__or2_1 _14257_ (.A(_07388_),
    .B(_07389_),
    .X(_07408_));
 sky130_fd_sc_hd__or2b_1 _14258_ (.A(_07373_),
    .B_N(_07384_),
    .X(_07409_));
 sky130_fd_sc_hd__nand2_1 _14259_ (.A(net569),
    .B(_07370_),
    .Y(_07410_));
 sky130_fd_sc_hd__or4_1 _14260_ (.A(_07311_),
    .B(_06737_),
    .C(net532),
    .D(_07366_),
    .X(_07411_));
 sky130_fd_sc_hd__o22ai_1 _14261_ (.A1(_06737_),
    .A2(net533),
    .B1(_07366_),
    .B2(_07311_),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_1 _14262_ (.A(_07411_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__a21o_1 _14263_ (.A1(_07369_),
    .A2(_07410_),
    .B1(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__nand3_1 _14264_ (.A(_07369_),
    .B(_07410_),
    .C(_07413_),
    .Y(_07415_));
 sky130_fd_sc_hd__nand2_1 _14265_ (.A(_07414_),
    .B(_07415_),
    .Y(_07416_));
 sky130_fd_sc_hd__or2b_1 _14266_ (.A(_07376_),
    .B_N(_07379_),
    .X(_07417_));
 sky130_fd_sc_hd__or2_1 _14267_ (.A(_07377_),
    .B(_07378_),
    .X(_07418_));
 sky130_fd_sc_hd__and2b_1 _14268_ (.A_N(_06867_),
    .B(_06880_),
    .X(_07419_));
 sky130_fd_sc_hd__or2_1 _14269_ (.A(_06931_),
    .B(_06859_),
    .X(_07420_));
 sky130_fd_sc_hd__xnor2_1 _14270_ (.A(_07419_),
    .B(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__nand2_1 _14271_ (.A(net569),
    .B(_07410_),
    .Y(_07422_));
 sky130_fd_sc_hd__and3_1 _14272_ (.A(_07418_),
    .B(_07421_),
    .C(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__xnor2_1 _14273_ (.A(_07417_),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__xor2_1 _14274_ (.A(_07416_),
    .B(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__a21oi_1 _14275_ (.A1(_07371_),
    .A2(_07409_),
    .B1(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__and3_1 _14276_ (.A(_07371_),
    .B(_07409_),
    .C(_07425_),
    .X(_07427_));
 sky130_fd_sc_hd__nor2_1 _14277_ (.A(_07426_),
    .B(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__o21a_1 _14278_ (.A1(_07374_),
    .A2(_07383_),
    .B1(_07381_),
    .X(_07429_));
 sky130_fd_sc_hd__inv_2 _14279_ (.A(_07429_),
    .Y(_07430_));
 sky130_fd_sc_hd__xnor2_1 _14280_ (.A(_07428_),
    .B(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__a21o_1 _14281_ (.A1(_07386_),
    .A2(_07408_),
    .B1(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__nand3_1 _14282_ (.A(_07386_),
    .B(_07408_),
    .C(_07431_),
    .Y(_07433_));
 sky130_fd_sc_hd__and2_2 _14283_ (.A(_07432_),
    .B(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__xnor2_4 _14284_ (.A(_07391_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__xnor2_4 _14285_ (.A(_07407_),
    .B(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__xnor2_4 _14286_ (.A(_07406_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__xnor2_4 _14287_ (.A(_07405_),
    .B(_07437_),
    .Y(_07438_));
 sky130_fd_sc_hd__buf_6 _14288_ (.A(_07438_),
    .X(_07439_));
 sky130_fd_sc_hd__or2_1 _14289_ (.A(_06859_),
    .B(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__nor2_1 _14290_ (.A(_07356_),
    .B(_07400_),
    .Y(_07441_));
 sky130_fd_sc_hd__xnor2_1 _14291_ (.A(_07440_),
    .B(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__xnor2_1 _14292_ (.A(_07404_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__clkbuf_4 _14293_ (.A(_06990_),
    .X(_07444_));
 sky130_fd_sc_hd__nand2_1 _14294_ (.A(_07362_),
    .B(_07397_),
    .Y(_07445_));
 sky130_fd_sc_hd__a21oi_1 _14295_ (.A1(_07428_),
    .A2(_07430_),
    .B1(_07426_),
    .Y(_07446_));
 sky130_fd_sc_hd__or2b_1 _14296_ (.A(_07416_),
    .B_N(_07424_),
    .X(_07447_));
 sky130_fd_sc_hd__o211a_1 _14297_ (.A1(_06737_),
    .A2(_07366_),
    .B1(_07000_),
    .C1(_06611_),
    .X(_07448_));
 sky130_fd_sc_hd__a21o_1 _14298_ (.A1(_07082_),
    .A2(_07419_),
    .B1(_06931_),
    .X(_07449_));
 sky130_fd_sc_hd__nor2_1 _14299_ (.A(_07414_),
    .B(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__and2_1 _14300_ (.A(_07414_),
    .B(_07449_),
    .X(_07451_));
 sky130_fd_sc_hd__o21ai_1 _14301_ (.A1(_07450_),
    .A2(_07451_),
    .B1(_07418_),
    .Y(_07452_));
 sky130_fd_sc_hd__xor2_1 _14302_ (.A(_07448_),
    .B(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__xnor2_1 _14303_ (.A(_07447_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__inv_2 _14304_ (.A(_07423_),
    .Y(_07455_));
 sky130_fd_sc_hd__o21a_1 _14305_ (.A1(_07417_),
    .A2(_07455_),
    .B1(_07422_),
    .X(_07456_));
 sky130_fd_sc_hd__xnor2_1 _14306_ (.A(_07454_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__xnor2_1 _14307_ (.A(_07446_),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__xnor2_1 _14308_ (.A(_07432_),
    .B(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__a21oi_1 _14309_ (.A1(_07407_),
    .A2(_07395_),
    .B1(_07435_),
    .Y(_07460_));
 sky130_fd_sc_hd__a21oi_1 _14310_ (.A1(_07391_),
    .A2(_07434_),
    .B1(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__o211a_1 _14311_ (.A1(_07445_),
    .A2(_07436_),
    .B1(_07459_),
    .C1(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__a21o_1 _14312_ (.A1(_07405_),
    .A2(_07437_),
    .B1(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__buf_6 _14313_ (.A(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__nor2_2 _14314_ (.A(_07444_),
    .B(net558),
    .Y(_07465_));
 sky130_fd_sc_hd__a21oi_2 _14315_ (.A1(_07405_),
    .A2(_07437_),
    .B1(_07462_),
    .Y(_07466_));
 sky130_fd_sc_hd__clkbuf_4 _14316_ (.A(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__nor2_2 _14317_ (.A(_07311_),
    .B(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__a22o_1 _14318_ (.A1(net3246),
    .A2(_07467_),
    .B1(_07468_),
    .B2(net586),
    .X(_07469_));
 sky130_fd_sc_hd__nand2_2 _14319_ (.A(_07268_),
    .B(_07467_),
    .Y(_07470_));
 sky130_fd_sc_hd__clkbuf_4 _14320_ (.A(_07366_),
    .X(_07471_));
 sky130_fd_sc_hd__nor2_1 _14321_ (.A(_07471_),
    .B(_07464_),
    .Y(_07472_));
 sky130_fd_sc_hd__xnor2_2 _14322_ (.A(_07470_),
    .B(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__clkbuf_4 _14323_ (.A(net534),
    .X(_07474_));
 sky130_fd_sc_hd__nor2_1 _14324_ (.A(_07474_),
    .B(_07439_),
    .Y(_07475_));
 sky130_fd_sc_hd__xor2_1 _14325_ (.A(_07473_),
    .B(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__nand2_1 _14326_ (.A(_07465_),
    .B(_07469_),
    .Y(_07477_));
 sky130_fd_sc_hd__xor2_1 _14327_ (.A(_07477_),
    .B(_07476_),
    .X(_07478_));
 sky130_fd_sc_hd__nor2_1 _14328_ (.A(_07367_),
    .B(net558),
    .Y(_07479_));
 sky130_fd_sc_hd__nor2_1 _14329_ (.A(_07471_),
    .B(_07439_),
    .Y(_07480_));
 sky130_fd_sc_hd__nor2_1 _14330_ (.A(_07474_),
    .B(_07400_),
    .Y(_07481_));
 sky130_fd_sc_hd__xnor2_1 _14331_ (.A(_07470_),
    .B(_07480_),
    .Y(_07482_));
 sky130_fd_sc_hd__and2_1 _14332_ (.A(_07481_),
    .B(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__a21oi_1 _14333_ (.A1(_07479_),
    .A2(_07480_),
    .B1(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__nor2_1 _14334_ (.A(_07478_),
    .B(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__a31o_1 _14335_ (.A1(_07465_),
    .A2(_07469_),
    .A3(_07476_),
    .B1(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__xor2_1 _14336_ (.A(_07443_),
    .B(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__a32o_1 _14337_ (.A1(_07361_),
    .A2(_07403_),
    .A3(_07487_),
    .B1(_07486_),
    .B2(_07443_),
    .X(_07488_));
 sky130_fd_sc_hd__nor2_1 _14338_ (.A(_07474_),
    .B(net558),
    .Y(_07489_));
 sky130_fd_sc_hd__a211o_1 _14339_ (.A1(_07268_),
    .A2(_07468_),
    .B1(_07472_),
    .C1(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__nand2_1 _14340_ (.A(_07479_),
    .B(_07472_),
    .Y(_07491_));
 sky130_fd_sc_hd__a21bo_1 _14341_ (.A1(_07473_),
    .A2(_07489_),
    .B1_N(_07491_),
    .X(_07492_));
 sky130_fd_sc_hd__or3_4 _14342_ (.A(_07474_),
    .B(_07471_),
    .C(net558),
    .X(_07493_));
 sky130_fd_sc_hd__nand2_1 _14343_ (.A(_07492_),
    .B(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__a21o_1 _14344_ (.A1(_07490_),
    .A2(_07494_),
    .B1(net7438),
    .X(_07495_));
 sky130_fd_sc_hd__and2b_1 _14345_ (.A_N(_07440_),
    .B(_07441_),
    .X(_07496_));
 sky130_fd_sc_hd__or2_1 _14346_ (.A(_07356_),
    .B(_07439_),
    .X(_07497_));
 sky130_fd_sc_hd__nand2_1 _14347_ (.A(_07082_),
    .B(_07467_),
    .Y(_07498_));
 sky130_fd_sc_hd__and2b_1 _14348_ (.A_N(_07497_),
    .B(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__or2b_1 _14349_ (.A(_07498_),
    .B_N(_07497_),
    .X(_07500_));
 sky130_fd_sc_hd__o31a_1 _14350_ (.A1(_07450_),
    .A2(_07496_),
    .A3(_07499_),
    .B1(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__and2_1 _14351_ (.A(_07495_),
    .B(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__nor2_1 _14352_ (.A(_07495_),
    .B(_07501_),
    .Y(_07503_));
 sky130_fd_sc_hd__or2_1 _14353_ (.A(_07502_),
    .B(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__and2_1 _14354_ (.A(_07478_),
    .B(_07484_),
    .X(_07505_));
 sky130_fd_sc_hd__or2_1 _14355_ (.A(_07485_),
    .B(_07505_),
    .X(_07506_));
 sky130_fd_sc_hd__a211o_1 _14356_ (.A1(net3246),
    .A2(_07468_),
    .B1(_07465_),
    .C1(_07311_),
    .X(_07507_));
 sky130_fd_sc_hd__or2b_1 _14357_ (.A(_07506_),
    .B_N(_07507_),
    .X(_07508_));
 sky130_fd_sc_hd__nand2_2 _14358_ (.A(net7757),
    .B(net558),
    .Y(_07509_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(_07473_),
    .B(_07475_),
    .Y(_07510_));
 sky130_fd_sc_hd__xnor2_1 _14360_ (.A(_07473_),
    .B(_07489_),
    .Y(_07511_));
 sky130_fd_sc_hd__a31o_1 _14361_ (.A1(_07491_),
    .A2(_07510_),
    .A3(_07511_),
    .B1(_07450_),
    .X(_07512_));
 sky130_fd_sc_hd__o211a_1 _14362_ (.A1(_07444_),
    .A2(_07509_),
    .B1(_07512_),
    .C1(net7757),
    .X(_07513_));
 sky130_fd_sc_hd__nand2_1 _14363_ (.A(_07361_),
    .B(_07403_),
    .Y(_07514_));
 sky130_fd_sc_hd__xnor2_1 _14364_ (.A(_07514_),
    .B(_07487_),
    .Y(_07515_));
 sky130_fd_sc_hd__xor2_1 _14365_ (.A(_07508_),
    .B(_07513_),
    .X(_07516_));
 sky130_fd_sc_hd__nand2_1 _14366_ (.A(_07515_),
    .B(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__o21a_1 _14367_ (.A1(_07508_),
    .A2(_07513_),
    .B1(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__xnor2_1 _14368_ (.A(_07504_),
    .B(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__xor2_1 _14369_ (.A(_07488_),
    .B(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__or2_1 _14370_ (.A(_06859_),
    .B(_07359_),
    .X(_07521_));
 sky130_fd_sc_hd__and2_1 _14371_ (.A(_07302_),
    .B(_07305_),
    .X(_07522_));
 sky130_fd_sc_hd__or2_2 _14372_ (.A(_07306_),
    .B(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__clkbuf_4 _14373_ (.A(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__nor3_1 _14374_ (.A(_07356_),
    .B(_07521_),
    .C(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__xnor2_1 _14375_ (.A(_07355_),
    .B(_07360_),
    .Y(_07526_));
 sky130_fd_sc_hd__or2_1 _14376_ (.A(_07361_),
    .B(_07403_),
    .X(_07527_));
 sky130_fd_sc_hd__nand2_1 _14377_ (.A(_07514_),
    .B(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__or2_1 _14378_ (.A(_07474_),
    .B(_07354_),
    .X(_07529_));
 sky130_fd_sc_hd__o22a_1 _14379_ (.A1(_07471_),
    .A2(_07400_),
    .B1(_07439_),
    .B2(_07367_),
    .X(_07530_));
 sky130_fd_sc_hd__nor2_1 _14380_ (.A(_07529_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__buf_2 _14381_ (.A(_06955_),
    .X(_07532_));
 sky130_fd_sc_hd__or3_2 _14382_ (.A(_06957_),
    .B(_07532_),
    .C(_07463_),
    .X(_07533_));
 sky130_fd_sc_hd__clkbuf_4 _14383_ (.A(_06957_),
    .X(_07534_));
 sky130_fd_sc_hd__a21oi_1 _14384_ (.A1(_07534_),
    .A2(_07532_),
    .B1(_07464_),
    .Y(_07535_));
 sky130_fd_sc_hd__and3_1 _14385_ (.A(_07533_),
    .B(_07535_),
    .C(_07465_),
    .X(_07536_));
 sky130_fd_sc_hd__a31o_1 _14386_ (.A1(net587),
    .A2(net3333),
    .A3(_07467_),
    .B1(_07536_),
    .X(_07537_));
 sky130_fd_sc_hd__nor2_1 _14387_ (.A(_07481_),
    .B(_07482_),
    .Y(_07538_));
 sky130_fd_sc_hd__or2_1 _14388_ (.A(_07483_),
    .B(_07538_),
    .X(_07539_));
 sky130_fd_sc_hd__xnor2_2 _14389_ (.A(_07537_),
    .B(_07539_),
    .Y(_07540_));
 sky130_fd_sc_hd__and2b_1 _14390_ (.A_N(_07539_),
    .B(_07537_),
    .X(_07541_));
 sky130_fd_sc_hd__a21oi_1 _14391_ (.A1(_07531_),
    .A2(_07540_),
    .B1(_07541_),
    .Y(_07542_));
 sky130_fd_sc_hd__nor2_1 _14392_ (.A(_07528_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__and2_1 _14393_ (.A(_07528_),
    .B(_07542_),
    .X(_07544_));
 sky130_fd_sc_hd__nor2_1 _14394_ (.A(_07543_),
    .B(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__a31o_1 _14395_ (.A1(_07525_),
    .A2(_07526_),
    .A3(_07545_),
    .B1(_07543_),
    .X(_07546_));
 sky130_fd_sc_hd__or2_1 _14396_ (.A(_07515_),
    .B(_07516_),
    .X(_07547_));
 sky130_fd_sc_hd__nand2_1 _14397_ (.A(_07517_),
    .B(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__nand2_1 _14398_ (.A(_07525_),
    .B(_07526_),
    .Y(_07549_));
 sky130_fd_sc_hd__xnor2_1 _14399_ (.A(_07549_),
    .B(_07545_),
    .Y(_07550_));
 sky130_fd_sc_hd__xor2_2 _14400_ (.A(_07465_),
    .B(_07469_),
    .X(_07551_));
 sky130_fd_sc_hd__xor2_2 _14401_ (.A(_07531_),
    .B(_07540_),
    .X(_07552_));
 sky130_fd_sc_hd__xnor2_1 _14402_ (.A(_07507_),
    .B(_07506_),
    .Y(_07553_));
 sky130_fd_sc_hd__and3_1 _14403_ (.A(_07551_),
    .B(_07552_),
    .C(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__a21oi_1 _14404_ (.A1(_07551_),
    .A2(_07552_),
    .B1(_07553_),
    .Y(_07555_));
 sky130_fd_sc_hd__nor2_1 _14405_ (.A(_07554_),
    .B(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__a21oi_1 _14406_ (.A1(_07550_),
    .A2(_07556_),
    .B1(_07554_),
    .Y(_07557_));
 sky130_fd_sc_hd__nor2_1 _14407_ (.A(_07548_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__and2_1 _14408_ (.A(_07548_),
    .B(_07557_),
    .X(_07559_));
 sky130_fd_sc_hd__nor2_1 _14409_ (.A(_07558_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__a21oi_1 _14410_ (.A1(_07546_),
    .A2(_07560_),
    .B1(_07558_),
    .Y(_07561_));
 sky130_fd_sc_hd__nor2_1 _14411_ (.A(_07520_),
    .B(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__o21bai_2 _14412_ (.A1(_07471_),
    .A2(_07509_),
    .B1_N(_07489_),
    .Y(_07563_));
 sky130_fd_sc_hd__and3_1 _14413_ (.A(_07467_),
    .B(_07500_),
    .C(_07494_),
    .X(_07564_));
 sky130_fd_sc_hd__a21o_1 _14414_ (.A1(_07493_),
    .A2(_07563_),
    .B1(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__nand3_4 _14415_ (.A(_07493_),
    .B(_07564_),
    .C(_07563_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_2 _14416_ (.A(_07502_),
    .B(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__a21boi_2 _14417_ (.A1(_07565_),
    .A2(_07567_),
    .B1_N(_07500_),
    .Y(_07568_));
 sky130_fd_sc_hd__or2b_1 _14418_ (.A(_07519_),
    .B_N(_07488_),
    .X(_07569_));
 sky130_fd_sc_hd__o21a_1 _14419_ (.A1(_07504_),
    .A2(_07518_),
    .B1(_07569_),
    .X(_07570_));
 sky130_fd_sc_hd__xor2_1 _14420_ (.A(_07568_),
    .B(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__and2_1 _14421_ (.A(_07562_),
    .B(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__nor2_1 _14422_ (.A(_07568_),
    .B(_07570_),
    .Y(_07573_));
 sky130_fd_sc_hd__and2_1 _14423_ (.A(_07467_),
    .B(_07493_),
    .X(_07574_));
 sky130_fd_sc_hd__nor2_1 _14424_ (.A(_07474_),
    .B(_07509_),
    .Y(_07575_));
 sky130_fd_sc_hd__o311a_2 _14425_ (.A1(net7438),
    .A2(_07574_),
    .A3(_07575_),
    .B1(_07494_),
    .C1(_07566_),
    .X(_07576_));
 sky130_fd_sc_hd__xnor2_2 _14426_ (.A(_07567_),
    .B(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__nand2_2 _14427_ (.A(_07573_),
    .B(_07577_),
    .Y(_07578_));
 sky130_fd_sc_hd__or2_1 _14428_ (.A(_07573_),
    .B(_07577_),
    .X(_07579_));
 sky130_fd_sc_hd__and2_1 _14429_ (.A(_07578_),
    .B(_07579_),
    .X(_07580_));
 sky130_fd_sc_hd__nand2_1 _14430_ (.A(_07572_),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__or2_1 _14431_ (.A(_07572_),
    .B(_07580_),
    .X(_07582_));
 sky130_fd_sc_hd__and2_1 _14432_ (.A(_07581_),
    .B(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__inv_2 _14433_ (.A(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__xnor2_2 _14434_ (.A(_07546_),
    .B(_07560_),
    .Y(_07585_));
 sky130_fd_sc_hd__xnor2_1 _14435_ (.A(_07550_),
    .B(_07556_),
    .Y(_07586_));
 sky130_fd_sc_hd__nor2_1 _14436_ (.A(_06859_),
    .B(_07524_),
    .Y(_07587_));
 sky130_fd_sc_hd__and2_1 _14437_ (.A(_07303_),
    .B(_07304_),
    .X(_07588_));
 sky130_fd_sc_hd__nor2_1 _14438_ (.A(_07305_),
    .B(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__clkbuf_4 _14439_ (.A(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__nor2_1 _14440_ (.A(_07356_),
    .B(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_1 _14441_ (.A(_07587_),
    .B(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__o21a_1 _14442_ (.A1(_07356_),
    .A2(_07524_),
    .B1(_07521_),
    .X(_07593_));
 sky130_fd_sc_hd__o21a_1 _14443_ (.A1(_07525_),
    .A2(_07593_),
    .B1(net7757),
    .X(_07594_));
 sky130_fd_sc_hd__nor2_1 _14444_ (.A(_07592_),
    .B(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__or2_1 _14445_ (.A(_07525_),
    .B(_07526_),
    .X(_07596_));
 sky130_fd_sc_hd__nand2_1 _14446_ (.A(_07549_),
    .B(_07596_),
    .Y(_07597_));
 sky130_fd_sc_hd__nand2_2 _14447_ (.A(_07533_),
    .B(_07535_),
    .Y(_07598_));
 sky130_fd_sc_hd__or3_1 _14448_ (.A(_07444_),
    .B(_07598_),
    .C(_07439_),
    .X(_07599_));
 sky130_fd_sc_hd__and2_1 _14449_ (.A(_07529_),
    .B(_07530_),
    .X(_07600_));
 sky130_fd_sc_hd__or2_1 _14450_ (.A(_07531_),
    .B(_07600_),
    .X(_07601_));
 sky130_fd_sc_hd__a21o_1 _14451_ (.A1(_07533_),
    .A2(_07599_),
    .B1(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__nand3_1 _14452_ (.A(_07533_),
    .B(_07599_),
    .C(_07601_),
    .Y(_07603_));
 sky130_fd_sc_hd__nand2_2 _14453_ (.A(_07602_),
    .B(_07603_),
    .Y(_07604_));
 sky130_fd_sc_hd__nor2_1 _14454_ (.A(_07474_),
    .B(_07358_),
    .Y(_07605_));
 sky130_fd_sc_hd__or2_1 _14455_ (.A(_07367_),
    .B(_07399_),
    .X(_07606_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_07366_),
    .B(_07353_),
    .Y(_07607_));
 sky130_fd_sc_hd__xnor2_2 _14457_ (.A(_07606_),
    .B(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__or3_1 _14458_ (.A(_07471_),
    .B(_07354_),
    .C(_07606_),
    .X(_07609_));
 sky130_fd_sc_hd__a21boi_4 _14459_ (.A1(_07605_),
    .A2(_07608_),
    .B1_N(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__o21a_1 _14460_ (.A1(_07604_),
    .A2(_07610_),
    .B1(_07602_),
    .X(_07611_));
 sky130_fd_sc_hd__nor2_1 _14461_ (.A(_07597_),
    .B(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__and2_1 _14462_ (.A(_07597_),
    .B(_07611_),
    .X(_07613_));
 sky130_fd_sc_hd__nor2_1 _14463_ (.A(_07612_),
    .B(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__xor2_1 _14464_ (.A(_07595_),
    .B(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__xnor2_1 _14465_ (.A(_07551_),
    .B(_07552_),
    .Y(_07616_));
 sky130_fd_sc_hd__xor2_4 _14466_ (.A(_07604_),
    .B(_07610_),
    .X(_07617_));
 sky130_fd_sc_hd__clkbuf_4 _14467_ (.A(_06922_),
    .X(_07618_));
 sky130_fd_sc_hd__a21oi_1 _14468_ (.A1(_07533_),
    .A2(_07535_),
    .B1(_07465_),
    .Y(_07619_));
 sky130_fd_sc_hd__o221a_2 _14469_ (.A1(_07618_),
    .A2(_07509_),
    .B1(_07619_),
    .B2(_07536_),
    .C1(_06611_),
    .X(_07620_));
 sky130_fd_sc_hd__nor2_2 _14470_ (.A(_07444_),
    .B(_07439_),
    .Y(_07621_));
 sky130_fd_sc_hd__xnor2_4 _14471_ (.A(_07598_),
    .B(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__and3b_2 _14472_ (.A_N(_06922_),
    .B(_07466_),
    .C(_06923_),
    .X(_07623_));
 sky130_fd_sc_hd__nor2_1 _14473_ (.A(_07618_),
    .B(_07464_),
    .Y(_07624_));
 sky130_fd_sc_hd__a21oi_1 _14474_ (.A1(_06923_),
    .A2(_07468_),
    .B1(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__nor2_2 _14475_ (.A(_07623_),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__a21oi_4 _14476_ (.A1(_07622_),
    .A2(_07626_),
    .B1(_07623_),
    .Y(_07627_));
 sky130_fd_sc_hd__xor2_4 _14477_ (.A(_07620_),
    .B(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__nor2_1 _14478_ (.A(_07620_),
    .B(_07627_),
    .Y(_07629_));
 sky130_fd_sc_hd__a21oi_1 _14479_ (.A1(_07617_),
    .A2(_07628_),
    .B1(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__xor2_1 _14480_ (.A(_07616_),
    .B(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__nor2_1 _14481_ (.A(_07616_),
    .B(_07630_),
    .Y(_07632_));
 sky130_fd_sc_hd__a21oi_1 _14482_ (.A1(_07615_),
    .A2(_07631_),
    .B1(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__xnor2_1 _14483_ (.A(_07586_),
    .B(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__a21o_1 _14484_ (.A1(_07595_),
    .A2(_07614_),
    .B1(_07612_),
    .X(_07635_));
 sky130_fd_sc_hd__or2b_1 _14485_ (.A(_07634_),
    .B_N(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__o21a_1 _14486_ (.A1(_07586_),
    .A2(_07633_),
    .B1(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__nor2_1 _14487_ (.A(_07585_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__and2_1 _14488_ (.A(_07520_),
    .B(_07561_),
    .X(_07639_));
 sky130_fd_sc_hd__nor2_1 _14489_ (.A(_07562_),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__xor2_1 _14490_ (.A(_07638_),
    .B(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__xor2_1 _14491_ (.A(_07635_),
    .B(_07634_),
    .X(_07642_));
 sky130_fd_sc_hd__xnor2_1 _14492_ (.A(_07615_),
    .B(_07631_),
    .Y(_07643_));
 sky130_fd_sc_hd__nor2_1 _14493_ (.A(_06859_),
    .B(_07590_),
    .Y(_07644_));
 sky130_fd_sc_hd__or2_1 _14494_ (.A(_07356_),
    .B(_07304_),
    .X(_07645_));
 sky130_fd_sc_hd__inv_2 _14495_ (.A(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__nand2_1 _14496_ (.A(_07644_),
    .B(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__xnor2_1 _14497_ (.A(_07587_),
    .B(_07591_),
    .Y(_07648_));
 sky130_fd_sc_hd__or2_2 _14498_ (.A(_07647_),
    .B(_07648_),
    .X(_07649_));
 sky130_fd_sc_hd__and2_1 _14499_ (.A(_07592_),
    .B(_07594_),
    .X(_07650_));
 sky130_fd_sc_hd__or2_2 _14500_ (.A(_07595_),
    .B(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__or4_4 _14501_ (.A(_06957_),
    .B(_07532_),
    .C(_07463_),
    .D(_07438_),
    .X(_07652_));
 sky130_fd_sc_hd__a2bb2o_1 _14502_ (.A1_N(_07438_),
    .A2_N(_07532_),
    .B1(net586),
    .B2(_07466_),
    .X(_07653_));
 sky130_fd_sc_hd__nor2_1 _14503_ (.A(_07444_),
    .B(_07400_),
    .Y(_07654_));
 sky130_fd_sc_hd__nand3_1 _14504_ (.A(_07652_),
    .B(_07653_),
    .C(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__xnor2_1 _14505_ (.A(_07605_),
    .B(_07608_),
    .Y(_07656_));
 sky130_fd_sc_hd__a21o_1 _14506_ (.A1(_07652_),
    .A2(_07655_),
    .B1(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__nand3_1 _14507_ (.A(_07652_),
    .B(_07655_),
    .C(_07656_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand2_2 _14508_ (.A(_07657_),
    .B(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__nor2_1 _14509_ (.A(_07474_),
    .B(_07523_),
    .Y(_07660_));
 sky130_fd_sc_hd__or2_1 _14510_ (.A(_07367_),
    .B(_07353_),
    .X(_07661_));
 sky130_fd_sc_hd__nor2_1 _14511_ (.A(_07366_),
    .B(_07358_),
    .Y(_07662_));
 sky130_fd_sc_hd__xnor2_2 _14512_ (.A(_07661_),
    .B(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__or3_1 _14513_ (.A(_07471_),
    .B(_07359_),
    .C(_07661_),
    .X(_07664_));
 sky130_fd_sc_hd__a21boi_4 _14514_ (.A1(_07660_),
    .A2(_07663_),
    .B1_N(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__o21a_2 _14515_ (.A1(_07659_),
    .A2(_07665_),
    .B1(_07657_),
    .X(_07666_));
 sky130_fd_sc_hd__xor2_4 _14516_ (.A(_07651_),
    .B(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__xnor2_4 _14517_ (.A(_07649_),
    .B(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__xnor2_4 _14518_ (.A(_07617_),
    .B(_07628_),
    .Y(_07669_));
 sky130_fd_sc_hd__xor2_4 _14519_ (.A(_07659_),
    .B(_07665_),
    .X(_07670_));
 sky130_fd_sc_hd__xnor2_4 _14520_ (.A(_07622_),
    .B(_07626_),
    .Y(_07671_));
 sky130_fd_sc_hd__a221oi_1 _14521_ (.A1(_06923_),
    .A2(_07467_),
    .B1(_07468_),
    .B2(_07090_),
    .C1(_07624_),
    .Y(_07672_));
 sky130_fd_sc_hd__a21o_1 _14522_ (.A1(_07652_),
    .A2(_07653_),
    .B1(_07654_),
    .X(_07673_));
 sky130_fd_sc_hd__nand2_1 _14523_ (.A(_07655_),
    .B(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__or3_2 _14524_ (.A(_07232_),
    .B(_06918_),
    .C(_07463_),
    .X(_07675_));
 sky130_fd_sc_hd__or3_4 _14525_ (.A(_07083_),
    .B(_06922_),
    .C(_07463_),
    .X(_07676_));
 sky130_fd_sc_hd__a21o_1 _14526_ (.A1(_07675_),
    .A2(_07676_),
    .B1(_07623_),
    .X(_07677_));
 sky130_fd_sc_hd__o21a_2 _14527_ (.A1(_07672_),
    .A2(_07674_),
    .B1(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__xor2_4 _14528_ (.A(_07671_),
    .B(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__nor2_1 _14529_ (.A(_07671_),
    .B(_07678_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21oi_4 _14530_ (.A1(_07670_),
    .A2(_07679_),
    .B1(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__xor2_4 _14531_ (.A(_07669_),
    .B(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__nor2_1 _14532_ (.A(_07669_),
    .B(_07681_),
    .Y(_07683_));
 sky130_fd_sc_hd__a21oi_1 _14533_ (.A1(_07668_),
    .A2(_07682_),
    .B1(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__xnor2_1 _14534_ (.A(_07643_),
    .B(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__or2b_1 _14535_ (.A(_07649_),
    .B_N(_07667_),
    .X(_07686_));
 sky130_fd_sc_hd__o21ai_2 _14536_ (.A1(_07651_),
    .A2(_07666_),
    .B1(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__or2b_1 _14537_ (.A(_07685_),
    .B_N(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__o21a_1 _14538_ (.A1(_07643_),
    .A2(_07684_),
    .B1(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__nor2_1 _14539_ (.A(_07642_),
    .B(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__xor2_2 _14540_ (.A(_07585_),
    .B(_07637_),
    .X(_07691_));
 sky130_fd_sc_hd__and2_1 _14541_ (.A(_07690_),
    .B(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__and2_1 _14542_ (.A(_07641_),
    .B(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__nor2_1 _14543_ (.A(_07641_),
    .B(_07692_),
    .Y(_07694_));
 sky130_fd_sc_hd__nor2_2 _14544_ (.A(_07693_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__xor2_2 _14545_ (.A(_07687_),
    .B(_07685_),
    .X(_07696_));
 sky130_fd_sc_hd__or4_4 _14546_ (.A(_06957_),
    .B(_06955_),
    .C(_07399_),
    .D(_07438_),
    .X(_07697_));
 sky130_fd_sc_hd__o22ai_2 _14547_ (.A1(_07532_),
    .A2(_07400_),
    .B1(_07439_),
    .B2(_07534_),
    .Y(_07698_));
 sky130_fd_sc_hd__nor2_1 _14548_ (.A(_06990_),
    .B(_07354_),
    .Y(_07699_));
 sky130_fd_sc_hd__nand3_1 _14549_ (.A(_07697_),
    .B(_07698_),
    .C(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__xnor2_1 _14550_ (.A(_07660_),
    .B(_07663_),
    .Y(_07701_));
 sky130_fd_sc_hd__a21o_1 _14551_ (.A1(_07697_),
    .A2(_07700_),
    .B1(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__nand3_1 _14552_ (.A(_07697_),
    .B(_07700_),
    .C(_07701_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_1 _14553_ (.A(_07702_),
    .B(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__nor2_1 _14554_ (.A(_07474_),
    .B(_07589_),
    .Y(_07705_));
 sky130_fd_sc_hd__or2_1 _14555_ (.A(_07367_),
    .B(_07358_),
    .X(_07706_));
 sky130_fd_sc_hd__nor2_1 _14556_ (.A(_07366_),
    .B(_07523_),
    .Y(_07707_));
 sky130_fd_sc_hd__xnor2_1 _14557_ (.A(_07706_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__or3_1 _14558_ (.A(_07471_),
    .B(_07524_),
    .C(_07706_),
    .X(_07709_));
 sky130_fd_sc_hd__a21boi_2 _14559_ (.A1(_07705_),
    .A2(_07708_),
    .B1_N(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__or2_1 _14560_ (.A(_07704_),
    .B(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__nand2_1 _14561_ (.A(_07647_),
    .B(_07648_),
    .Y(_07712_));
 sky130_fd_sc_hd__nand2_1 _14562_ (.A(_07649_),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__a21oi_4 _14563_ (.A1(_07702_),
    .A2(_07711_),
    .B1(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__xnor2_4 _14564_ (.A(_07668_),
    .B(_07682_),
    .Y(_07715_));
 sky130_fd_sc_hd__and3_1 _14565_ (.A(_07702_),
    .B(_07711_),
    .C(_07713_),
    .X(_07716_));
 sky130_fd_sc_hd__nor2_1 _14566_ (.A(_07714_),
    .B(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__xor2_2 _14567_ (.A(_07670_),
    .B(_07679_),
    .X(_07718_));
 sky130_fd_sc_hd__xor2_2 _14568_ (.A(_07704_),
    .B(_07710_),
    .X(_07719_));
 sky130_fd_sc_hd__or2b_1 _14569_ (.A(_07672_),
    .B_N(_07677_),
    .X(_07720_));
 sky130_fd_sc_hd__xnor2_2 _14570_ (.A(_07674_),
    .B(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__a21oi_2 _14571_ (.A1(_07083_),
    .A2(_07618_),
    .B1(_07464_),
    .Y(_07722_));
 sky130_fd_sc_hd__nand2_2 _14572_ (.A(_06865_),
    .B(_07467_),
    .Y(_07723_));
 sky130_fd_sc_hd__or2_2 _14573_ (.A(_07618_),
    .B(_07438_),
    .X(_07724_));
 sky130_fd_sc_hd__o21ai_4 _14574_ (.A1(_07723_),
    .A2(_07724_),
    .B1(_07675_),
    .Y(_07725_));
 sky130_fd_sc_hd__a21o_1 _14575_ (.A1(_07697_),
    .A2(_07698_),
    .B1(_07699_),
    .X(_07726_));
 sky130_fd_sc_hd__and2_2 _14576_ (.A(_07700_),
    .B(_07726_),
    .X(_07727_));
 sky130_fd_sc_hd__nand2_1 _14577_ (.A(_07676_),
    .B(_07722_),
    .Y(_07728_));
 sky130_fd_sc_hd__xnor2_2 _14578_ (.A(_07728_),
    .B(_07725_),
    .Y(_07729_));
 sky130_fd_sc_hd__a32oi_4 _14579_ (.A1(_07676_),
    .A2(_07722_),
    .A3(_07725_),
    .B1(_07727_),
    .B2(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__xor2_2 _14580_ (.A(_07721_),
    .B(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__nor2_1 _14581_ (.A(_07721_),
    .B(_07730_),
    .Y(_07732_));
 sky130_fd_sc_hd__a21oi_2 _14582_ (.A1(_07719_),
    .A2(_07731_),
    .B1(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__xnor2_2 _14583_ (.A(_07718_),
    .B(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__and2b_1 _14584_ (.A_N(_07733_),
    .B(_07718_),
    .X(_07735_));
 sky130_fd_sc_hd__a21oi_2 _14585_ (.A1(_07717_),
    .A2(_07734_),
    .B1(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__xor2_4 _14586_ (.A(_07715_),
    .B(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__nor2_1 _14587_ (.A(_07715_),
    .B(_07736_),
    .Y(_07738_));
 sky130_fd_sc_hd__a21oi_2 _14588_ (.A1(_07714_),
    .A2(_07737_),
    .B1(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__nor2_1 _14589_ (.A(_07696_),
    .B(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_1 _14590_ (.A(_07642_),
    .B(_07689_),
    .Y(_07741_));
 sky130_fd_sc_hd__and2b_1 _14591_ (.A_N(_07690_),
    .B(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__xnor2_4 _14592_ (.A(_07714_),
    .B(_07737_),
    .Y(_07743_));
 sky130_fd_sc_hd__or2_1 _14593_ (.A(_06955_),
    .B(_07353_),
    .X(_07744_));
 sky130_fd_sc_hd__or3_1 _14594_ (.A(_07534_),
    .B(_07400_),
    .C(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__nor2_1 _14595_ (.A(_07534_),
    .B(_07399_),
    .Y(_07746_));
 sky130_fd_sc_hd__xnor2_1 _14596_ (.A(_07746_),
    .B(_07744_),
    .Y(_07747_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(_06990_),
    .B(_07359_),
    .Y(_07748_));
 sky130_fd_sc_hd__nand2_1 _14598_ (.A(_07747_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__xnor2_1 _14599_ (.A(_07705_),
    .B(_07708_),
    .Y(_07750_));
 sky130_fd_sc_hd__a21o_1 _14600_ (.A1(_07745_),
    .A2(_07749_),
    .B1(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__nand3_1 _14601_ (.A(_07745_),
    .B(_07749_),
    .C(_07750_),
    .Y(_07752_));
 sky130_fd_sc_hd__nand2_1 _14602_ (.A(_07751_),
    .B(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__or2_1 _14603_ (.A(_07367_),
    .B(_07523_),
    .X(_07754_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(_07474_),
    .B(_07304_),
    .Y(_07755_));
 sky130_fd_sc_hd__nor2_1 _14605_ (.A(_07366_),
    .B(_07589_),
    .Y(_07756_));
 sky130_fd_sc_hd__xnor2_1 _14606_ (.A(_07754_),
    .B(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__nand2_1 _14607_ (.A(_07755_),
    .B(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__o31a_1 _14608_ (.A1(_07471_),
    .A2(_07590_),
    .A3(_07754_),
    .B1(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__or2_1 _14609_ (.A(_07753_),
    .B(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__or2_1 _14610_ (.A(_07644_),
    .B(_07646_),
    .X(_07761_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_07647_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__a21oi_2 _14612_ (.A1(_07751_),
    .A2(_07760_),
    .B1(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__xnor2_2 _14613_ (.A(_07717_),
    .B(_07734_),
    .Y(_07764_));
 sky130_fd_sc_hd__and3_1 _14614_ (.A(_07751_),
    .B(_07760_),
    .C(_07762_),
    .X(_07765_));
 sky130_fd_sc_hd__nor2_1 _14615_ (.A(_07763_),
    .B(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__xnor2_2 _14616_ (.A(_07719_),
    .B(_07731_),
    .Y(_07767_));
 sky130_fd_sc_hd__xor2_2 _14617_ (.A(_07753_),
    .B(_07759_),
    .X(_07768_));
 sky130_fd_sc_hd__xnor2_4 _14618_ (.A(_07727_),
    .B(_07729_),
    .Y(_07769_));
 sky130_fd_sc_hd__or2_1 _14619_ (.A(_07747_),
    .B(_07748_),
    .X(_07770_));
 sky130_fd_sc_hd__and2_1 _14620_ (.A(_07749_),
    .B(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__xnor2_2 _14621_ (.A(_07723_),
    .B(_07724_),
    .Y(_07772_));
 sky130_fd_sc_hd__nor2_1 _14622_ (.A(_07618_),
    .B(_07400_),
    .Y(_07773_));
 sky130_fd_sc_hd__buf_2 _14623_ (.A(_06918_),
    .X(_07774_));
 sky130_fd_sc_hd__a2bb2o_1 _14624_ (.A1_N(_07439_),
    .A2_N(_07774_),
    .B1(_07090_),
    .B2(_07466_),
    .X(_07775_));
 sky130_fd_sc_hd__or4_4 _14625_ (.A(_07232_),
    .B(_06918_),
    .C(_07464_),
    .D(_07438_),
    .X(_07776_));
 sky130_fd_sc_hd__a21bo_4 _14626_ (.A1(_07773_),
    .A2(_07775_),
    .B1_N(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__xnor2_4 _14627_ (.A(_07772_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__and2b_1 _14628_ (.A_N(_07772_),
    .B(_07777_),
    .X(_07779_));
 sky130_fd_sc_hd__a21o_1 _14629_ (.A1(_07771_),
    .A2(_07778_),
    .B1(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__xnor2_2 _14630_ (.A(_07769_),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__or2b_1 _14631_ (.A(_07780_),
    .B_N(_07769_),
    .X(_07782_));
 sky130_fd_sc_hd__a21boi_4 _14632_ (.A1(_07768_),
    .A2(_07781_),
    .B1_N(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__xor2_2 _14633_ (.A(_07767_),
    .B(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__nor2_1 _14634_ (.A(_07767_),
    .B(_07783_),
    .Y(_07785_));
 sky130_fd_sc_hd__a21oi_2 _14635_ (.A1(_07766_),
    .A2(_07784_),
    .B1(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__xor2_2 _14636_ (.A(_07764_),
    .B(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__nor2_1 _14637_ (.A(_07764_),
    .B(_07786_),
    .Y(_07788_));
 sky130_fd_sc_hd__a21oi_2 _14638_ (.A1(_07763_),
    .A2(_07787_),
    .B1(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__nor2_1 _14639_ (.A(_07743_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__xor2_2 _14640_ (.A(_07696_),
    .B(_07739_),
    .X(_07791_));
 sky130_fd_sc_hd__and2_1 _14641_ (.A(_07790_),
    .B(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__nor2_1 _14642_ (.A(_07740_),
    .B(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__xnor2_1 _14643_ (.A(_07742_),
    .B(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__xor2_4 _14644_ (.A(_07743_),
    .B(_07789_),
    .X(_07795_));
 sky130_fd_sc_hd__xnor2_2 _14645_ (.A(_07763_),
    .B(_07787_),
    .Y(_07796_));
 sky130_fd_sc_hd__nor2_1 _14646_ (.A(_07534_),
    .B(_07353_),
    .Y(_07797_));
 sky130_fd_sc_hd__nor2_1 _14647_ (.A(_07532_),
    .B(_07358_),
    .Y(_07798_));
 sky130_fd_sc_hd__nand2_1 _14648_ (.A(_07797_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__xnor2_1 _14649_ (.A(_07797_),
    .B(_07798_),
    .Y(_07800_));
 sky130_fd_sc_hd__or3_1 _14650_ (.A(_07444_),
    .B(_07523_),
    .C(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__xnor2_1 _14651_ (.A(_07755_),
    .B(_07757_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand3_1 _14652_ (.A(_07799_),
    .B(_07801_),
    .C(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__or2_1 _14653_ (.A(_07367_),
    .B(_07590_),
    .X(_07804_));
 sky130_fd_sc_hd__clkbuf_4 _14654_ (.A(_07304_),
    .X(_07805_));
 sky130_fd_sc_hd__nor2_1 _14655_ (.A(_07471_),
    .B(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__and2b_1 _14656_ (.A_N(_07804_),
    .B(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__a21o_1 _14657_ (.A1(_07799_),
    .A2(_07801_),
    .B1(_07802_),
    .X(_07808_));
 sky130_fd_sc_hd__a21boi_1 _14658_ (.A1(_07803_),
    .A2(_07807_),
    .B1_N(_07808_),
    .Y(_07809_));
 sky130_fd_sc_hd__nor2_1 _14659_ (.A(_06859_),
    .B(_07805_),
    .Y(_07810_));
 sky130_fd_sc_hd__nor2b_1 _14660_ (.A(_07809_),
    .B_N(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__xnor2_2 _14661_ (.A(_07766_),
    .B(_07784_),
    .Y(_07812_));
 sky130_fd_sc_hd__and2b_1 _14662_ (.A_N(_07810_),
    .B(_07809_),
    .X(_07813_));
 sky130_fd_sc_hd__nor2_1 _14663_ (.A(_07811_),
    .B(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__xnor2_2 _14664_ (.A(_07768_),
    .B(_07781_),
    .Y(_07815_));
 sky130_fd_sc_hd__nand2_1 _14665_ (.A(_07808_),
    .B(_07803_),
    .Y(_07816_));
 sky130_fd_sc_hd__xnor2_1 _14666_ (.A(_07816_),
    .B(_07807_),
    .Y(_07817_));
 sky130_fd_sc_hd__xnor2_2 _14667_ (.A(_07771_),
    .B(_07778_),
    .Y(_07818_));
 sky130_fd_sc_hd__o21ai_1 _14668_ (.A1(_07444_),
    .A2(_07524_),
    .B1(_07800_),
    .Y(_07819_));
 sky130_fd_sc_hd__and2_1 _14669_ (.A(_07801_),
    .B(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__nand3_1 _14670_ (.A(_07776_),
    .B(_07773_),
    .C(_07775_),
    .Y(_07821_));
 sky130_fd_sc_hd__a21o_1 _14671_ (.A1(_07776_),
    .A2(_07775_),
    .B1(_07773_),
    .X(_07822_));
 sky130_fd_sc_hd__nor2_1 _14672_ (.A(_07618_),
    .B(_07354_),
    .Y(_07823_));
 sky130_fd_sc_hd__o22ai_2 _14673_ (.A1(_07774_),
    .A2(_07400_),
    .B1(_07439_),
    .B2(_07232_),
    .Y(_07824_));
 sky130_fd_sc_hd__or4_4 _14674_ (.A(_07232_),
    .B(_07774_),
    .C(_07400_),
    .D(_07438_),
    .X(_07825_));
 sky130_fd_sc_hd__a21bo_1 _14675_ (.A1(_07823_),
    .A2(_07824_),
    .B1_N(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__a21o_1 _14676_ (.A1(_07821_),
    .A2(_07822_),
    .B1(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__nand3_1 _14677_ (.A(_07821_),
    .B(_07822_),
    .C(_07826_),
    .Y(_07828_));
 sky130_fd_sc_hd__a21boi_2 _14678_ (.A1(_07820_),
    .A2(_07827_),
    .B1_N(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__xor2_2 _14679_ (.A(_07818_),
    .B(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__nor2_1 _14680_ (.A(_07818_),
    .B(_07829_),
    .Y(_07831_));
 sky130_fd_sc_hd__a21oi_2 _14681_ (.A1(_07817_),
    .A2(_07830_),
    .B1(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__xor2_2 _14682_ (.A(_07815_),
    .B(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__nor2_1 _14683_ (.A(_07815_),
    .B(_07832_),
    .Y(_07834_));
 sky130_fd_sc_hd__a21oi_2 _14684_ (.A1(_07814_),
    .A2(_07833_),
    .B1(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__xor2_2 _14685_ (.A(_07812_),
    .B(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__nor2_1 _14686_ (.A(_07812_),
    .B(_07835_),
    .Y(_07837_));
 sky130_fd_sc_hd__a21oi_2 _14687_ (.A1(_07811_),
    .A2(_07836_),
    .B1(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__nor2_1 _14688_ (.A(_07796_),
    .B(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__and2_1 _14689_ (.A(_07795_),
    .B(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__nor2_1 _14690_ (.A(_07790_),
    .B(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__xnor2_2 _14691_ (.A(_07791_),
    .B(_07841_),
    .Y(_07842_));
 sky130_fd_sc_hd__xor2_2 _14692_ (.A(_07796_),
    .B(_07838_),
    .X(_07843_));
 sky130_fd_sc_hd__or2_1 _14693_ (.A(_07532_),
    .B(_07523_),
    .X(_07844_));
 sky130_fd_sc_hd__or3_1 _14694_ (.A(_07534_),
    .B(_07359_),
    .C(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__nor2_1 _14695_ (.A(_07534_),
    .B(_07359_),
    .Y(_07846_));
 sky130_fd_sc_hd__xnor2_1 _14696_ (.A(_07846_),
    .B(_07844_),
    .Y(_07847_));
 sky130_fd_sc_hd__nor2_1 _14697_ (.A(_07444_),
    .B(_07590_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand2_1 _14698_ (.A(_07847_),
    .B(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__xor2_1 _14699_ (.A(_07804_),
    .B(_07806_),
    .X(_07850_));
 sky130_fd_sc_hd__a21oi_2 _14700_ (.A1(_07845_),
    .A2(_07849_),
    .B1(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__xnor2_1 _14701_ (.A(_07817_),
    .B(_07830_),
    .Y(_07852_));
 sky130_fd_sc_hd__and3_1 _14702_ (.A(_07845_),
    .B(_07849_),
    .C(_07850_),
    .X(_07853_));
 sky130_fd_sc_hd__nor2_1 _14703_ (.A(_07851_),
    .B(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand3_1 _14704_ (.A(_07828_),
    .B(_07820_),
    .C(_07827_),
    .Y(_07855_));
 sky130_fd_sc_hd__a21o_1 _14705_ (.A1(_07828_),
    .A2(_07827_),
    .B1(_07820_),
    .X(_07856_));
 sky130_fd_sc_hd__or2_1 _14706_ (.A(_07847_),
    .B(_07848_),
    .X(_07857_));
 sky130_fd_sc_hd__and2_1 _14707_ (.A(_07849_),
    .B(_07857_),
    .X(_07858_));
 sky130_fd_sc_hd__nand3_1 _14708_ (.A(_07825_),
    .B(_07823_),
    .C(_07824_),
    .Y(_07859_));
 sky130_fd_sc_hd__a21o_1 _14709_ (.A1(_07825_),
    .A2(_07824_),
    .B1(_07823_),
    .X(_07860_));
 sky130_fd_sc_hd__nor2_1 _14710_ (.A(_07618_),
    .B(_07359_),
    .Y(_07861_));
 sky130_fd_sc_hd__or2_1 _14711_ (.A(_07232_),
    .B(_07399_),
    .X(_07862_));
 sky130_fd_sc_hd__nor2_1 _14712_ (.A(_06918_),
    .B(_07354_),
    .Y(_07863_));
 sky130_fd_sc_hd__xnor2_1 _14713_ (.A(_07862_),
    .B(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__or3_1 _14714_ (.A(_07774_),
    .B(_07354_),
    .C(_07862_),
    .X(_07865_));
 sky130_fd_sc_hd__a21bo_1 _14715_ (.A1(_07861_),
    .A2(_07864_),
    .B1_N(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__a21o_1 _14716_ (.A1(_07859_),
    .A2(_07860_),
    .B1(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__and3_1 _14717_ (.A(_07859_),
    .B(_07860_),
    .C(_07866_),
    .X(_07868_));
 sky130_fd_sc_hd__a21o_1 _14718_ (.A1(_07858_),
    .A2(_07867_),
    .B1(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__a21o_1 _14719_ (.A1(_07855_),
    .A2(_07856_),
    .B1(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__and3_1 _14720_ (.A(_07855_),
    .B(_07856_),
    .C(_07869_),
    .X(_07871_));
 sky130_fd_sc_hd__a21oi_1 _14721_ (.A1(_07854_),
    .A2(_07870_),
    .B1(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_1 _14722_ (.A(_07852_),
    .B(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__nor2_1 _14723_ (.A(_07852_),
    .B(_07872_),
    .Y(_07874_));
 sky130_fd_sc_hd__a21oi_1 _14724_ (.A1(_07851_),
    .A2(_07873_),
    .B1(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__xnor2_1 _14725_ (.A(_07814_),
    .B(_07833_),
    .Y(_07876_));
 sky130_fd_sc_hd__xor2_1 _14726_ (.A(_07811_),
    .B(_07836_),
    .X(_07877_));
 sky130_fd_sc_hd__nor3b_2 _14727_ (.A(_07875_),
    .B(_07876_),
    .C_N(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__and2_1 _14728_ (.A(_07843_),
    .B(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__xor2_1 _14729_ (.A(_07876_),
    .B(_07875_),
    .X(_07880_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_07877_),
    .B(_07880_),
    .Y(_07881_));
 sky130_fd_sc_hd__xor2_2 _14731_ (.A(_07843_),
    .B(net78),
    .X(_07882_));
 sky130_fd_sc_hd__and2b_1 _14732_ (.A_N(_07874_),
    .B(_07873_),
    .X(_07883_));
 sky130_fd_sc_hd__xor2_1 _14733_ (.A(_07851_),
    .B(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__and2b_1 _14734_ (.A_N(_07868_),
    .B(_07867_),
    .X(_07885_));
 sky130_fd_sc_hd__xnor2_1 _14735_ (.A(_07858_),
    .B(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__nor2_1 _14736_ (.A(_07534_),
    .B(_07524_),
    .Y(_07887_));
 sky130_fd_sc_hd__nor2_1 _14737_ (.A(_07532_),
    .B(_07590_),
    .Y(_07888_));
 sky130_fd_sc_hd__xnor2_1 _14738_ (.A(_07887_),
    .B(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__nor2_1 _14739_ (.A(_07444_),
    .B(_07805_),
    .Y(_07890_));
 sky130_fd_sc_hd__xnor2_1 _14740_ (.A(_07889_),
    .B(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__xnor2_1 _14741_ (.A(_07861_),
    .B(_07864_),
    .Y(_07892_));
 sky130_fd_sc_hd__or2_1 _14742_ (.A(_07232_),
    .B(_07354_),
    .X(_07893_));
 sky130_fd_sc_hd__nor2_1 _14743_ (.A(_07618_),
    .B(_07524_),
    .Y(_07894_));
 sky130_fd_sc_hd__nor2_1 _14744_ (.A(_07774_),
    .B(_07359_),
    .Y(_07895_));
 sky130_fd_sc_hd__xnor2_1 _14745_ (.A(_07893_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand2_1 _14746_ (.A(_07894_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__o31a_1 _14747_ (.A1(_07774_),
    .A2(_07359_),
    .A3(_07893_),
    .B1(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__nand2_1 _14748_ (.A(_07892_),
    .B(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__nor2_1 _14749_ (.A(_07892_),
    .B(_07898_),
    .Y(_07900_));
 sky130_fd_sc_hd__a21oi_1 _14750_ (.A1(_07891_),
    .A2(_07899_),
    .B1(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__or2_1 _14751_ (.A(_07886_),
    .B(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(_07887_),
    .B(_07888_),
    .Y(_07903_));
 sky130_fd_sc_hd__o31a_1 _14753_ (.A1(_07444_),
    .A2(_07805_),
    .A3(_07889_),
    .B1(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__or3_1 _14754_ (.A(_07367_),
    .B(_07805_),
    .C(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__o21ai_1 _14755_ (.A1(_07367_),
    .A2(_07805_),
    .B1(_07904_),
    .Y(_07906_));
 sky130_fd_sc_hd__and2_1 _14756_ (.A(_07905_),
    .B(_07906_),
    .X(_07907_));
 sky130_fd_sc_hd__nand2_1 _14757_ (.A(_07886_),
    .B(_07901_),
    .Y(_07908_));
 sky130_fd_sc_hd__and2_1 _14758_ (.A(_07902_),
    .B(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__nand2_1 _14759_ (.A(_07907_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__and2b_1 _14760_ (.A_N(_07871_),
    .B(_07870_),
    .X(_07911_));
 sky130_fd_sc_hd__xnor2_1 _14761_ (.A(_07854_),
    .B(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__a21oi_1 _14762_ (.A1(_07902_),
    .A2(_07910_),
    .B1(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__and3_1 _14763_ (.A(_07912_),
    .B(_07902_),
    .C(_07910_),
    .X(_07914_));
 sky130_fd_sc_hd__or3_1 _14764_ (.A(_07905_),
    .B(_07913_),
    .C(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__or2b_1 _14765_ (.A(_07913_),
    .B_N(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__and4_1 _14766_ (.A(_07877_),
    .B(_07884_),
    .C(_07916_),
    .D(_07880_),
    .X(_07917_));
 sky130_fd_sc_hd__xnor2_2 _14767_ (.A(_07882_),
    .B(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__or2_1 _14768_ (.A(_07534_),
    .B(_07590_),
    .X(_07919_));
 sky130_fd_sc_hd__or3_1 _14769_ (.A(_07532_),
    .B(_07805_),
    .C(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__o21ai_1 _14770_ (.A1(_07532_),
    .A2(_07805_),
    .B1(_07919_),
    .Y(_07921_));
 sky130_fd_sc_hd__nand2_1 _14771_ (.A(_07920_),
    .B(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__xnor2_1 _14772_ (.A(_07894_),
    .B(_07896_),
    .Y(_07923_));
 sky130_fd_sc_hd__nor2_1 _14773_ (.A(_07618_),
    .B(_07590_),
    .Y(_07924_));
 sky130_fd_sc_hd__or2_1 _14774_ (.A(_07232_),
    .B(_07359_),
    .X(_07925_));
 sky130_fd_sc_hd__nor2_1 _14775_ (.A(_07774_),
    .B(_07524_),
    .Y(_07926_));
 sky130_fd_sc_hd__xnor2_1 _14776_ (.A(_07925_),
    .B(_07926_),
    .Y(_07927_));
 sky130_fd_sc_hd__or3_1 _14777_ (.A(_07774_),
    .B(_07524_),
    .C(_07925_),
    .X(_07928_));
 sky130_fd_sc_hd__a21boi_1 _14778_ (.A1(_07924_),
    .A2(_07927_),
    .B1_N(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__or2_1 _14779_ (.A(_07923_),
    .B(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__nand2_1 _14780_ (.A(_07923_),
    .B(_07929_),
    .Y(_07931_));
 sky130_fd_sc_hd__nand2_1 _14781_ (.A(_07930_),
    .B(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__or2_1 _14782_ (.A(_07922_),
    .B(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__nand2_1 _14783_ (.A(_07922_),
    .B(_07932_),
    .Y(_07934_));
 sky130_fd_sc_hd__and2_1 _14784_ (.A(_07933_),
    .B(_07934_),
    .X(_07935_));
 sky130_fd_sc_hd__xnor2_1 _14785_ (.A(_07924_),
    .B(_07927_),
    .Y(_07936_));
 sky130_fd_sc_hd__or2_1 _14786_ (.A(_07232_),
    .B(_07524_),
    .X(_07937_));
 sky130_fd_sc_hd__nor2_1 _14787_ (.A(_07618_),
    .B(_07805_),
    .Y(_07938_));
 sky130_fd_sc_hd__nor2_1 _14788_ (.A(_07774_),
    .B(_07590_),
    .Y(_07939_));
 sky130_fd_sc_hd__xnor2_1 _14789_ (.A(_07937_),
    .B(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand2_1 _14790_ (.A(_07938_),
    .B(_07940_),
    .Y(_07941_));
 sky130_fd_sc_hd__o31a_1 _14791_ (.A1(_07774_),
    .A2(_07590_),
    .A3(_07937_),
    .B1(_07941_),
    .X(_07942_));
 sky130_fd_sc_hd__nor2_1 _14792_ (.A(_07534_),
    .B(_07805_),
    .Y(_07943_));
 sky130_fd_sc_hd__xor2_1 _14793_ (.A(_07936_),
    .B(_07942_),
    .X(_07944_));
 sky130_fd_sc_hd__nand2_1 _14794_ (.A(_07943_),
    .B(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__o21ai_1 _14795_ (.A1(_07936_),
    .A2(_07942_),
    .B1(_07945_),
    .Y(_07946_));
 sky130_fd_sc_hd__and3_1 _14796_ (.A(_07205_),
    .B(_07305_),
    .C(_07941_),
    .X(_07947_));
 sky130_fd_sc_hd__o211a_1 _14797_ (.A1(_07938_),
    .A2(_07940_),
    .B1(_07945_),
    .C1(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__o221a_1 _14798_ (.A1(_07943_),
    .A2(_07944_),
    .B1(_07946_),
    .B2(_07935_),
    .C1(_07948_),
    .X(_07949_));
 sky130_fd_sc_hd__a21oi_1 _14799_ (.A1(_07935_),
    .A2(_07946_),
    .B1(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__and2b_1 _14800_ (.A_N(_07900_),
    .B(_07899_),
    .X(_07951_));
 sky130_fd_sc_hd__xnor2_1 _14801_ (.A(_07891_),
    .B(_07951_),
    .Y(_07952_));
 sky130_fd_sc_hd__and3_1 _14802_ (.A(_07952_),
    .B(_07930_),
    .C(_07933_),
    .X(_07953_));
 sky130_fd_sc_hd__a21oi_1 _14803_ (.A1(_07920_),
    .A2(_07950_),
    .B1(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__a21oi_1 _14804_ (.A1(_07930_),
    .A2(_07933_),
    .B1(_07952_),
    .Y(_07955_));
 sky130_fd_sc_hd__o21bai_1 _14805_ (.A1(_07920_),
    .A2(_07950_),
    .B1_N(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__or2_1 _14806_ (.A(_07907_),
    .B(_07909_),
    .X(_07957_));
 sky130_fd_sc_hd__and2_1 _14807_ (.A(_07910_),
    .B(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__o21ai_1 _14808_ (.A1(_07913_),
    .A2(_07914_),
    .B1(_07905_),
    .Y(_07959_));
 sky130_fd_sc_hd__o2111a_1 _14809_ (.A1(_07954_),
    .A2(_07956_),
    .B1(_07958_),
    .C1(_07959_),
    .D1(_07915_),
    .X(_07960_));
 sky130_fd_sc_hd__o21ai_1 _14810_ (.A1(_07884_),
    .A2(_07916_),
    .B1(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2_1 _14811_ (.A(_07882_),
    .B(_07917_),
    .Y(_07962_));
 sky130_fd_sc_hd__o31ai_2 _14812_ (.A1(_07881_),
    .A2(_07918_),
    .A3(_07961_),
    .B1(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__nor2_2 _14813_ (.A(_07839_),
    .B(_07879_),
    .Y(_07964_));
 sky130_fd_sc_hd__xnor2_4 _14814_ (.A(_07795_),
    .B(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__a22o_1 _14815_ (.A1(_07795_),
    .A2(_07879_),
    .B1(_07963_),
    .B2(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__a22o_1 _14816_ (.A1(_07791_),
    .A2(_07840_),
    .B1(_07842_),
    .B2(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__a22o_1 _14817_ (.A1(_07742_),
    .A2(_07792_),
    .B1(_07794_),
    .B2(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__a21oi_1 _14818_ (.A1(_07740_),
    .A2(_07741_),
    .B1(_07690_),
    .Y(_07969_));
 sky130_fd_sc_hd__xnor2_1 _14819_ (.A(_07691_),
    .B(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__a32o_2 _14820_ (.A1(_07691_),
    .A2(_07740_),
    .A3(_07742_),
    .B1(_07968_),
    .B2(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__and2_1 _14821_ (.A(_07638_),
    .B(_07640_),
    .X(_07972_));
 sky130_fd_sc_hd__nor2_1 _14822_ (.A(_07562_),
    .B(_07571_),
    .Y(_07973_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(_07572_),
    .B(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__xnor2_1 _14824_ (.A(_07972_),
    .B(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__inv_2 _14825_ (.A(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__o21a_1 _14826_ (.A1(_07972_),
    .A2(_07693_),
    .B1(_07974_),
    .X(_07977_));
 sky130_fd_sc_hd__a31oi_4 _14827_ (.A1(_07695_),
    .A2(_07971_),
    .A3(_07976_),
    .B1(_07977_),
    .Y(_07978_));
 sky130_fd_sc_hd__nand2_2 _14828_ (.A(_07494_),
    .B(_07566_),
    .Y(_07979_));
 sky130_fd_sc_hd__o21a_1 _14829_ (.A1(_07467_),
    .A2(_07575_),
    .B1(_07498_),
    .X(_07980_));
 sky130_fd_sc_hd__o21a_2 _14830_ (.A1(net7438),
    .A2(_07980_),
    .B1(_07493_),
    .X(_07981_));
 sky130_fd_sc_hd__a32oi_4 _14831_ (.A1(_07502_),
    .A2(_07566_),
    .A3(_07576_),
    .B1(_07981_),
    .B2(_07979_),
    .Y(_07982_));
 sky130_fd_sc_hd__o21ai_4 _14832_ (.A1(_07979_),
    .A2(_07981_),
    .B1(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__xnor2_4 _14833_ (.A(_07578_),
    .B(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__a21o_1 _14834_ (.A1(_07578_),
    .A2(_07581_),
    .B1(_07983_),
    .X(_07985_));
 sky130_fd_sc_hd__o31ai_4 _14835_ (.A1(_07584_),
    .A2(_07978_),
    .A3(_07984_),
    .B1(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__o211a_1 _14836_ (.A1(_07356_),
    .A2(_07509_),
    .B1(_07498_),
    .C1(net7757),
    .X(_07987_));
 sky130_fd_sc_hd__nand3_2 _14837_ (.A(_07493_),
    .B(_07982_),
    .C(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__xor2_2 _14838_ (.A(_07986_),
    .B(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__nand2_1 _14839_ (.A(_06690_),
    .B(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__buf_2 _14840_ (.A(net7434),
    .X(_07991_));
 sky130_fd_sc_hd__o21ai_2 _14841_ (.A1(_07584_),
    .A2(_07978_),
    .B1(_07581_),
    .Y(_07992_));
 sky130_fd_sc_hd__xnor2_4 _14842_ (.A(_07984_),
    .B(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__nand2_1 _14843_ (.A(_07991_),
    .B(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__buf_2 _14844_ (.A(_06707_),
    .X(_07995_));
 sky130_fd_sc_hd__a21o_1 _14845_ (.A1(_07695_),
    .A2(_07971_),
    .B1(_07693_),
    .X(_07996_));
 sky130_fd_sc_hd__xnor2_1 _14846_ (.A(_07996_),
    .B(_07976_),
    .Y(_07997_));
 sky130_fd_sc_hd__xnor2_1 _14847_ (.A(_07584_),
    .B(_07978_),
    .Y(_07998_));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(_07997_),
    .A1(_07998_),
    .S(_06690_),
    .X(_07999_));
 sky130_fd_sc_hd__and2_1 _14849_ (.A(_07995_),
    .B(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__a31o_1 _14850_ (.A1(_06678_),
    .A2(_07990_),
    .A3(_07994_),
    .B1(_08000_),
    .X(_08001_));
 sky130_fd_sc_hd__and3_1 _14851_ (.A(net7434),
    .B(_07986_),
    .C(_07988_),
    .X(_08002_));
 sky130_fd_sc_hd__o21a_1 _14852_ (.A1(net7438),
    .A2(_08002_),
    .B1(_06707_),
    .X(_08003_));
 sky130_fd_sc_hd__nor2_1 _14853_ (.A(_06664_),
    .B(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__a21o_1 _14854_ (.A1(_06664_),
    .A2(_08001_),
    .B1(_08004_),
    .X(_08005_));
 sky130_fd_sc_hd__buf_2 _14855_ (.A(_07995_),
    .X(_08006_));
 sky130_fd_sc_hd__xor2_2 _14856_ (.A(_07695_),
    .B(_07971_),
    .X(_08007_));
 sky130_fd_sc_hd__and2_1 _14857_ (.A(net7908),
    .B(_08007_),
    .X(_08008_));
 sky130_fd_sc_hd__xnor2_1 _14858_ (.A(_07968_),
    .B(_07970_),
    .Y(_08009_));
 sky130_fd_sc_hd__nor2_1 _14859_ (.A(net7908),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__xnor2_2 _14860_ (.A(_07966_),
    .B(_07842_),
    .Y(_08011_));
 sky130_fd_sc_hd__xnor2_1 _14861_ (.A(_07967_),
    .B(_07794_),
    .Y(_08012_));
 sky130_fd_sc_hd__nor2_1 _14862_ (.A(net7434),
    .B(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__o21ba_1 _14863_ (.A1(_06690_),
    .A2(_08011_),
    .B1_N(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__nand2_1 _14864_ (.A(_08006_),
    .B(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__o31a_1 _14865_ (.A1(_08006_),
    .A2(_08008_),
    .A3(_08010_),
    .B1(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__xor2_4 _14866_ (.A(net527),
    .B(_07965_),
    .X(_08017_));
 sky130_fd_sc_hd__nor2_1 _14867_ (.A(_07881_),
    .B(_07961_),
    .Y(_08018_));
 sky130_fd_sc_hd__xnor2_2 _14868_ (.A(_07918_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__and2_1 _14869_ (.A(net7434),
    .B(_08019_),
    .X(_08020_));
 sky130_fd_sc_hd__a21o_1 _14870_ (.A1(_06690_),
    .A2(_08017_),
    .B1(_08020_),
    .X(_08021_));
 sky130_fd_sc_hd__a31o_1 _14871_ (.A1(_06664_),
    .A2(_06678_),
    .A3(_08021_),
    .B1(net7566),
    .X(_08022_));
 sky130_fd_sc_hd__a21oi_1 _14872_ (.A1(net7891),
    .A2(_08016_),
    .B1(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__a211o_1 _14873_ (.A1(net7566),
    .A2(_08005_),
    .B1(_08023_),
    .C1(_06589_),
    .X(_08024_));
 sky130_fd_sc_hd__nand2_2 _14874_ (.A(_06625_),
    .B(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__and4b_2 _14875_ (.A_N(net4931),
    .B(net4027),
    .C(_04622_),
    .D(_06207_),
    .X(_08026_));
 sky130_fd_sc_hd__buf_4 _14876_ (.A(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__mux2_1 _14877_ (.A0(net4315),
    .A1(_08025_),
    .S(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__clkbuf_1 _14878_ (.A(_08028_),
    .X(_00391_));
 sky130_fd_sc_hd__nor2_1 _14879_ (.A(net7908),
    .B(_07998_),
    .Y(_08029_));
 sky130_fd_sc_hd__a211o_1 _14880_ (.A1(_06690_),
    .A2(_07993_),
    .B1(_08029_),
    .C1(_06678_),
    .X(_08030_));
 sky130_fd_sc_hd__and3_2 _14881_ (.A(net7908),
    .B(_07986_),
    .C(_07988_),
    .X(_08031_));
 sky130_fd_sc_hd__a211o_1 _14882_ (.A1(_07991_),
    .A2(_07989_),
    .B1(_08031_),
    .C1(_06707_),
    .X(_08032_));
 sky130_fd_sc_hd__a31o_1 _14883_ (.A1(_06664_),
    .A2(_08030_),
    .A3(_08032_),
    .B1(net7457),
    .X(_08033_));
 sky130_fd_sc_hd__nand2_1 _14884_ (.A(_07991_),
    .B(_08007_),
    .Y(_08034_));
 sky130_fd_sc_hd__o21a_1 _14885_ (.A1(_07991_),
    .A2(_07997_),
    .B1(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__nor2_1 _14886_ (.A(net7434),
    .B(_08009_),
    .Y(_08036_));
 sky130_fd_sc_hd__nor2_1 _14887_ (.A(net7908),
    .B(_08012_),
    .Y(_08037_));
 sky130_fd_sc_hd__nor3_1 _14888_ (.A(_06678_),
    .B(_08036_),
    .C(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__a211o_1 _14889_ (.A1(_06678_),
    .A2(_08035_),
    .B1(_08038_),
    .C1(_06664_),
    .X(_08039_));
 sky130_fd_sc_hd__nor2_1 _14890_ (.A(net7434),
    .B(_08011_),
    .Y(_08040_));
 sky130_fd_sc_hd__a21oi_1 _14891_ (.A1(_07991_),
    .A2(_08017_),
    .B1(_08040_),
    .Y(_08041_));
 sky130_fd_sc_hd__nand2_1 _14892_ (.A(net7908),
    .B(_08019_),
    .Y(_08042_));
 sky130_fd_sc_hd__a21o_1 _14893_ (.A1(_08006_),
    .A2(_08042_),
    .B1(_06838_),
    .X(_08043_));
 sky130_fd_sc_hd__a21o_1 _14894_ (.A1(_06678_),
    .A2(_08041_),
    .B1(_08043_),
    .X(_08044_));
 sky130_fd_sc_hd__a31oi_1 _14895_ (.A1(net7568),
    .A2(_08039_),
    .A3(_08044_),
    .B1(_06589_),
    .Y(_08045_));
 sky130_fd_sc_hd__clkbuf_1 _14896_ (.A(_06626_),
    .X(_08046_));
 sky130_fd_sc_hd__clkbuf_4 _14897_ (.A(net6162),
    .X(_08047_));
 sky130_fd_sc_hd__a21o_2 _14898_ (.A1(_08033_),
    .A2(_08045_),
    .B1(_08047_),
    .X(_08048_));
 sky130_fd_sc_hd__mux2_1 _14899_ (.A0(net4310),
    .A1(_08048_),
    .S(_08027_),
    .X(_08049_));
 sky130_fd_sc_hd__clkbuf_1 _14900_ (.A(net4311),
    .X(_00392_));
 sky130_fd_sc_hd__nor3_1 _14901_ (.A(net7438),
    .B(_07995_),
    .C(_08002_),
    .Y(_08050_));
 sky130_fd_sc_hd__a311o_2 _14902_ (.A1(_07995_),
    .A2(_07990_),
    .A3(_07994_),
    .B1(_08050_),
    .C1(net7891),
    .X(_08051_));
 sky130_fd_sc_hd__nand2_1 _14903_ (.A(net7566),
    .B(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__nor2_1 _14904_ (.A(_08008_),
    .B(_08010_),
    .Y(_08053_));
 sky130_fd_sc_hd__mux2_1 _14905_ (.A0(_07999_),
    .A1(_08053_),
    .S(_07995_),
    .X(_08054_));
 sky130_fd_sc_hd__nand2_1 _14906_ (.A(_08006_),
    .B(_08021_),
    .Y(_08055_));
 sky130_fd_sc_hd__o211a_1 _14907_ (.A1(_08006_),
    .A2(_08014_),
    .B1(_08055_),
    .C1(_06663_),
    .X(_08056_));
 sky130_fd_sc_hd__a21o_1 _14908_ (.A1(_06838_),
    .A2(_08054_),
    .B1(_08056_),
    .X(_08057_));
 sky130_fd_sc_hd__nand2_1 _14909_ (.A(net7568),
    .B(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__a31o_1 _14910_ (.A1(net7433),
    .A2(_08052_),
    .A3(_08058_),
    .B1(_08047_),
    .X(_08059_));
 sky130_fd_sc_hd__mux2_1 _14911_ (.A0(net4455),
    .A1(_08059_),
    .S(_08027_),
    .X(_08060_));
 sky130_fd_sc_hd__clkbuf_1 _14912_ (.A(net4456),
    .X(_00393_));
 sky130_fd_sc_hd__a21o_1 _14913_ (.A1(_07991_),
    .A2(_07989_),
    .B1(_08031_),
    .X(_08061_));
 sky130_fd_sc_hd__a31o_1 _14914_ (.A1(_06664_),
    .A2(_08006_),
    .A3(_08061_),
    .B1(net7457),
    .X(_08062_));
 sky130_fd_sc_hd__nand2_1 _14915_ (.A(_08006_),
    .B(_08035_),
    .Y(_08063_));
 sky130_fd_sc_hd__a211o_1 _14916_ (.A1(_06690_),
    .A2(_07993_),
    .B1(_08029_),
    .C1(_07995_),
    .X(_08064_));
 sky130_fd_sc_hd__nand2_1 _14917_ (.A(_07995_),
    .B(_08041_),
    .Y(_08065_));
 sky130_fd_sc_hd__o311a_1 _14918_ (.A1(_07995_),
    .A2(_08036_),
    .A3(_08037_),
    .B1(_08065_),
    .C1(net7843),
    .X(_08066_));
 sky130_fd_sc_hd__a311o_1 _14919_ (.A1(net7891),
    .A2(_08063_),
    .A3(_08064_),
    .B1(_08066_),
    .C1(net7566),
    .X(_08067_));
 sky130_fd_sc_hd__clkbuf_4 _14920_ (.A(net7436),
    .X(_08068_));
 sky130_fd_sc_hd__buf_4 _14921_ (.A(net7771),
    .X(_08069_));
 sky130_fd_sc_hd__a21bo_1 _14922_ (.A1(net7434),
    .A2(_08017_),
    .B1_N(_08042_),
    .X(_08070_));
 sky130_fd_sc_hd__nand2_1 _14923_ (.A(_08069_),
    .B(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__nor2_1 _14924_ (.A(net7458),
    .B(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21o_1 _14925_ (.A1(_08068_),
    .A2(_08072_),
    .B1(net6162),
    .X(_08073_));
 sky130_fd_sc_hd__a31o_2 _14926_ (.A1(net7433),
    .A2(_08062_),
    .A3(_08067_),
    .B1(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__mux2_1 _14927_ (.A0(net4435),
    .A1(_08074_),
    .S(_08027_),
    .X(_08075_));
 sky130_fd_sc_hd__clkbuf_1 _14928_ (.A(_08075_),
    .X(_00394_));
 sky130_fd_sc_hd__nor2_1 _14929_ (.A(net7891),
    .B(_08016_),
    .Y(_08076_));
 sky130_fd_sc_hd__a211o_1 _14930_ (.A1(net7891),
    .A2(_08001_),
    .B1(_08076_),
    .C1(net7566),
    .X(_08077_));
 sky130_fd_sc_hd__and2_1 _14931_ (.A(net7843),
    .B(_08003_),
    .X(_08078_));
 sky130_fd_sc_hd__nand2_1 _14932_ (.A(net7566),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__a21o_1 _14933_ (.A1(_08077_),
    .A2(_08079_),
    .B1(_06589_),
    .X(_08080_));
 sky130_fd_sc_hd__nand2_1 _14934_ (.A(net7908),
    .B(_08017_),
    .Y(_08081_));
 sky130_fd_sc_hd__o21ai_1 _14935_ (.A1(net7908),
    .A2(_08011_),
    .B1(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__mux2_1 _14936_ (.A0(_08020_),
    .A1(_08082_),
    .S(_08069_),
    .X(_08083_));
 sky130_fd_sc_hd__and2_1 _14937_ (.A(net7759),
    .B(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__a21oi_1 _14938_ (.A1(_08068_),
    .A2(_08084_),
    .B1(_08047_),
    .Y(_08085_));
 sky130_fd_sc_hd__nand2_2 _14939_ (.A(_08080_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__mux2_1 _14940_ (.A0(net4382),
    .A1(_08086_),
    .S(_08027_),
    .X(_08087_));
 sky130_fd_sc_hd__clkbuf_1 _14941_ (.A(_08087_),
    .X(_00395_));
 sky130_fd_sc_hd__a21o_1 _14942_ (.A1(_08030_),
    .A2(_08032_),
    .B1(net7843),
    .X(_08088_));
 sky130_fd_sc_hd__a21o_1 _14943_ (.A1(_06678_),
    .A2(_08035_),
    .B1(_08038_),
    .X(_08089_));
 sky130_fd_sc_hd__nand2_1 _14944_ (.A(net7433),
    .B(net7457),
    .Y(_08090_));
 sky130_fd_sc_hd__a21oi_1 _14945_ (.A1(_06664_),
    .A2(_08089_),
    .B1(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__clkbuf_4 _14946_ (.A(net7759),
    .X(_08092_));
 sky130_fd_sc_hd__or2_1 _14947_ (.A(_08037_),
    .B(_08040_),
    .X(_08093_));
 sky130_fd_sc_hd__mux2_1 _14948_ (.A0(_08070_),
    .A1(_08093_),
    .S(_08069_),
    .X(_08094_));
 sky130_fd_sc_hd__and2_1 _14949_ (.A(_08092_),
    .B(_08094_),
    .X(_08095_));
 sky130_fd_sc_hd__a221o_2 _14950_ (.A1(_08088_),
    .A2(_08091_),
    .B1(_08095_),
    .B2(_08068_),
    .C1(net6162),
    .X(_08096_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(net4374),
    .A1(_08096_),
    .S(_08027_),
    .X(_08097_));
 sky130_fd_sc_hd__clkbuf_1 _14952_ (.A(_08097_),
    .X(_00396_));
 sky130_fd_sc_hd__a31o_1 _14953_ (.A1(_08006_),
    .A2(_07990_),
    .A3(_07994_),
    .B1(_08050_),
    .X(_08098_));
 sky130_fd_sc_hd__a21o_1 _14954_ (.A1(_06664_),
    .A2(_08054_),
    .B1(_08090_),
    .X(_08099_));
 sky130_fd_sc_hd__a21o_1 _14955_ (.A1(net7891),
    .A2(_08098_),
    .B1(_08099_),
    .X(_08100_));
 sky130_fd_sc_hd__or2_1 _14956_ (.A(_08013_),
    .B(_08010_),
    .X(_08101_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(_08082_),
    .A1(_08101_),
    .S(_08069_),
    .X(_08102_));
 sky130_fd_sc_hd__and3_1 _14958_ (.A(_07995_),
    .B(_07991_),
    .C(_08019_),
    .X(_08103_));
 sky130_fd_sc_hd__mux2_1 _14959_ (.A0(_08102_),
    .A1(_08103_),
    .S(net7458),
    .X(_08104_));
 sky130_fd_sc_hd__a21oi_1 _14960_ (.A1(_08068_),
    .A2(_08104_),
    .B1(net6162),
    .Y(_08105_));
 sky130_fd_sc_hd__nand2_2 _14961_ (.A(_08100_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(net4473),
    .A1(_08106_),
    .S(_08027_),
    .X(_08107_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_08107_),
    .X(_00397_));
 sky130_fd_sc_hd__inv_2 _14964_ (.A(_08090_),
    .Y(_08108_));
 sky130_fd_sc_hd__a21o_1 _14965_ (.A1(_08006_),
    .A2(_08061_),
    .B1(_06664_),
    .X(_08109_));
 sky130_fd_sc_hd__a21o_1 _14966_ (.A1(_08063_),
    .A2(_08064_),
    .B1(net7891),
    .X(_08110_));
 sky130_fd_sc_hd__a21o_1 _14967_ (.A1(_07991_),
    .A2(_08007_),
    .B1(_08036_),
    .X(_08111_));
 sky130_fd_sc_hd__nand2_1 _14968_ (.A(_08069_),
    .B(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand2_1 _14969_ (.A(_06721_),
    .B(_08093_),
    .Y(_08113_));
 sky130_fd_sc_hd__and2_1 _14970_ (.A(net7458),
    .B(_08071_),
    .X(_08114_));
 sky130_fd_sc_hd__a31oi_2 _14971_ (.A1(_08092_),
    .A2(_08112_),
    .A3(_08113_),
    .B1(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__a21o_1 _14972_ (.A1(_08068_),
    .A2(_08115_),
    .B1(net6162),
    .X(_08116_));
 sky130_fd_sc_hd__a31o_2 _14973_ (.A1(_08108_),
    .A2(_08109_),
    .A3(_08110_),
    .B1(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__mux2_1 _14974_ (.A0(net4353),
    .A1(_08117_),
    .S(_08027_),
    .X(_08118_));
 sky130_fd_sc_hd__clkbuf_1 _14975_ (.A(net4354),
    .X(_00398_));
 sky130_fd_sc_hd__a211o_1 _14976_ (.A1(_06664_),
    .A2(_08001_),
    .B1(_08004_),
    .C1(_08090_),
    .X(_08119_));
 sky130_fd_sc_hd__xnor2_1 _14977_ (.A(_07996_),
    .B(_07975_),
    .Y(_08120_));
 sky130_fd_sc_hd__a21o_1 _14978_ (.A1(_07991_),
    .A2(_08120_),
    .B1(_08008_),
    .X(_08121_));
 sky130_fd_sc_hd__mux2_1 _14979_ (.A0(_08101_),
    .A1(_08121_),
    .S(_08069_),
    .X(_08122_));
 sky130_fd_sc_hd__mux2_1 _14980_ (.A0(_08083_),
    .A1(_08122_),
    .S(_08092_),
    .X(_08123_));
 sky130_fd_sc_hd__a21oi_1 _14981_ (.A1(_08068_),
    .A2(_08123_),
    .B1(net6162),
    .Y(_08124_));
 sky130_fd_sc_hd__nand2_1 _14982_ (.A(net7439),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__mux2_1 _14983_ (.A0(net3505),
    .A1(_08125_),
    .S(_08027_),
    .X(_08126_));
 sky130_fd_sc_hd__clkbuf_1 _14984_ (.A(_08126_),
    .X(_00399_));
 sky130_fd_sc_hd__and3_1 _14985_ (.A(_06663_),
    .B(_08030_),
    .C(_08032_),
    .X(_08127_));
 sky130_fd_sc_hd__a21o_1 _14986_ (.A1(_06690_),
    .A2(_08120_),
    .B1(_08029_),
    .X(_08128_));
 sky130_fd_sc_hd__mux4_2 _14987_ (.A0(_08070_),
    .A1(_08093_),
    .A2(_08111_),
    .A3(_08128_),
    .S0(_08069_),
    .S1(net7759),
    .X(_08129_));
 sky130_fd_sc_hd__a221o_4 _14988_ (.A1(_08127_),
    .A2(_08108_),
    .B1(_08129_),
    .B2(net7436),
    .C1(net6162),
    .X(_08130_));
 sky130_fd_sc_hd__mux2_1 _14989_ (.A0(net4393),
    .A1(net7437),
    .S(_08027_),
    .X(_08131_));
 sky130_fd_sc_hd__clkbuf_1 _14990_ (.A(_08131_),
    .X(_00400_));
 sky130_fd_sc_hd__xnor2_1 _14991_ (.A(_07583_),
    .B(_07978_),
    .Y(_08132_));
 sky130_fd_sc_hd__mux4_2 _14992_ (.A0(_08120_),
    .A1(_08132_),
    .A2(_07993_),
    .A3(_08007_),
    .S0(_06690_),
    .S1(_06707_),
    .X(_08133_));
 sky130_fd_sc_hd__nand2_1 _14993_ (.A(net7458),
    .B(_08102_),
    .Y(_08134_));
 sky130_fd_sc_hd__a21boi_2 _14994_ (.A1(_08092_),
    .A2(_08133_),
    .B1_N(_08134_),
    .Y(_08135_));
 sky130_fd_sc_hd__a21oi_1 _14995_ (.A1(_06734_),
    .A2(_08103_),
    .B1(net3457),
    .Y(_08136_));
 sky130_fd_sc_hd__o221ai_4 _14996_ (.A1(net7566),
    .A2(_08051_),
    .B1(_08135_),
    .B2(net7836),
    .C1(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__buf_4 _14997_ (.A(_08026_),
    .X(_08138_));
 sky130_fd_sc_hd__mux2_1 _14998_ (.A0(net4405),
    .A1(_08137_),
    .S(_08138_),
    .X(_08139_));
 sky130_fd_sc_hd__clkbuf_1 _14999_ (.A(_08139_),
    .X(_00401_));
 sky130_fd_sc_hd__and3_1 _15000_ (.A(net7843),
    .B(_07995_),
    .C(_08061_),
    .X(_08140_));
 sky130_fd_sc_hd__mux2_4 _15001_ (.A0(_07989_),
    .A1(_07993_),
    .S(_06690_),
    .X(_08141_));
 sky130_fd_sc_hd__mux4_2 _15002_ (.A0(_08093_),
    .A1(_08111_),
    .A2(_08128_),
    .A3(_08141_),
    .S0(_08069_),
    .S1(net7759),
    .X(_08142_));
 sky130_fd_sc_hd__a21o_1 _15003_ (.A1(_06734_),
    .A2(_08072_),
    .B1(net3457),
    .X(_08143_));
 sky130_fd_sc_hd__a221o_2 _15004_ (.A1(net7457),
    .A2(_08140_),
    .B1(_08142_),
    .B2(net7436),
    .C1(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__mux2_1 _15005_ (.A0(net4451),
    .A1(_08144_),
    .S(_08138_),
    .X(_08145_));
 sky130_fd_sc_hd__clkbuf_1 _15006_ (.A(_08145_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _15007_ (.A0(_08132_),
    .A1(_07993_),
    .S(_07991_),
    .X(_08146_));
 sky130_fd_sc_hd__a21o_1 _15008_ (.A1(_06690_),
    .A2(_07989_),
    .B1(_08002_),
    .X(_08147_));
 sky130_fd_sc_hd__mux2_1 _15009_ (.A0(_08146_),
    .A1(_08147_),
    .S(_08069_),
    .X(_08148_));
 sky130_fd_sc_hd__mux2_2 _15010_ (.A0(_08122_),
    .A1(_08148_),
    .S(_08092_),
    .X(_08149_));
 sky130_fd_sc_hd__clkbuf_4 _15011_ (.A(_06734_),
    .X(_08150_));
 sky130_fd_sc_hd__a221o_1 _15012_ (.A1(net7457),
    .A2(_08078_),
    .B1(_08084_),
    .B2(_08150_),
    .C1(net6162),
    .X(_08151_));
 sky130_fd_sc_hd__a21o_4 _15013_ (.A1(_08068_),
    .A2(_08149_),
    .B1(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__mux2_1 _15014_ (.A0(net4372),
    .A1(_08152_),
    .S(_08138_),
    .X(_08153_));
 sky130_fd_sc_hd__clkbuf_1 _15015_ (.A(_08153_),
    .X(_00403_));
 sky130_fd_sc_hd__mux4_1 _15016_ (.A0(_08031_),
    .A1(_08128_),
    .A2(_08141_),
    .A3(_08111_),
    .S0(net7458),
    .S1(net7478),
    .X(_08154_));
 sky130_fd_sc_hd__a221o_4 _15017_ (.A1(_08150_),
    .A2(_08095_),
    .B1(_08154_),
    .B2(_08068_),
    .C1(net6162),
    .X(_08155_));
 sky130_fd_sc_hd__mux2_1 _15018_ (.A0(net4423),
    .A1(_08155_),
    .S(_08138_),
    .X(_08156_));
 sky130_fd_sc_hd__clkbuf_1 _15019_ (.A(_08156_),
    .X(_00404_));
 sky130_fd_sc_hd__and2_1 _15020_ (.A(net7478),
    .B(_08147_),
    .X(_08157_));
 sky130_fd_sc_hd__or2_1 _15021_ (.A(net7759),
    .B(_08133_),
    .X(_08158_));
 sky130_fd_sc_hd__o211a_1 _15022_ (.A1(net7458),
    .A2(_08157_),
    .B1(_08158_),
    .C1(_08068_),
    .X(_08159_));
 sky130_fd_sc_hd__a211o_2 _15023_ (.A1(_08150_),
    .A2(_08104_),
    .B1(_08159_),
    .C1(net6162),
    .X(_08160_));
 sky130_fd_sc_hd__mux2_1 _15024_ (.A0(net4378),
    .A1(_08160_),
    .S(_08138_),
    .X(_08161_));
 sky130_fd_sc_hd__clkbuf_1 _15025_ (.A(_08161_),
    .X(_00405_));
 sky130_fd_sc_hd__inv_2 _15026_ (.A(net5684),
    .Y(_08162_));
 sky130_fd_sc_hd__mux2_1 _15027_ (.A0(_08128_),
    .A1(_08141_),
    .S(_08069_),
    .X(_08163_));
 sky130_fd_sc_hd__nand2_1 _15028_ (.A(_08006_),
    .B(_08031_),
    .Y(_08164_));
 sky130_fd_sc_hd__a21oi_1 _15029_ (.A1(_08092_),
    .A2(_08164_),
    .B1(net7836),
    .Y(_08165_));
 sky130_fd_sc_hd__o21ai_2 _15030_ (.A1(_08092_),
    .A2(_08163_),
    .B1(_08165_),
    .Y(_08166_));
 sky130_fd_sc_hd__a21oi_2 _15031_ (.A1(_08150_),
    .A2(_08115_),
    .B1(_08047_),
    .Y(_08167_));
 sky130_fd_sc_hd__and2_1 _15032_ (.A(_08166_),
    .B(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__mux2_1 _15033_ (.A0(net3064),
    .A1(_08168_),
    .S(_08026_),
    .X(_08169_));
 sky130_fd_sc_hd__inv_2 _15034_ (.A(net5686),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _15035_ (.A(net7757),
    .B(_08092_),
    .Y(_08170_));
 sky130_fd_sc_hd__o211a_1 _15036_ (.A1(_08092_),
    .A2(_08148_),
    .B1(net7430),
    .C1(_06715_),
    .X(_08171_));
 sky130_fd_sc_hd__a31o_1 _15037_ (.A1(net7431),
    .A2(_06714_),
    .A3(_08123_),
    .B1(_08171_),
    .X(_08172_));
 sky130_fd_sc_hd__a21o_2 _15038_ (.A1(_06589_),
    .A2(_08172_),
    .B1(_08047_),
    .X(_08173_));
 sky130_fd_sc_hd__mux2_1 _15039_ (.A0(net4368),
    .A1(_08173_),
    .S(_08138_),
    .X(_08174_));
 sky130_fd_sc_hd__clkbuf_1 _15040_ (.A(_08174_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _15041_ (.A0(_08031_),
    .A1(_08141_),
    .S(net7478),
    .X(_08175_));
 sky130_fd_sc_hd__nor2_2 _15042_ (.A(_08092_),
    .B(net7836),
    .Y(_08176_));
 sky130_fd_sc_hd__a221o_2 _15043_ (.A1(_08150_),
    .A2(_08129_),
    .B1(_08175_),
    .B2(_08176_),
    .C1(_08047_),
    .X(_08177_));
 sky130_fd_sc_hd__mux2_1 _15044_ (.A0(net4386),
    .A1(_08177_),
    .S(_08138_),
    .X(_08178_));
 sky130_fd_sc_hd__clkbuf_1 _15045_ (.A(_08178_),
    .X(_00408_));
 sky130_fd_sc_hd__nand2_1 _15046_ (.A(_08157_),
    .B(_08176_),
    .Y(_08179_));
 sky130_fd_sc_hd__o311a_2 _15047_ (.A1(net7433),
    .A2(_06715_),
    .A3(_08135_),
    .B1(_08179_),
    .C1(_06625_),
    .X(_08180_));
 sky130_fd_sc_hd__inv_2 _15048_ (.A(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__mux2_1 _15049_ (.A0(net4431),
    .A1(_08181_),
    .S(_08138_),
    .X(_08182_));
 sky130_fd_sc_hd__clkbuf_1 _15050_ (.A(_08182_),
    .X(_00409_));
 sky130_fd_sc_hd__inv_2 _15051_ (.A(_08164_),
    .Y(_08183_));
 sky130_fd_sc_hd__a221o_1 _15052_ (.A1(_08150_),
    .A2(_08142_),
    .B1(_08183_),
    .B2(_08176_),
    .C1(_08047_),
    .X(_08184_));
 sky130_fd_sc_hd__mux2_1 _15053_ (.A0(net4380),
    .A1(_08184_),
    .S(_08138_),
    .X(_08185_));
 sky130_fd_sc_hd__clkbuf_1 _15054_ (.A(_08185_),
    .X(_00410_));
 sky130_fd_sc_hd__a21o_1 _15055_ (.A1(_08150_),
    .A2(_08149_),
    .B1(_08047_),
    .X(_08186_));
 sky130_fd_sc_hd__mux2_1 _15056_ (.A0(net4586),
    .A1(_08186_),
    .S(_08138_),
    .X(_08187_));
 sky130_fd_sc_hd__clkbuf_1 _15057_ (.A(_08187_),
    .X(_00411_));
 sky130_fd_sc_hd__and3_1 _15058_ (.A(_06625_),
    .B(_08150_),
    .C(_08154_),
    .X(_08188_));
 sky130_fd_sc_hd__mux2_1 _15059_ (.A0(net4332),
    .A1(_08188_),
    .S(_08026_),
    .X(_08189_));
 sky130_fd_sc_hd__clkbuf_1 _15060_ (.A(_08189_),
    .X(_00412_));
 sky130_fd_sc_hd__clkbuf_4 _15061_ (.A(_06386_),
    .X(_08190_));
 sky130_fd_sc_hd__clkbuf_4 _15062_ (.A(_06344_),
    .X(_08191_));
 sky130_fd_sc_hd__mux2_1 _15063_ (.A0(net4568),
    .A1(net4475),
    .S(_08191_),
    .X(_08192_));
 sky130_fd_sc_hd__inv_2 _15064_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .Y(_08193_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(net3722),
    .B(_06386_),
    .Y(_08194_));
 sky130_fd_sc_hd__clkbuf_8 _15066_ (.A(_04624_),
    .X(_08195_));
 sky130_fd_sc_hd__clkbuf_4 _15067_ (.A(_08195_),
    .X(_01622_));
 sky130_fd_sc_hd__o211a_1 _15068_ (.A1(_08190_),
    .A2(_08192_),
    .B1(net3723),
    .C1(_01622_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _15069_ (.A0(net4507),
    .A1(net4467),
    .S(_08191_),
    .X(_08196_));
 sky130_fd_sc_hd__inv_2 _15070_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_08197_));
 sky130_fd_sc_hd__nand2_1 _15071_ (.A(net3539),
    .B(_06386_),
    .Y(_08198_));
 sky130_fd_sc_hd__o211a_1 _15072_ (.A1(_08190_),
    .A2(_08196_),
    .B1(net3540),
    .C1(_01622_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _15073_ (.A0(net4689),
    .A1(net4687),
    .S(_08191_),
    .X(_08199_));
 sky130_fd_sc_hd__nor2_2 _15074_ (.A(_06203_),
    .B(_06384_),
    .Y(_08200_));
 sky130_fd_sc_hd__buf_2 _15075_ (.A(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__or2_1 _15076_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_08201_),
    .X(_08202_));
 sky130_fd_sc_hd__o211a_1 _15077_ (.A1(_08190_),
    .A2(_08199_),
    .B1(net6139),
    .C1(_01622_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _15078_ (.A0(net4528),
    .A1(net4499),
    .S(_08191_),
    .X(_08203_));
 sky130_fd_sc_hd__or2_1 _15079_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08201_),
    .X(_08204_));
 sky130_fd_sc_hd__o211a_1 _15080_ (.A1(_08190_),
    .A2(_08203_),
    .B1(net6092),
    .C1(_01622_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _15081_ (.A0(net4597),
    .A1(net4591),
    .S(_08191_),
    .X(_08205_));
 sky130_fd_sc_hd__or2_1 _15082_ (.A(net3206),
    .B(_08201_),
    .X(_08206_));
 sky130_fd_sc_hd__o211a_1 _15083_ (.A1(_08190_),
    .A2(_08205_),
    .B1(net3207),
    .C1(_01622_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _15084_ (.A0(net4556),
    .A1(net4511),
    .S(_08191_),
    .X(_08207_));
 sky130_fd_sc_hd__or2_1 _15085_ (.A(net3356),
    .B(_08201_),
    .X(_08208_));
 sky130_fd_sc_hd__o211a_1 _15086_ (.A1(_08190_),
    .A2(_08207_),
    .B1(net3357),
    .C1(_01622_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _15087_ (.A0(net4560),
    .A1(net4491),
    .S(_08191_),
    .X(_08209_));
 sky130_fd_sc_hd__or2_1 _15088_ (.A(net3262),
    .B(_08201_),
    .X(_08210_));
 sky130_fd_sc_hd__o211a_1 _15089_ (.A1(_08190_),
    .A2(_08209_),
    .B1(net3263),
    .C1(_01622_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _15090_ (.A0(net3462),
    .A1(net3284),
    .S(_08191_),
    .X(_08211_));
 sky130_fd_sc_hd__or2_1 _15091_ (.A(net645),
    .B(_08201_),
    .X(_08212_));
 sky130_fd_sc_hd__o211a_1 _15092_ (.A1(_08190_),
    .A2(net3463),
    .B1(net6204),
    .C1(_01622_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _15093_ (.A0(net3200),
    .A1(net3184),
    .S(_08191_),
    .X(_08213_));
 sky130_fd_sc_hd__or2_1 _15094_ (.A(net6253),
    .B(_08201_),
    .X(_08214_));
 sky130_fd_sc_hd__buf_2 _15095_ (.A(_08195_),
    .X(_08215_));
 sky130_fd_sc_hd__o211a_1 _15096_ (.A1(_08190_),
    .A2(net3201),
    .B1(net6254),
    .C1(_08215_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _15097_ (.A0(net3417),
    .A1(net3221),
    .S(_08191_),
    .X(_08216_));
 sky130_fd_sc_hd__or2_1 _15098_ (.A(net6278),
    .B(_08201_),
    .X(_08217_));
 sky130_fd_sc_hd__o211a_1 _15099_ (.A1(_08190_),
    .A2(net3067),
    .B1(net6279),
    .C1(_08215_),
    .X(_00422_));
 sky130_fd_sc_hd__buf_2 _15100_ (.A(_06386_),
    .X(_08218_));
 sky130_fd_sc_hd__clkbuf_4 _15101_ (.A(_06344_),
    .X(_08219_));
 sky130_fd_sc_hd__mux2_1 _15102_ (.A0(net3047),
    .A1(net3233),
    .S(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__or2_1 _15103_ (.A(net6281),
    .B(_08201_),
    .X(_08221_));
 sky130_fd_sc_hd__o211a_1 _15104_ (.A1(_08218_),
    .A2(net3048),
    .B1(net6282),
    .C1(_08215_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _15105_ (.A0(net3186),
    .A1(net3174),
    .S(_08219_),
    .X(_08222_));
 sky130_fd_sc_hd__clkbuf_2 _15106_ (.A(_08200_),
    .X(_08223_));
 sky130_fd_sc_hd__or2_1 _15107_ (.A(net6259),
    .B(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__o211a_1 _15108_ (.A1(_08218_),
    .A2(net3187),
    .B1(net6260),
    .C1(_08215_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _15109_ (.A0(net3460),
    .A1(net3054),
    .S(_08219_),
    .X(_08225_));
 sky130_fd_sc_hd__or2_1 _15110_ (.A(net4783),
    .B(_08223_),
    .X(_08226_));
 sky130_fd_sc_hd__o211a_1 _15111_ (.A1(_08218_),
    .A2(net3055),
    .B1(net4784),
    .C1(_08215_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _15112_ (.A0(net3166),
    .A1(net3314),
    .S(_08219_),
    .X(_08227_));
 sky130_fd_sc_hd__or2_1 _15113_ (.A(net4581),
    .B(_08223_),
    .X(_08228_));
 sky130_fd_sc_hd__o211a_1 _15114_ (.A1(_08218_),
    .A2(net3167),
    .B1(net4582),
    .C1(_08215_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _15115_ (.A0(net4501),
    .A1(net4613),
    .S(_08219_),
    .X(_08229_));
 sky130_fd_sc_hd__or2_1 _15116_ (.A(net6123),
    .B(_08223_),
    .X(_08230_));
 sky130_fd_sc_hd__o211a_1 _15117_ (.A1(_08218_),
    .A2(_08229_),
    .B1(net3631),
    .C1(_08215_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _15118_ (.A0(net4403),
    .A1(net4458),
    .S(_08219_),
    .X(_08231_));
 sky130_fd_sc_hd__or2_1 _15119_ (.A(net6098),
    .B(_08223_),
    .X(_08232_));
 sky130_fd_sc_hd__o211a_1 _15120_ (.A1(_08218_),
    .A2(_08231_),
    .B1(net3223),
    .C1(_08215_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _15121_ (.A0(net4433),
    .A1(net4483),
    .S(_08219_),
    .X(_08233_));
 sky130_fd_sc_hd__or2_1 _15122_ (.A(net6148),
    .B(_08223_),
    .X(_08234_));
 sky130_fd_sc_hd__o211a_1 _15123_ (.A1(_08218_),
    .A2(_08233_),
    .B1(net3628),
    .C1(_08215_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _15124_ (.A0(net4558),
    .A1(net4573),
    .S(_08219_),
    .X(_08235_));
 sky130_fd_sc_hd__or2_1 _15125_ (.A(net6150),
    .B(_08223_),
    .X(_08236_));
 sky130_fd_sc_hd__o211a_1 _15126_ (.A1(_08218_),
    .A2(_08235_),
    .B1(net3719),
    .C1(_08215_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(net4599),
    .A1(net4513),
    .S(_08219_),
    .X(_08237_));
 sky130_fd_sc_hd__or2_1 _15128_ (.A(net6146),
    .B(_08223_),
    .X(_08238_));
 sky130_fd_sc_hd__buf_4 _15129_ (.A(_08195_),
    .X(_08239_));
 sky130_fd_sc_hd__o211a_1 _15130_ (.A1(_08218_),
    .A2(_08237_),
    .B1(net3773),
    .C1(_08239_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _15131_ (.A0(net4497),
    .A1(net4437),
    .S(_08219_),
    .X(_08240_));
 sky130_fd_sc_hd__or2_1 _15132_ (.A(net6134),
    .B(_08223_),
    .X(_08241_));
 sky130_fd_sc_hd__o211a_1 _15133_ (.A1(_08218_),
    .A2(_08240_),
    .B1(net6136),
    .C1(_08239_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _15134_ (.A0(net3691),
    .A1(net3058),
    .S(_06344_),
    .X(_08242_));
 sky130_fd_sc_hd__or2_1 _15135_ (.A(net4779),
    .B(_08223_),
    .X(_08243_));
 sky130_fd_sc_hd__o211a_1 _15136_ (.A1(_06386_),
    .A2(net3692),
    .B1(net4780),
    .C1(_08239_),
    .X(_00433_));
 sky130_fd_sc_hd__o21a_1 _15137_ (.A1(net4577),
    .A2(_06343_),
    .B1(net4342),
    .X(_08244_));
 sky130_fd_sc_hd__nand2_1 _15138_ (.A(net4828),
    .B(_06386_),
    .Y(_08245_));
 sky130_fd_sc_hd__o211a_1 _15139_ (.A1(_06386_),
    .A2(net2960),
    .B1(net4829),
    .C1(_08239_),
    .X(_00434_));
 sky130_fd_sc_hd__buf_4 _15140_ (.A(_04621_),
    .X(_08246_));
 sky130_fd_sc_hd__or4b_1 _15141_ (.A(net4909),
    .B(net2982),
    .C(net4027),
    .D_N(net4931),
    .X(_08247_));
 sky130_fd_sc_hd__nor2_1 _15142_ (.A(_08246_),
    .B(net4932),
    .Y(_08248_));
 sky130_fd_sc_hd__buf_4 _15143_ (.A(net4933),
    .X(_08249_));
 sky130_fd_sc_hd__mux2_1 _15144_ (.A0(net4566),
    .A1(_08025_),
    .S(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__clkbuf_1 _15145_ (.A(_08250_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _15146_ (.A0(net4579),
    .A1(_08048_),
    .S(_08249_),
    .X(_08251_));
 sky130_fd_sc_hd__clkbuf_1 _15147_ (.A(net4580),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _15148_ (.A0(net4570),
    .A1(_08059_),
    .S(_08249_),
    .X(_08252_));
 sky130_fd_sc_hd__clkbuf_1 _15149_ (.A(net4571),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _15150_ (.A0(net4727),
    .A1(_08074_),
    .S(_08249_),
    .X(_08253_));
 sky130_fd_sc_hd__clkbuf_1 _15151_ (.A(_08253_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _15152_ (.A0(net4370),
    .A1(_08086_),
    .S(_08249_),
    .X(_08254_));
 sky130_fd_sc_hd__clkbuf_1 _15153_ (.A(_08254_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _15154_ (.A0(net4719),
    .A1(_08096_),
    .S(_08249_),
    .X(_08255_));
 sky130_fd_sc_hd__clkbuf_1 _15155_ (.A(_08255_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _15156_ (.A0(net4399),
    .A1(_08106_),
    .S(_08249_),
    .X(_08256_));
 sky130_fd_sc_hd__clkbuf_1 _15157_ (.A(_08256_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(net4716),
    .A1(_08117_),
    .S(_08249_),
    .X(_08257_));
 sky130_fd_sc_hd__clkbuf_1 _15159_ (.A(net4717),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _15160_ (.A0(net3419),
    .A1(_08125_),
    .S(_08249_),
    .X(_08258_));
 sky130_fd_sc_hd__clkbuf_1 _15161_ (.A(_08258_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _15162_ (.A0(net4714),
    .A1(net7437),
    .S(_08249_),
    .X(_08259_));
 sky130_fd_sc_hd__clkbuf_1 _15163_ (.A(_08259_),
    .X(_00444_));
 sky130_fd_sc_hd__buf_4 _15164_ (.A(net4933),
    .X(_08260_));
 sky130_fd_sc_hd__mux2_1 _15165_ (.A0(net4362),
    .A1(_08137_),
    .S(_08260_),
    .X(_08261_));
 sky130_fd_sc_hd__clkbuf_1 _15166_ (.A(_08261_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _15167_ (.A0(net4334),
    .A1(_08144_),
    .S(_08260_),
    .X(_08262_));
 sky130_fd_sc_hd__clkbuf_1 _15168_ (.A(_08262_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _15169_ (.A0(net4411),
    .A1(_08152_),
    .S(_08260_),
    .X(_08263_));
 sky130_fd_sc_hd__clkbuf_1 _15170_ (.A(_08263_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _15171_ (.A0(net4349),
    .A1(_08155_),
    .S(_08260_),
    .X(_08264_));
 sky130_fd_sc_hd__clkbuf_1 _15172_ (.A(_08264_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _15173_ (.A0(net4417),
    .A1(_08160_),
    .S(_08260_),
    .X(_08265_));
 sky130_fd_sc_hd__clkbuf_1 _15174_ (.A(_08265_),
    .X(_00449_));
 sky130_fd_sc_hd__inv_2 _15175_ (.A(net3272),
    .Y(_08266_));
 sky130_fd_sc_hd__mux2_1 _15176_ (.A0(net3273),
    .A1(_08168_),
    .S(net4933),
    .X(_08267_));
 sky130_fd_sc_hd__inv_2 _15177_ (.A(net4934),
    .Y(_00450_));
 sky130_fd_sc_hd__mux2_1 _15178_ (.A0(net4593),
    .A1(_08173_),
    .S(_08260_),
    .X(_08268_));
 sky130_fd_sc_hd__clkbuf_1 _15179_ (.A(_08268_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _15180_ (.A0(net4639),
    .A1(_08177_),
    .S(_08260_),
    .X(_08269_));
 sky130_fd_sc_hd__clkbuf_1 _15181_ (.A(_08269_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _15182_ (.A0(net4530),
    .A1(_08181_),
    .S(_08260_),
    .X(_08270_));
 sky130_fd_sc_hd__clkbuf_1 _15183_ (.A(_08270_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _15184_ (.A0(net4619),
    .A1(_08184_),
    .S(_08260_),
    .X(_08271_));
 sky130_fd_sc_hd__clkbuf_1 _15185_ (.A(_08271_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _15186_ (.A0(net4605),
    .A1(_08186_),
    .S(_08260_),
    .X(_08272_));
 sky130_fd_sc_hd__clkbuf_1 _15187_ (.A(_08272_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _15188_ (.A0(net4575),
    .A1(_08188_),
    .S(net4933),
    .X(_08273_));
 sky130_fd_sc_hd__clkbuf_1 _15189_ (.A(_08273_),
    .X(_00456_));
 sky130_fd_sc_hd__buf_4 _15190_ (.A(net89),
    .X(_08274_));
 sky130_fd_sc_hd__buf_4 _15191_ (.A(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__buf_4 _15192_ (.A(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__and2_1 _15193_ (.A(_08276_),
    .B(net4095),
    .X(_08277_));
 sky130_fd_sc_hd__clkbuf_1 _15194_ (.A(net4096),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _15195_ (.A(net65),
    .B(net4007),
    .Y(_00458_));
 sky130_fd_sc_hd__and2_1 _15196_ (.A(_08276_),
    .B(net4045),
    .X(_08278_));
 sky130_fd_sc_hd__clkbuf_1 _15197_ (.A(net4046),
    .X(_00459_));
 sky130_fd_sc_hd__buf_4 _15198_ (.A(_08275_),
    .X(_08279_));
 sky130_fd_sc_hd__and2_1 _15199_ (.A(_08279_),
    .B(net4066),
    .X(_08280_));
 sky130_fd_sc_hd__clkbuf_1 _15200_ (.A(net4067),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _15201_ (.A(_08279_),
    .B(net4083),
    .X(_08281_));
 sky130_fd_sc_hd__clkbuf_1 _15202_ (.A(net4084),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _15203_ (.A(_08279_),
    .B(net4078),
    .X(_08282_));
 sky130_fd_sc_hd__clkbuf_1 _15204_ (.A(net4079),
    .X(_00462_));
 sky130_fd_sc_hd__o21bai_1 _15205_ (.A1(_06382_),
    .A2(_06359_),
    .B1_N(_06267_),
    .Y(_08283_));
 sky130_fd_sc_hd__a2bb2o_1 _15206_ (.A1_N(_06381_),
    .A2_N(_08283_),
    .B1(_06267_),
    .B2(net1054),
    .X(_08284_));
 sky130_fd_sc_hd__mux2_1 _15207_ (.A0(_08284_),
    .A1(net1068),
    .S(net3622),
    .X(_08285_));
 sky130_fd_sc_hd__and2_1 _15208_ (.A(net3508),
    .B(_06384_),
    .X(_08286_));
 sky130_fd_sc_hd__mux2_1 _15209_ (.A0(_04693_),
    .A1(net3623),
    .S(net3509),
    .X(_08287_));
 sky130_fd_sc_hd__and2_1 _15210_ (.A(_08195_),
    .B(net3624),
    .X(_08288_));
 sky130_fd_sc_hd__clkbuf_1 _15211_ (.A(net3625),
    .X(_00463_));
 sky130_fd_sc_hd__a2bb2o_1 _15212_ (.A1_N(_06367_),
    .A2_N(_08283_),
    .B1(_06267_),
    .B2(net1312),
    .X(_08289_));
 sky130_fd_sc_hd__mux2_1 _15213_ (.A0(_08289_),
    .A1(net1008),
    .S(_06258_),
    .X(_08290_));
 sky130_fd_sc_hd__mux2_1 _15214_ (.A0(_04692_),
    .A1(_08290_),
    .S(net3509),
    .X(_08291_));
 sky130_fd_sc_hd__and2_1 _15215_ (.A(_08195_),
    .B(net3510),
    .X(_08292_));
 sky130_fd_sc_hd__clkbuf_1 _15216_ (.A(net3511),
    .X(_00464_));
 sky130_fd_sc_hd__buf_4 _15217_ (.A(net4087),
    .X(_08293_));
 sky130_fd_sc_hd__o211a_1 _15218_ (.A1(net4088),
    .A2(_08201_),
    .B1(_06387_),
    .C1(_08239_),
    .X(_00465_));
 sky130_fd_sc_hd__nor2_2 _15219_ (.A(net3507),
    .B(_04818_),
    .Y(_08294_));
 sky130_fd_sc_hd__clkbuf_4 _15220_ (.A(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__buf_4 _15221_ (.A(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__nand2b_4 _15222_ (.A_N(net3535),
    .B(_06207_),
    .Y(_08297_));
 sky130_fd_sc_hd__clkbuf_8 _15223_ (.A(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__clkbuf_8 _15224_ (.A(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__clkbuf_4 _15225_ (.A(net4086),
    .X(_08300_));
 sky130_fd_sc_hd__mux2_1 _15226_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__mux2_2 _15227_ (.A0(_08048_),
    .A1(net7464),
    .S(_08295_),
    .X(_08302_));
 sky130_fd_sc_hd__and3_2 _15228_ (.A(net3506),
    .B(net3534),
    .C(_06207_),
    .X(_08303_));
 sky130_fd_sc_hd__buf_4 _15229_ (.A(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__clkbuf_8 _15230_ (.A(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__and3b_2 _15231_ (.A_N(_04627_),
    .B(_06207_),
    .C(_04626_),
    .X(_08306_));
 sky130_fd_sc_hd__clkbuf_8 _15232_ (.A(_08306_),
    .X(_08307_));
 sky130_fd_sc_hd__a21o_1 _15233_ (.A1(net4310),
    .A2(_08305_),
    .B1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__a21oi_2 _15234_ (.A1(_08299_),
    .A2(_08302_),
    .B1(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__buf_2 _15235_ (.A(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__buf_4 _15236_ (.A(_08306_),
    .X(_08311_));
 sky130_fd_sc_hd__buf_6 _15237_ (.A(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__clkbuf_4 _15238_ (.A(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__clkbuf_8 _15239_ (.A(_08299_),
    .X(_08314_));
 sky130_fd_sc_hd__nand2_2 _15240_ (.A(net7552),
    .B(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__or2_1 _15241_ (.A(_08313_),
    .B(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__clkbuf_4 _15242_ (.A(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__or2_2 _15243_ (.A(_08310_),
    .B(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__or2_2 _15244_ (.A(net3507),
    .B(_04818_),
    .X(_08319_));
 sky130_fd_sc_hd__buf_4 _15245_ (.A(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__mux2_1 _15246_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(_08300_),
    .X(_08321_));
 sky130_fd_sc_hd__nor2_1 _15247_ (.A(_08320_),
    .B(net7589),
    .Y(_08322_));
 sky130_fd_sc_hd__a31o_1 _15248_ (.A1(_06625_),
    .A2(_08024_),
    .A3(_08320_),
    .B1(net7590),
    .X(_08323_));
 sky130_fd_sc_hd__nor2_1 _15249_ (.A(net4315),
    .B(_08299_),
    .Y(_08324_));
 sky130_fd_sc_hd__a211o_2 _15250_ (.A1(_08299_),
    .A2(_08323_),
    .B1(_08324_),
    .C1(_08312_),
    .X(_08325_));
 sky130_fd_sc_hd__clkbuf_4 _15251_ (.A(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__buf_4 _15252_ (.A(_08307_),
    .X(_08327_));
 sky130_fd_sc_hd__buf_4 _15253_ (.A(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__nand2_2 _15254_ (.A(net7476),
    .B(_08314_),
    .Y(_08329_));
 sky130_fd_sc_hd__or2_1 _15255_ (.A(_08328_),
    .B(net7477),
    .X(_08330_));
 sky130_fd_sc_hd__clkbuf_4 _15256_ (.A(_08330_),
    .X(_08331_));
 sky130_fd_sc_hd__or3_2 _15257_ (.A(_08318_),
    .B(_08326_),
    .C(_08331_),
    .X(_08332_));
 sky130_fd_sc_hd__xor2_1 _15258_ (.A(net3024),
    .B(net4355),
    .X(_08333_));
 sky130_fd_sc_hd__mux2_1 _15259_ (.A0(_08333_),
    .A1(net3024),
    .S(_06177_),
    .X(_08334_));
 sky130_fd_sc_hd__mux2_1 _15260_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_08334_),
    .S(_08303_),
    .X(_08335_));
 sky130_fd_sc_hd__and2_1 _15261_ (.A(_06523_),
    .B(_06524_),
    .X(_08336_));
 sky130_fd_sc_hd__or4_1 _15262_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .C(_06427_),
    .D(_06418_),
    .X(_08337_));
 sky130_fd_sc_hd__or4_1 _15263_ (.A(_06510_),
    .B(_06507_),
    .C(_06497_),
    .D(net7401),
    .X(_08338_));
 sky130_fd_sc_hd__and4b_1 _15264_ (.A_N(net7402),
    .B(_06492_),
    .C(_06500_),
    .D(_06482_),
    .X(_08339_));
 sky130_fd_sc_hd__nor2_1 _15265_ (.A(_06470_),
    .B(_06489_),
    .Y(_08340_));
 sky130_fd_sc_hd__a41o_2 _15266_ (.A1(_06535_),
    .A2(_08336_),
    .A3(net7403),
    .A4(_08340_),
    .B1(_06570_),
    .X(_08341_));
 sky130_fd_sc_hd__nor2_1 _15267_ (.A(net4306),
    .B(net4335),
    .Y(_08342_));
 sky130_fd_sc_hd__and2_1 _15268_ (.A(net4306),
    .B(net4335),
    .X(_08343_));
 sky130_fd_sc_hd__or3_1 _15269_ (.A(_08341_),
    .B(_08342_),
    .C(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__a21oi_1 _15270_ (.A1(net4306),
    .A2(_08341_),
    .B1(_06209_),
    .Y(_08345_));
 sky130_fd_sc_hd__a2bb2o_2 _15271_ (.A1_N(_08311_),
    .A2_N(net7761),
    .B1(_08344_),
    .B2(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__buf_2 _15272_ (.A(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__nor2_1 _15273_ (.A(net4086),
    .B(_06152_),
    .Y(_08348_));
 sky130_fd_sc_hd__a211o_1 _15274_ (.A1(_08300_),
    .A2(_06492_),
    .B1(_08319_),
    .C1(net7510),
    .X(_08349_));
 sky130_fd_sc_hd__a21o_1 _15275_ (.A1(_08119_),
    .A2(_08124_),
    .B1(_08294_),
    .X(_08350_));
 sky130_fd_sc_hd__a21o_4 _15276_ (.A1(net7511),
    .A2(_08350_),
    .B1(_08304_),
    .X(_08351_));
 sky130_fd_sc_hd__a21oi_4 _15277_ (.A1(net3392),
    .A2(_08305_),
    .B1(_08307_),
    .Y(_08352_));
 sky130_fd_sc_hd__a2bb2o_4 _15278_ (.A1_N(net3397),
    .A2_N(_06209_),
    .B1(_08351_),
    .B2(_08352_),
    .X(_08353_));
 sky130_fd_sc_hd__or3_1 _15279_ (.A(net4893),
    .B(net3024),
    .C(net4355),
    .X(_08354_));
 sky130_fd_sc_hd__o21ai_1 _15280_ (.A1(net3024),
    .A2(net4355),
    .B1(net4893),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_1 _15281_ (.A(_08354_),
    .B(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__inv_2 _15282_ (.A(net2940),
    .Y(_08357_));
 sky130_fd_sc_hd__mux2_1 _15283_ (.A0(_08356_),
    .A1(_08357_),
    .S(_06177_),
    .X(_08358_));
 sky130_fd_sc_hd__or2_1 _15284_ (.A(_08297_),
    .B(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__a21oi_1 _15285_ (.A1(net3206),
    .A2(_08297_),
    .B1(_08307_),
    .Y(_08360_));
 sky130_fd_sc_hd__inv_2 _15286_ (.A(net5463),
    .Y(_08361_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(_08361_),
    .B(_08342_),
    .Y(_08362_));
 sky130_fd_sc_hd__or2_1 _15288_ (.A(_08361_),
    .B(_08342_),
    .X(_08363_));
 sky130_fd_sc_hd__nand2_1 _15289_ (.A(_08362_),
    .B(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__mux2_1 _15290_ (.A0(_08364_),
    .A1(_08361_),
    .S(_08341_),
    .X(_08365_));
 sky130_fd_sc_hd__a22o_2 _15291_ (.A1(_08359_),
    .A2(net7779),
    .B1(_08365_),
    .B2(_08311_),
    .X(_08366_));
 sky130_fd_sc_hd__buf_2 _15292_ (.A(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__inv_2 _15293_ (.A(_06171_),
    .Y(_08368_));
 sky130_fd_sc_hd__mux2_1 _15294_ (.A0(net7809),
    .A1(_06497_),
    .S(net4086),
    .X(_08369_));
 sky130_fd_sc_hd__mux2_1 _15295_ (.A0(_08117_),
    .A1(net7810),
    .S(_08294_),
    .X(_08370_));
 sky130_fd_sc_hd__a21o_1 _15296_ (.A1(net3057),
    .A2(_08303_),
    .B1(_08306_),
    .X(_08371_));
 sky130_fd_sc_hd__a21oi_4 _15297_ (.A1(_08298_),
    .A2(_08370_),
    .B1(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__o21bai_4 _15298_ (.A1(net3172),
    .A2(_06209_),
    .B1_N(_08372_),
    .Y(_08373_));
 sky130_fd_sc_hd__o22ai_1 _15299_ (.A1(_08347_),
    .A2(_08353_),
    .B1(_08367_),
    .B2(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__or2_1 _15300_ (.A(net2942),
    .B(_08354_),
    .X(_08375_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(net2942),
    .B(_08354_),
    .Y(_08376_));
 sky130_fd_sc_hd__and2_1 _15302_ (.A(_08375_),
    .B(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__mux2_1 _15303_ (.A0(_08377_),
    .A1(net2942),
    .S(_06178_),
    .X(_08378_));
 sky130_fd_sc_hd__buf_4 _15304_ (.A(_08304_),
    .X(_08379_));
 sky130_fd_sc_hd__mux2_1 _15305_ (.A0(net3356),
    .A1(_08378_),
    .S(_08379_),
    .X(_08380_));
 sky130_fd_sc_hd__buf_4 _15306_ (.A(net7404),
    .X(_08381_));
 sky130_fd_sc_hd__nand2_1 _15307_ (.A(net4338),
    .B(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__or2_1 _15308_ (.A(net4338),
    .B(_08362_),
    .X(_08383_));
 sky130_fd_sc_hd__nand2_1 _15309_ (.A(net4338),
    .B(_08362_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand2_1 _15310_ (.A(_08383_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__o21a_1 _15311_ (.A1(_08381_),
    .A2(_08385_),
    .B1(_08327_),
    .X(_08386_));
 sky130_fd_sc_hd__a2bb2o_4 _15312_ (.A1_N(_08312_),
    .A2_N(_08380_),
    .B1(_08382_),
    .B2(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__nor2_1 _15313_ (.A(_08300_),
    .B(_06162_),
    .Y(_08388_));
 sky130_fd_sc_hd__a211o_1 _15314_ (.A1(_08300_),
    .A2(_06500_),
    .B1(_08320_),
    .C1(_08388_),
    .X(_08389_));
 sky130_fd_sc_hd__a21o_1 _15315_ (.A1(_08100_),
    .A2(_08105_),
    .B1(_08294_),
    .X(_08390_));
 sky130_fd_sc_hd__a21o_2 _15316_ (.A1(net7777),
    .A2(_08390_),
    .B1(_08304_),
    .X(_08391_));
 sky130_fd_sc_hd__a21oi_1 _15317_ (.A1(net3315),
    .A2(_08305_),
    .B1(_08311_),
    .Y(_08392_));
 sky130_fd_sc_hd__a2bb2o_2 _15318_ (.A1_N(net3149),
    .A2_N(_06210_),
    .B1(_08391_),
    .B2(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__buf_2 _15319_ (.A(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__nor2_1 _15320_ (.A(_08387_),
    .B(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__or4_1 _15321_ (.A(_08346_),
    .B(_08353_),
    .C(_08366_),
    .D(_08373_),
    .X(_08396_));
 sky130_fd_sc_hd__a21bo_1 _15322_ (.A1(_08374_),
    .A2(_08395_),
    .B1_N(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__xor2_1 _15323_ (.A(net4294),
    .B(_08375_),
    .X(_08398_));
 sky130_fd_sc_hd__mux2_1 _15324_ (.A0(_08398_),
    .A1(net4294),
    .S(_06177_),
    .X(_08399_));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(net3262),
    .A1(_08399_),
    .S(_08303_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_1 _15326_ (.A(net2935),
    .B(_08341_),
    .Y(_08401_));
 sky130_fd_sc_hd__xnor2_1 _15327_ (.A(net2935),
    .B(_08383_),
    .Y(_08402_));
 sky130_fd_sc_hd__o21a_1 _15328_ (.A1(_08341_),
    .A2(_08402_),
    .B1(_08307_),
    .X(_08403_));
 sky130_fd_sc_hd__a2bb2o_2 _15329_ (.A1_N(_08307_),
    .A2_N(_08400_),
    .B1(_08401_),
    .B2(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__buf_2 _15330_ (.A(_08404_),
    .X(_08405_));
 sky130_fd_sc_hd__mux2_1 _15331_ (.A0(_06156_),
    .A1(_06507_),
    .S(net4086),
    .X(_08406_));
 sky130_fd_sc_hd__mux2_1 _15332_ (.A0(_08096_),
    .A1(net7775),
    .S(_08294_),
    .X(_08407_));
 sky130_fd_sc_hd__a21o_1 _15333_ (.A1(net3115),
    .A2(_08304_),
    .B1(_08306_),
    .X(_08408_));
 sky130_fd_sc_hd__a21oi_4 _15334_ (.A1(_08298_),
    .A2(_08407_),
    .B1(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__o21bai_4 _15335_ (.A1(net3216),
    .A2(_06210_),
    .B1_N(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__clkbuf_4 _15336_ (.A(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__or3_1 _15337_ (.A(net3003),
    .B(net4294),
    .C(_08375_),
    .X(_08412_));
 sky130_fd_sc_hd__o21ai_1 _15338_ (.A1(net4294),
    .A2(_08375_),
    .B1(net3003),
    .Y(_08413_));
 sky130_fd_sc_hd__and2_1 _15339_ (.A(_08412_),
    .B(_08413_),
    .X(_08414_));
 sky130_fd_sc_hd__mux2_1 _15340_ (.A0(_08414_),
    .A1(net3003),
    .S(_06177_),
    .X(_08415_));
 sky130_fd_sc_hd__mux2_1 _15341_ (.A0(net645),
    .A1(_08415_),
    .S(_08303_),
    .X(_08416_));
 sky130_fd_sc_hd__nand2_1 _15342_ (.A(net4300),
    .B(net7404),
    .Y(_08417_));
 sky130_fd_sc_hd__or3_1 _15343_ (.A(net4300),
    .B(net2935),
    .C(_08383_),
    .X(_08418_));
 sky130_fd_sc_hd__o21ai_1 _15344_ (.A1(net2935),
    .A2(_08383_),
    .B1(net4300),
    .Y(_08419_));
 sky130_fd_sc_hd__nand2_1 _15345_ (.A(_08418_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__o21a_1 _15346_ (.A1(net7404),
    .A2(_08420_),
    .B1(_08306_),
    .X(_08421_));
 sky130_fd_sc_hd__a2bb2o_4 _15347_ (.A1_N(_08307_),
    .A2_N(_08416_),
    .B1(_08417_),
    .B2(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__or4_1 _15348_ (.A(_08393_),
    .B(_08405_),
    .C(_08411_),
    .D(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__clkbuf_4 _15349_ (.A(_08422_),
    .X(_08424_));
 sky130_fd_sc_hd__o22ai_1 _15350_ (.A1(_08394_),
    .A2(_08405_),
    .B1(_08411_),
    .B2(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand2_1 _15351_ (.A(_08423_),
    .B(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__mux2_1 _15352_ (.A0(_06163_),
    .A1(_06510_),
    .S(_08300_),
    .X(_08427_));
 sky130_fd_sc_hd__nand2_1 _15353_ (.A(_08295_),
    .B(net7766),
    .Y(_08428_));
 sky130_fd_sc_hd__a21o_1 _15354_ (.A1(_08080_),
    .A2(_08085_),
    .B1(_08295_),
    .X(_08429_));
 sky130_fd_sc_hd__a21o_2 _15355_ (.A1(_08428_),
    .A2(_08429_),
    .B1(_08305_),
    .X(_08430_));
 sky130_fd_sc_hd__a21oi_2 _15356_ (.A1(net4382),
    .A2(_08379_),
    .B1(_08311_),
    .Y(_08431_));
 sky130_fd_sc_hd__a2bb2o_2 _15357_ (.A1_N(net3102),
    .A2_N(_06210_),
    .B1(_08430_),
    .B2(_08431_),
    .X(_08432_));
 sky130_fd_sc_hd__clkbuf_4 _15358_ (.A(_08432_),
    .X(_08433_));
 sky130_fd_sc_hd__or2_1 _15359_ (.A(net4063),
    .B(_08412_),
    .X(_08434_));
 sky130_fd_sc_hd__nand2_1 _15360_ (.A(net4063),
    .B(_08412_),
    .Y(_08435_));
 sky130_fd_sc_hd__and2_1 _15361_ (.A(_08434_),
    .B(_08435_),
    .X(_08436_));
 sky130_fd_sc_hd__mux2_1 _15362_ (.A0(_08436_),
    .A1(net4063),
    .S(_06178_),
    .X(_08437_));
 sky130_fd_sc_hd__mux2_1 _15363_ (.A0(net6253),
    .A1(_08437_),
    .S(_08305_),
    .X(_08438_));
 sky130_fd_sc_hd__or2_1 _15364_ (.A(net3008),
    .B(_08418_),
    .X(_08439_));
 sky130_fd_sc_hd__nand2_1 _15365_ (.A(net3008),
    .B(_08418_),
    .Y(_08440_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_08439_),
    .B(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__nor2_1 _15367_ (.A(_08381_),
    .B(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a211o_1 _15368_ (.A1(net3008),
    .A2(_08381_),
    .B1(_08442_),
    .C1(_06209_),
    .X(_08443_));
 sky130_fd_sc_hd__o21ai_4 _15369_ (.A1(_08312_),
    .A2(_08438_),
    .B1(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__nor2_1 _15370_ (.A(_08433_),
    .B(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__xnor2_2 _15371_ (.A(_08426_),
    .B(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__xnor2_2 _15372_ (.A(_08397_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__or4_1 _15373_ (.A(_08405_),
    .B(_08411_),
    .C(_08422_),
    .D(_08432_),
    .X(_08448_));
 sky130_fd_sc_hd__clkbuf_4 _15374_ (.A(_08405_),
    .X(_08449_));
 sky130_fd_sc_hd__o22ai_2 _15375_ (.A1(_08449_),
    .A2(_08411_),
    .B1(_08424_),
    .B2(_08433_),
    .Y(_08450_));
 sky130_fd_sc_hd__mux2_1 _15376_ (.A0(_06165_),
    .A1(_06418_),
    .S(net4086),
    .X(_08451_));
 sky130_fd_sc_hd__mux2_1 _15377_ (.A0(_08074_),
    .A1(net7773),
    .S(_08295_),
    .X(_08452_));
 sky130_fd_sc_hd__a21o_1 _15378_ (.A1(net3193),
    .A2(_08304_),
    .B1(_08307_),
    .X(_08453_));
 sky130_fd_sc_hd__a21oi_4 _15379_ (.A1(_08298_),
    .A2(_08452_),
    .B1(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__o21bai_4 _15380_ (.A1(net3332),
    .A2(_06210_),
    .B1_N(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__clkbuf_4 _15381_ (.A(_08455_),
    .X(_08456_));
 sky130_fd_sc_hd__nor2_1 _15382_ (.A(_08444_),
    .B(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__nand3_1 _15383_ (.A(_08448_),
    .B(_08450_),
    .C(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__nand2_1 _15384_ (.A(_08448_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__and2b_1 _15385_ (.A_N(_08447_),
    .B(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__a21o_1 _15386_ (.A1(_08397_),
    .A2(_08446_),
    .B1(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__nor2_2 _15387_ (.A(_08325_),
    .B(_08331_),
    .Y(_08462_));
 sky130_fd_sc_hd__xnor2_4 _15388_ (.A(_08318_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__xor2_1 _15389_ (.A(net4358),
    .B(_08434_),
    .X(_08464_));
 sky130_fd_sc_hd__mux2_1 _15390_ (.A0(_08464_),
    .A1(net4358),
    .S(_06178_),
    .X(_08465_));
 sky130_fd_sc_hd__mux2_1 _15391_ (.A0(net695),
    .A1(_08465_),
    .S(_08305_),
    .X(_08466_));
 sky130_fd_sc_hd__xnor2_1 _15392_ (.A(net3028),
    .B(_08439_),
    .Y(_08467_));
 sky130_fd_sc_hd__nor2_1 _15393_ (.A(_08381_),
    .B(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__a211o_1 _15394_ (.A1(net3028),
    .A2(_08381_),
    .B1(_08468_),
    .C1(_06209_),
    .X(_08469_));
 sky130_fd_sc_hd__o21ai_4 _15395_ (.A1(_08312_),
    .A2(_08466_),
    .B1(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__buf_2 _15396_ (.A(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__nor2_1 _15397_ (.A(_08433_),
    .B(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__or3_4 _15398_ (.A(net4288),
    .B(net4358),
    .C(_08434_),
    .X(_08473_));
 sky130_fd_sc_hd__o21ai_1 _15399_ (.A1(net4358),
    .A2(_08434_),
    .B1(net4288),
    .Y(_08474_));
 sky130_fd_sc_hd__and2_1 _15400_ (.A(_08473_),
    .B(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__mux2_1 _15401_ (.A0(_08475_),
    .A1(net4288),
    .S(_06178_),
    .X(_08476_));
 sky130_fd_sc_hd__nand2_1 _15402_ (.A(_08379_),
    .B(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__a21oi_1 _15403_ (.A1(net7939),
    .A2(_08298_),
    .B1(_08327_),
    .Y(_08478_));
 sky130_fd_sc_hd__or3_4 _15404_ (.A(net4105),
    .B(net3028),
    .C(_08439_),
    .X(_08479_));
 sky130_fd_sc_hd__o21ai_1 _15405_ (.A1(net3028),
    .A2(_08439_),
    .B1(net4105),
    .Y(_08480_));
 sky130_fd_sc_hd__nand2_1 _15406_ (.A(_08479_),
    .B(_08480_),
    .Y(_08481_));
 sky130_fd_sc_hd__mux2_1 _15407_ (.A0(_08481_),
    .A1(_04846_),
    .S(_08381_),
    .X(_08482_));
 sky130_fd_sc_hd__a22o_2 _15408_ (.A1(_08477_),
    .A2(_08478_),
    .B1(_08482_),
    .B2(_08327_),
    .X(_08483_));
 sky130_fd_sc_hd__buf_2 _15409_ (.A(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__nor2_1 _15410_ (.A(_08456_),
    .B(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__xnor2_1 _15411_ (.A(_08472_),
    .B(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__mux2_1 _15412_ (.A0(_06166_),
    .A1(_06427_),
    .S(net4086),
    .X(_08487_));
 sky130_fd_sc_hd__mux2_1 _15413_ (.A0(_08059_),
    .A1(net7764),
    .S(_08295_),
    .X(_08488_));
 sky130_fd_sc_hd__a21o_1 _15414_ (.A1(net3217),
    .A2(_08304_),
    .B1(_08307_),
    .X(_08489_));
 sky130_fd_sc_hd__a21o_4 _15415_ (.A1(_08299_),
    .A2(_08488_),
    .B1(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__or2_1 _15416_ (.A(net3470),
    .B(_06209_),
    .X(_08491_));
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(_08490_),
    .B(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__clkbuf_4 _15418_ (.A(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__nand2_1 _15419_ (.A(net6259),
    .B(_08299_),
    .Y(_08494_));
 sky130_fd_sc_hd__o31a_1 _15420_ (.A1(_06178_),
    .A2(_08314_),
    .A3(_08473_),
    .B1(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__or3_1 _15421_ (.A(_06210_),
    .B(_08381_),
    .C(_08479_),
    .X(_08496_));
 sky130_fd_sc_hd__o21a_2 _15422_ (.A1(_08328_),
    .A2(_08495_),
    .B1(_08496_),
    .X(_08497_));
 sky130_fd_sc_hd__buf_2 _15423_ (.A(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__or2_1 _15424_ (.A(_08493_),
    .B(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__xnor2_1 _15425_ (.A(_08486_),
    .B(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__o21bai_4 _15426_ (.A1(net3492),
    .A2(_06210_),
    .B1_N(_08309_),
    .Y(_08501_));
 sky130_fd_sc_hd__or2_1 _15427_ (.A(_08497_),
    .B(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__or4_1 _15428_ (.A(_08455_),
    .B(_08470_),
    .C(_08483_),
    .D(_08493_),
    .X(_08503_));
 sky130_fd_sc_hd__o22ai_1 _15429_ (.A1(_08456_),
    .A2(_08470_),
    .B1(_08484_),
    .B2(_08493_),
    .Y(_08504_));
 sky130_fd_sc_hd__nand2_1 _15430_ (.A(_08503_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21a_1 _15431_ (.A1(_08502_),
    .A2(_08505_),
    .B1(_08503_),
    .X(_08506_));
 sky130_fd_sc_hd__nor2_1 _15432_ (.A(_08500_),
    .B(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__nand2_1 _15433_ (.A(_08500_),
    .B(_08506_),
    .Y(_08508_));
 sky130_fd_sc_hd__and2b_1 _15434_ (.A_N(_08507_),
    .B(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__xor2_2 _15435_ (.A(_08463_),
    .B(_08509_),
    .X(_08510_));
 sky130_fd_sc_hd__xnor2_2 _15436_ (.A(_08461_),
    .B(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__nor2_1 _15437_ (.A(_08317_),
    .B(_08326_),
    .Y(_08512_));
 sky130_fd_sc_hd__xnor2_1 _15438_ (.A(_08502_),
    .B(_08505_),
    .Y(_08513_));
 sky130_fd_sc_hd__a21boi_4 _15439_ (.A1(net3471),
    .A2(_08328_),
    .B1_N(_08325_),
    .Y(_08514_));
 sky130_fd_sc_hd__or2_1 _15440_ (.A(_08497_),
    .B(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__clkbuf_4 _15441_ (.A(_08484_),
    .X(_08516_));
 sky130_fd_sc_hd__clkbuf_4 _15442_ (.A(_08501_),
    .X(_08517_));
 sky130_fd_sc_hd__or2_1 _15443_ (.A(_08470_),
    .B(_08492_),
    .X(_08518_));
 sky130_fd_sc_hd__o21a_1 _15444_ (.A1(_08516_),
    .A2(_08517_),
    .B1(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__or3_1 _15445_ (.A(_08516_),
    .B(_08501_),
    .C(_08518_),
    .X(_08520_));
 sky130_fd_sc_hd__o21a_1 _15446_ (.A1(_08515_),
    .A2(_08519_),
    .B1(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__xor2_1 _15447_ (.A(_08513_),
    .B(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__nor2_1 _15448_ (.A(_08513_),
    .B(_08521_),
    .Y(_08523_));
 sky130_fd_sc_hd__a21o_1 _15449_ (.A1(_08512_),
    .A2(_08522_),
    .B1(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__or2b_1 _15450_ (.A(_08511_),
    .B_N(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__a21boi_1 _15451_ (.A1(_08461_),
    .A2(_08510_),
    .B1_N(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__or2_1 _15452_ (.A(_08332_),
    .B(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__inv_2 _15453_ (.A(_08527_),
    .Y(_08528_));
 sky130_fd_sc_hd__clkbuf_4 _15454_ (.A(_08373_),
    .X(_08529_));
 sky130_fd_sc_hd__o22ai_2 _15455_ (.A1(_08353_),
    .A2(_08405_),
    .B1(_08424_),
    .B2(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__nor2_1 _15456_ (.A(_08394_),
    .B(_08444_),
    .Y(_08531_));
 sky130_fd_sc_hd__or4_1 _15457_ (.A(_08353_),
    .B(_08373_),
    .C(_08405_),
    .D(_08422_),
    .X(_08532_));
 sky130_fd_sc_hd__a21bo_1 _15458_ (.A1(_08530_),
    .A2(_08531_),
    .B1_N(_08532_),
    .X(_08533_));
 sky130_fd_sc_hd__o21ai_1 _15459_ (.A1(_08130_),
    .A2(_08137_),
    .B1(_08144_),
    .Y(_08534_));
 sky130_fd_sc_hd__or3_1 _15460_ (.A(_08130_),
    .B(_08137_),
    .C(_08144_),
    .X(_08535_));
 sky130_fd_sc_hd__a21o_1 _15461_ (.A1(_08534_),
    .A2(_08535_),
    .B1(_08295_),
    .X(_08536_));
 sky130_fd_sc_hd__nand2_1 _15462_ (.A(_08300_),
    .B(_06470_),
    .Y(_08537_));
 sky130_fd_sc_hd__o211a_1 _15463_ (.A1(_04646_),
    .A2(_06174_),
    .B1(_08294_),
    .C1(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__nor2_1 _15464_ (.A(_08304_),
    .B(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__a22o_4 _15465_ (.A1(net3210),
    .A2(_08305_),
    .B1(_08536_),
    .B2(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__nand2_1 _15466_ (.A(net3041),
    .B(_08327_),
    .Y(_08541_));
 sky130_fd_sc_hd__a21boi_2 _15467_ (.A1(_06210_),
    .A2(_08540_),
    .B1_N(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__xor2_1 _15468_ (.A(_08130_),
    .B(_08137_),
    .X(_08543_));
 sky130_fd_sc_hd__nor2_1 _15469_ (.A(_08300_),
    .B(net8016),
    .Y(_08544_));
 sky130_fd_sc_hd__a211o_1 _15470_ (.A1(_08300_),
    .A2(_06482_),
    .B1(_08320_),
    .C1(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__o21a_4 _15471_ (.A1(_08295_),
    .A2(_08543_),
    .B1(_08545_),
    .X(_08546_));
 sky130_fd_sc_hd__o21ai_2 _15472_ (.A1(net3161),
    .A2(_08298_),
    .B1(_06209_),
    .Y(_08547_));
 sky130_fd_sc_hd__a21o_4 _15473_ (.A1(_08299_),
    .A2(_08546_),
    .B1(_08547_),
    .X(_08548_));
 sky130_fd_sc_hd__nand2_1 _15474_ (.A(net3065),
    .B(_08327_),
    .Y(_08549_));
 sky130_fd_sc_hd__and2_2 _15475_ (.A(_08548_),
    .B(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__or4_2 _15476_ (.A(_08347_),
    .B(_08367_),
    .C(_08542_),
    .D(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__nand2_1 _15477_ (.A(_08300_),
    .B(_06489_),
    .Y(_08552_));
 sky130_fd_sc_hd__o21a_1 _15478_ (.A1(net4086),
    .A2(_06151_),
    .B1(_08294_),
    .X(_08553_));
 sky130_fd_sc_hd__a22o_1 _15479_ (.A1(_08130_),
    .A2(_08320_),
    .B1(_08552_),
    .B2(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__nor2_1 _15480_ (.A(net3148),
    .B(_08297_),
    .Y(_08555_));
 sky130_fd_sc_hd__a211o_4 _15481_ (.A1(_08298_),
    .A2(_08554_),
    .B1(_08555_),
    .C1(_08307_),
    .X(_08556_));
 sky130_fd_sc_hd__a21boi_4 _15482_ (.A1(net3171),
    .A2(_08312_),
    .B1_N(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__or2_1 _15483_ (.A(_08387_),
    .B(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__clkbuf_4 _15484_ (.A(_08347_),
    .X(_08559_));
 sky130_fd_sc_hd__clkbuf_4 _15485_ (.A(_08367_),
    .X(_08560_));
 sky130_fd_sc_hd__o22ai_1 _15486_ (.A1(_08559_),
    .A2(_08542_),
    .B1(_08550_),
    .B2(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__nand3b_1 _15487_ (.A_N(_08558_),
    .B(_08561_),
    .C(_08551_),
    .Y(_08562_));
 sky130_fd_sc_hd__or4_1 _15488_ (.A(_08353_),
    .B(_08405_),
    .C(_08424_),
    .D(_08557_),
    .X(_08563_));
 sky130_fd_sc_hd__clkbuf_4 _15489_ (.A(_08353_),
    .X(_08564_));
 sky130_fd_sc_hd__clkbuf_4 _15490_ (.A(_08557_),
    .X(_08565_));
 sky130_fd_sc_hd__o22ai_2 _15491_ (.A1(_08564_),
    .A2(_08424_),
    .B1(_08565_),
    .B2(_08449_),
    .Y(_08566_));
 sky130_fd_sc_hd__nand2_1 _15492_ (.A(_08563_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__nor2_1 _15493_ (.A(_08529_),
    .B(_08444_),
    .Y(_08568_));
 sky130_fd_sc_hd__xor2_1 _15494_ (.A(_08567_),
    .B(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__a21o_1 _15495_ (.A1(_08551_),
    .A2(_08562_),
    .B1(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__nand3_1 _15496_ (.A(_08551_),
    .B(_08562_),
    .C(_08569_),
    .Y(_08571_));
 sky130_fd_sc_hd__nand2_1 _15497_ (.A(_08570_),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__xnor2_2 _15498_ (.A(_08533_),
    .B(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__clkbuf_4 _15499_ (.A(_08542_),
    .X(_08574_));
 sky130_fd_sc_hd__o21a_4 _15500_ (.A1(_08130_),
    .A2(_08137_),
    .B1(_08144_),
    .X(_08575_));
 sky130_fd_sc_hd__xnor2_2 _15501_ (.A(_08152_),
    .B(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_1 _15502_ (.A(_04646_),
    .B(_08336_),
    .Y(_08577_));
 sky130_fd_sc_hd__o211a_2 _15503_ (.A1(_04646_),
    .A2(net8126),
    .B1(_08295_),
    .C1(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__a211o_2 _15504_ (.A1(_08320_),
    .A2(_08576_),
    .B1(_08578_),
    .C1(_08305_),
    .X(_08579_));
 sky130_fd_sc_hd__o21a_1 _15505_ (.A1(net3114),
    .A2(_08299_),
    .B1(_06210_),
    .X(_08580_));
 sky130_fd_sc_hd__a22oi_4 _15506_ (.A1(net3162),
    .A2(_08328_),
    .B1(_08579_),
    .B2(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__clkbuf_4 _15507_ (.A(_08581_),
    .X(_08582_));
 sky130_fd_sc_hd__or4_1 _15508_ (.A(_08559_),
    .B(_08560_),
    .C(_08574_),
    .D(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__clkbuf_4 _15509_ (.A(_08559_),
    .X(_08584_));
 sky130_fd_sc_hd__o22ai_2 _15510_ (.A1(_08560_),
    .A2(_08574_),
    .B1(_08582_),
    .B2(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__nand2_1 _15511_ (.A(_08583_),
    .B(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__clkbuf_4 _15512_ (.A(_08387_),
    .X(_08587_));
 sky130_fd_sc_hd__clkbuf_4 _15513_ (.A(_08550_),
    .X(_08588_));
 sky130_fd_sc_hd__nor2_1 _15514_ (.A(_08587_),
    .B(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__xnor2_2 _15515_ (.A(_08586_),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__inv_2 _15516_ (.A(_08155_),
    .Y(_08591_));
 sky130_fd_sc_hd__nor2_1 _15517_ (.A(_08152_),
    .B(_08575_),
    .Y(_08592_));
 sky130_fd_sc_hd__xnor2_2 _15518_ (.A(_08591_),
    .B(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_1 _15519_ (.A(_04646_),
    .B(_06535_),
    .Y(_08594_));
 sky130_fd_sc_hd__o211a_2 _15520_ (.A1(_04646_),
    .A2(_06138_),
    .B1(_08295_),
    .C1(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__a211o_4 _15521_ (.A1(_08320_),
    .A2(_08593_),
    .B1(_08595_),
    .C1(_08379_),
    .X(_08596_));
 sky130_fd_sc_hd__o21a_2 _15522_ (.A1(net3169),
    .A2(_08298_),
    .B1(_06209_),
    .X(_08597_));
 sky130_fd_sc_hd__and2_1 _15523_ (.A(net3046),
    .B(_08312_),
    .X(_08598_));
 sky130_fd_sc_hd__a21o_1 _15524_ (.A1(_08596_),
    .A2(_08597_),
    .B1(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__mux2_1 _15525_ (.A0(net4355),
    .A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .S(_08297_),
    .X(_08600_));
 sky130_fd_sc_hd__or2_1 _15526_ (.A(_08311_),
    .B(net7769),
    .X(_08601_));
 sky130_fd_sc_hd__o21a_1 _15527_ (.A1(net4335),
    .A2(_06211_),
    .B1(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__nand2_1 _15528_ (.A(_08599_),
    .B(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__a21oi_1 _15529_ (.A1(_08068_),
    .A2(_08149_),
    .B1(_08151_),
    .Y(_08604_));
 sky130_fd_sc_hd__a211oi_1 _15530_ (.A1(_08150_),
    .A2(_08104_),
    .B1(_08159_),
    .C1(_08047_),
    .Y(_08605_));
 sky130_fd_sc_hd__a31o_1 _15531_ (.A1(_08604_),
    .A2(_08591_),
    .A3(_08534_),
    .B1(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__or4_4 _15532_ (.A(_08152_),
    .B(_08155_),
    .C(_08160_),
    .D(_08575_),
    .X(_08607_));
 sky130_fd_sc_hd__mux2_1 _15533_ (.A0(_06133_),
    .A1(_06570_),
    .S(net4086),
    .X(_08608_));
 sky130_fd_sc_hd__o21a_4 _15534_ (.A1(_08319_),
    .A2(_08608_),
    .B1(_08297_),
    .X(_08609_));
 sky130_fd_sc_hd__inv_2 _15535_ (.A(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__a31o_4 _15536_ (.A1(_08320_),
    .A2(_08606_),
    .A3(_08607_),
    .B1(_08610_),
    .X(_08611_));
 sky130_fd_sc_hd__or4_4 _15537_ (.A(net3539),
    .B(_08327_),
    .C(_08379_),
    .D(_08611_),
    .X(_08612_));
 sky130_fd_sc_hd__nor2_2 _15538_ (.A(net3722),
    .B(_08304_),
    .Y(_08613_));
 sky130_fd_sc_hd__and4_1 _15539_ (.A(_08604_),
    .B(_08591_),
    .C(_08605_),
    .D(_08534_),
    .X(_08614_));
 sky130_fd_sc_hd__nand2_2 _15540_ (.A(_08166_),
    .B(_08167_),
    .Y(_08615_));
 sky130_fd_sc_hd__o41a_1 _15541_ (.A1(_08152_),
    .A2(_08155_),
    .A3(_08160_),
    .A4(_08575_),
    .B1(_08615_),
    .X(_08616_));
 sky130_fd_sc_hd__a311o_1 _15542_ (.A1(_08166_),
    .A2(_08167_),
    .A3(_08614_),
    .B1(_08616_),
    .C1(_08296_),
    .X(_08617_));
 sky130_fd_sc_hd__a22o_4 _15543_ (.A1(net3063),
    .A2(_08379_),
    .B1(_08609_),
    .B2(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__and3_1 _15544_ (.A(_06211_),
    .B(_08613_),
    .C(_08618_),
    .X(_08619_));
 sky130_fd_sc_hd__xor2_2 _15545_ (.A(_08612_),
    .B(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__xor2_2 _15546_ (.A(_08603_),
    .B(_08620_),
    .X(_08621_));
 sky130_fd_sc_hd__inv_2 _15547_ (.A(_08597_),
    .Y(_08622_));
 sky130_fd_sc_hd__nand2_1 _15548_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08298_),
    .Y(_08623_));
 sky130_fd_sc_hd__or4b_4 _15549_ (.A(_08622_),
    .B(_08612_),
    .C(net7444),
    .D_N(_08596_),
    .X(_08624_));
 sky130_fd_sc_hd__o21ai_4 _15550_ (.A1(net4335),
    .A2(_06210_),
    .B1(_08601_),
    .Y(_08625_));
 sky130_fd_sc_hd__clkbuf_4 _15551_ (.A(_08625_),
    .X(_08626_));
 sky130_fd_sc_hd__nor2_1 _15552_ (.A(_08581_),
    .B(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__buf_2 _15553_ (.A(_08379_),
    .X(_08628_));
 sky130_fd_sc_hd__nand2_1 _15554_ (.A(net3120),
    .B(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__a21o_1 _15555_ (.A1(_08629_),
    .A2(_08611_),
    .B1(_08312_),
    .X(_08630_));
 sky130_fd_sc_hd__nor2_2 _15556_ (.A(net3539),
    .B(_08304_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand2_4 _15557_ (.A(_06208_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__buf_4 _15558_ (.A(_08320_),
    .X(_08633_));
 sky130_fd_sc_hd__a21oi_4 _15559_ (.A1(_08633_),
    .A2(_08593_),
    .B1(_08595_),
    .Y(_08634_));
 sky130_fd_sc_hd__o22ai_2 _15560_ (.A1(_08630_),
    .A2(net7444),
    .B1(_08632_),
    .B2(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__nand3_2 _15561_ (.A(_08624_),
    .B(_08627_),
    .C(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_1 _15562_ (.A(_08624_),
    .B(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__xor2_2 _15563_ (.A(_08621_),
    .B(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__xnor2_2 _15564_ (.A(_08590_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__a21o_1 _15565_ (.A1(_08624_),
    .A2(_08635_),
    .B1(_08627_),
    .X(_08640_));
 sky130_fd_sc_hd__nand2_2 _15566_ (.A(_06211_),
    .B(_08540_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand2_1 _15567_ (.A(_08641_),
    .B(_08541_),
    .Y(_08642_));
 sky130_fd_sc_hd__a21oi_4 _15568_ (.A1(_08320_),
    .A2(_08576_),
    .B1(_08578_),
    .Y(_08643_));
 sky130_fd_sc_hd__nor2_1 _15569_ (.A(_08643_),
    .B(_08632_),
    .Y(_08644_));
 sky130_fd_sc_hd__a31o_1 _15570_ (.A1(_08596_),
    .A2(_08597_),
    .A3(_08613_),
    .B1(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__and4_1 _15571_ (.A(_08596_),
    .B(_08597_),
    .C(_08613_),
    .D(_08644_),
    .X(_08646_));
 sky130_fd_sc_hd__a31o_1 _15572_ (.A1(_08642_),
    .A2(_08602_),
    .A3(_08645_),
    .B1(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__nand3_1 _15573_ (.A(_08636_),
    .B(_08640_),
    .C(_08647_),
    .Y(_08648_));
 sky130_fd_sc_hd__a21bo_1 _15574_ (.A1(_08551_),
    .A2(_08561_),
    .B1_N(_08558_),
    .X(_08649_));
 sky130_fd_sc_hd__and2_1 _15575_ (.A(_08562_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__a21o_1 _15576_ (.A1(_08636_),
    .A2(_08640_),
    .B1(_08647_),
    .X(_08651_));
 sky130_fd_sc_hd__and3_1 _15577_ (.A(_08648_),
    .B(_08650_),
    .C(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__a31o_1 _15578_ (.A1(_08636_),
    .A2(_08640_),
    .A3(_08647_),
    .B1(_08652_),
    .X(_08653_));
 sky130_fd_sc_hd__xnor2_2 _15579_ (.A(_08639_),
    .B(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__xnor2_2 _15580_ (.A(_08573_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__a21oi_1 _15581_ (.A1(_08648_),
    .A2(_08651_),
    .B1(_08650_),
    .Y(_08656_));
 sky130_fd_sc_hd__or4b_1 _15582_ (.A(_08542_),
    .B(_08626_),
    .C(_08646_),
    .D_N(_08645_),
    .X(_08657_));
 sky130_fd_sc_hd__nand4_1 _15583_ (.A(_08596_),
    .B(_08597_),
    .C(_08613_),
    .D(_08644_),
    .Y(_08658_));
 sky130_fd_sc_hd__a22o_1 _15584_ (.A1(_08642_),
    .A2(_08602_),
    .B1(_08658_),
    .B2(_08645_),
    .X(_08659_));
 sky130_fd_sc_hd__or4b_1 _15585_ (.A(net3722),
    .B(_08327_),
    .C(_08379_),
    .D_N(_08579_),
    .X(_08660_));
 sky130_fd_sc_hd__nand2_1 _15586_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08298_),
    .Y(_08661_));
 sky130_fd_sc_hd__or3b_1 _15587_ (.A(_08327_),
    .B(net4954),
    .C_N(_08540_),
    .X(_08662_));
 sky130_fd_sc_hd__nand2_1 _15588_ (.A(_06209_),
    .B(_08613_),
    .Y(_08663_));
 sky130_fd_sc_hd__clkbuf_4 _15589_ (.A(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__nor2_4 _15590_ (.A(_08311_),
    .B(net4954),
    .Y(_08665_));
 sky130_fd_sc_hd__and4bb_1 _15591_ (.A_N(_08664_),
    .B_N(_08643_),
    .C(_08540_),
    .D(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__a21oi_2 _15592_ (.A1(_08660_),
    .A2(_08662_),
    .B1(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__nor2_1 _15593_ (.A(_08550_),
    .B(_08625_),
    .Y(_08668_));
 sky130_fd_sc_hd__a21o_1 _15594_ (.A1(_08667_),
    .A2(_08668_),
    .B1(_08666_),
    .X(_08669_));
 sky130_fd_sc_hd__a21o_1 _15595_ (.A1(_08657_),
    .A2(_08659_),
    .B1(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__nor2_1 _15596_ (.A(_08367_),
    .B(_08557_),
    .Y(_08671_));
 sky130_fd_sc_hd__a21oi_1 _15597_ (.A1(_08548_),
    .A2(_08549_),
    .B1(_08347_),
    .Y(_08672_));
 sky130_fd_sc_hd__xor2_1 _15598_ (.A(_08671_),
    .B(_08672_),
    .X(_08673_));
 sky130_fd_sc_hd__nor2_1 _15599_ (.A(_08564_),
    .B(_08387_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_1 _15600_ (.A(_08673_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__or2_1 _15601_ (.A(_08673_),
    .B(_08674_),
    .X(_08676_));
 sky130_fd_sc_hd__and2_1 _15602_ (.A(_08675_),
    .B(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__nand3_1 _15603_ (.A(_08657_),
    .B(_08659_),
    .C(_08669_),
    .Y(_08678_));
 sky130_fd_sc_hd__a21boi_1 _15604_ (.A1(_08670_),
    .A2(_08677_),
    .B1_N(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__o21ai_2 _15605_ (.A1(_08652_),
    .A2(_08656_),
    .B1(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__or4_1 _15606_ (.A(_08529_),
    .B(_08393_),
    .C(_08405_),
    .D(_08422_),
    .X(_08681_));
 sky130_fd_sc_hd__o22ai_1 _15607_ (.A1(_08529_),
    .A2(_08449_),
    .B1(_08424_),
    .B2(_08394_),
    .Y(_08682_));
 sky130_fd_sc_hd__and2_1 _15608_ (.A(_08681_),
    .B(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__clkbuf_4 _15609_ (.A(_08444_),
    .X(_08684_));
 sky130_fd_sc_hd__nor2_1 _15610_ (.A(_08411_),
    .B(_08684_),
    .Y(_08685_));
 sky130_fd_sc_hd__nand2_1 _15611_ (.A(_08683_),
    .B(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_1 _15612_ (.A(_08681_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_1 _15613_ (.A(_08671_),
    .B(_08672_),
    .Y(_08688_));
 sky130_fd_sc_hd__nand2_1 _15614_ (.A(_08532_),
    .B(_08530_),
    .Y(_08689_));
 sky130_fd_sc_hd__xor2_1 _15615_ (.A(_08689_),
    .B(_08531_),
    .X(_08690_));
 sky130_fd_sc_hd__a21o_1 _15616_ (.A1(_08688_),
    .A2(_08675_),
    .B1(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__nand3_1 _15617_ (.A(_08688_),
    .B(_08675_),
    .C(_08690_),
    .Y(_08692_));
 sky130_fd_sc_hd__and2_1 _15618_ (.A(_08691_),
    .B(_08692_),
    .X(_08693_));
 sky130_fd_sc_hd__xor2_1 _15619_ (.A(_08687_),
    .B(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__or3_4 _15620_ (.A(_08652_),
    .B(_08656_),
    .C(_08679_),
    .X(_08695_));
 sky130_fd_sc_hd__a21boi_2 _15621_ (.A1(_08680_),
    .A2(_08694_),
    .B1_N(_08695_),
    .Y(_08696_));
 sky130_fd_sc_hd__xor2_1 _15622_ (.A(_08655_),
    .B(_08696_),
    .X(_08697_));
 sky130_fd_sc_hd__nor2_1 _15623_ (.A(_08313_),
    .B(_08315_),
    .Y(_08698_));
 sky130_fd_sc_hd__nand2_1 _15624_ (.A(_08698_),
    .B(_08490_),
    .Y(_08699_));
 sky130_fd_sc_hd__or2_1 _15625_ (.A(_08310_),
    .B(_08331_),
    .X(_08700_));
 sky130_fd_sc_hd__nor2_4 _15626_ (.A(_08328_),
    .B(_08329_),
    .Y(_08701_));
 sky130_fd_sc_hd__nand2_1 _15627_ (.A(_08701_),
    .B(_08490_),
    .Y(_08702_));
 sky130_fd_sc_hd__nor2_1 _15628_ (.A(_08318_),
    .B(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__a21o_1 _15629_ (.A1(_08699_),
    .A2(_08700_),
    .B1(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__nand2_4 _15630_ (.A(net6123),
    .B(_08314_),
    .Y(_08705_));
 sky130_fd_sc_hd__or2_1 _15631_ (.A(_08313_),
    .B(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__buf_2 _15632_ (.A(_08706_),
    .X(_08707_));
 sky130_fd_sc_hd__clkbuf_4 _15633_ (.A(_08707_),
    .X(_08708_));
 sky130_fd_sc_hd__nor2_1 _15634_ (.A(_08326_),
    .B(_08708_),
    .Y(_08709_));
 sky130_fd_sc_hd__xnor2_2 _15635_ (.A(_08704_),
    .B(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__or2_1 _15636_ (.A(_08410_),
    .B(_08470_),
    .X(_08711_));
 sky130_fd_sc_hd__or3_1 _15637_ (.A(_08433_),
    .B(_08484_),
    .C(_08711_),
    .X(_08712_));
 sky130_fd_sc_hd__o21ai_1 _15638_ (.A1(_08433_),
    .A2(_08516_),
    .B1(_08711_),
    .Y(_08713_));
 sky130_fd_sc_hd__and2_1 _15639_ (.A(_08712_),
    .B(_08713_),
    .X(_08714_));
 sky130_fd_sc_hd__nor2_1 _15640_ (.A(_08456_),
    .B(_08498_),
    .Y(_08715_));
 sky130_fd_sc_hd__xnor2_1 _15641_ (.A(_08714_),
    .B(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__buf_4 _15642_ (.A(_08498_),
    .X(_08717_));
 sky130_fd_sc_hd__nand2_1 _15643_ (.A(_08472_),
    .B(_08485_),
    .Y(_08718_));
 sky130_fd_sc_hd__o31a_1 _15644_ (.A1(_08486_),
    .A2(_08493_),
    .A3(_08717_),
    .B1(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__nand2_1 _15645_ (.A(_08716_),
    .B(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__nor2_1 _15646_ (.A(_08716_),
    .B(_08719_),
    .Y(_08721_));
 sky130_fd_sc_hd__a21o_1 _15647_ (.A1(_08710_),
    .A2(_08720_),
    .B1(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__nand2_1 _15648_ (.A(_08687_),
    .B(_08693_),
    .Y(_08723_));
 sky130_fd_sc_hd__clkbuf_4 _15649_ (.A(_08454_),
    .X(_08724_));
 sky130_fd_sc_hd__o21ai_1 _15650_ (.A1(_08317_),
    .A2(_08724_),
    .B1(_08702_),
    .Y(_08725_));
 sky130_fd_sc_hd__or3_2 _15651_ (.A(_08331_),
    .B(_08454_),
    .C(_08699_),
    .X(_08726_));
 sky130_fd_sc_hd__nor2_1 _15652_ (.A(_08310_),
    .B(_08707_),
    .Y(_08727_));
 sky130_fd_sc_hd__nand3_1 _15653_ (.A(_08725_),
    .B(_08726_),
    .C(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21o_1 _15654_ (.A1(_08725_),
    .A2(_08726_),
    .B1(_08727_),
    .X(_08729_));
 sky130_fd_sc_hd__and2_1 _15655_ (.A(_08728_),
    .B(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__or4_1 _15656_ (.A(_08394_),
    .B(_08411_),
    .C(_08470_),
    .D(_08484_),
    .X(_08731_));
 sky130_fd_sc_hd__o22ai_1 _15657_ (.A1(_08394_),
    .A2(_08471_),
    .B1(_08484_),
    .B2(_08411_),
    .Y(_08732_));
 sky130_fd_sc_hd__nand2_1 _15658_ (.A(_08731_),
    .B(_08732_),
    .Y(_08733_));
 sky130_fd_sc_hd__or2_1 _15659_ (.A(_08433_),
    .B(_08497_),
    .X(_08734_));
 sky130_fd_sc_hd__xnor2_1 _15660_ (.A(_08733_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__o21a_1 _15661_ (.A1(_08433_),
    .A2(_08516_),
    .B1(_08711_),
    .X(_08736_));
 sky130_fd_sc_hd__o31a_1 _15662_ (.A1(_08456_),
    .A2(_08498_),
    .A3(_08736_),
    .B1(_08712_),
    .X(_08737_));
 sky130_fd_sc_hd__nor2_1 _15663_ (.A(_08735_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__and2_1 _15664_ (.A(_08735_),
    .B(_08737_),
    .X(_08739_));
 sky130_fd_sc_hd__nor2_1 _15665_ (.A(_08738_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__xnor2_1 _15666_ (.A(_08730_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__a21o_1 _15667_ (.A1(_08691_),
    .A2(_08723_),
    .B1(_08741_),
    .X(_08742_));
 sky130_fd_sc_hd__nand3_1 _15668_ (.A(_08691_),
    .B(_08723_),
    .C(_08741_),
    .Y(_08743_));
 sky130_fd_sc_hd__nand2_1 _15669_ (.A(_08742_),
    .B(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__xnor2_1 _15670_ (.A(_08722_),
    .B(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__xnor2_1 _15671_ (.A(_08697_),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__and3_1 _15672_ (.A(_08695_),
    .B(_08680_),
    .C(_08694_),
    .X(_08747_));
 sky130_fd_sc_hd__a21oi_1 _15673_ (.A1(_08695_),
    .A2(_08680_),
    .B1(_08694_),
    .Y(_08748_));
 sky130_fd_sc_hd__or2_4 _15674_ (.A(_08747_),
    .B(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__nand2_1 _15675_ (.A(_08678_),
    .B(_08670_),
    .Y(_08750_));
 sky130_fd_sc_hd__xor2_2 _15676_ (.A(_08750_),
    .B(_08677_),
    .X(_08751_));
 sky130_fd_sc_hd__xnor2_2 _15677_ (.A(_08667_),
    .B(_08668_),
    .Y(_08752_));
 sky130_fd_sc_hd__or4b_2 _15678_ (.A(_08548_),
    .B(net4954),
    .C(_08664_),
    .D_N(_08540_),
    .X(_08753_));
 sky130_fd_sc_hd__a21oi_4 _15679_ (.A1(_08314_),
    .A2(_08546_),
    .B1(_08547_),
    .Y(_08754_));
 sky130_fd_sc_hd__nor2_4 _15680_ (.A(_08327_),
    .B(net7444),
    .Y(_08755_));
 sky130_fd_sc_hd__a22o_1 _15681_ (.A1(_08754_),
    .A2(_08631_),
    .B1(_08755_),
    .B2(_08540_),
    .X(_08756_));
 sky130_fd_sc_hd__nor2_1 _15682_ (.A(_08557_),
    .B(_08625_),
    .Y(_08757_));
 sky130_fd_sc_hd__nand3_1 _15683_ (.A(_08753_),
    .B(_08756_),
    .C(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__nand2_1 _15684_ (.A(_08753_),
    .B(_08758_),
    .Y(_08759_));
 sky130_fd_sc_hd__xnor2_2 _15685_ (.A(_08752_),
    .B(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__or4_1 _15686_ (.A(_08347_),
    .B(_08353_),
    .C(_08367_),
    .D(_08557_),
    .X(_08761_));
 sky130_fd_sc_hd__o22ai_2 _15687_ (.A1(_08564_),
    .A2(_08560_),
    .B1(_08565_),
    .B2(_08559_),
    .Y(_08762_));
 sky130_fd_sc_hd__nand2_1 _15688_ (.A(_08761_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__nor2_1 _15689_ (.A(_08529_),
    .B(_08587_),
    .Y(_08764_));
 sky130_fd_sc_hd__xnor2_2 _15690_ (.A(_08763_),
    .B(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__and2b_1 _15691_ (.A_N(_08752_),
    .B(_08759_),
    .X(_08766_));
 sky130_fd_sc_hd__a21oi_2 _15692_ (.A1(_08760_),
    .A2(_08765_),
    .B1(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__xor2_2 _15693_ (.A(_08751_),
    .B(_08767_),
    .X(_08768_));
 sky130_fd_sc_hd__a21bo_1 _15694_ (.A1(_08425_),
    .A2(_08445_),
    .B1_N(_08423_),
    .X(_08769_));
 sky130_fd_sc_hd__a21bo_1 _15695_ (.A1(_08762_),
    .A2(_08764_),
    .B1_N(_08761_),
    .X(_08770_));
 sky130_fd_sc_hd__or2_1 _15696_ (.A(_08683_),
    .B(_08685_),
    .X(_08771_));
 sky130_fd_sc_hd__nand2_1 _15697_ (.A(_08686_),
    .B(_08771_),
    .Y(_08772_));
 sky130_fd_sc_hd__xor2_2 _15698_ (.A(_08770_),
    .B(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__xnor2_2 _15699_ (.A(_08769_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__nor2_1 _15700_ (.A(_08751_),
    .B(_08767_),
    .Y(_08775_));
 sky130_fd_sc_hd__a21oi_2 _15701_ (.A1(_08768_),
    .A2(_08774_),
    .B1(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__xor2_4 _15702_ (.A(_08749_),
    .B(_08776_),
    .X(_08777_));
 sky130_fd_sc_hd__a21oi_2 _15703_ (.A1(_08463_),
    .A2(_08508_),
    .B1(_08507_),
    .Y(_08778_));
 sky130_fd_sc_hd__or2b_1 _15704_ (.A(_08772_),
    .B_N(_08770_),
    .X(_08779_));
 sky130_fd_sc_hd__or2b_1 _15705_ (.A(_08773_),
    .B_N(_08769_),
    .X(_08780_));
 sky130_fd_sc_hd__nand2_2 _15706_ (.A(_08779_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__and2b_1 _15707_ (.A_N(_08721_),
    .B(_08720_),
    .X(_08782_));
 sky130_fd_sc_hd__xnor2_2 _15708_ (.A(_08710_),
    .B(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__xnor2_2 _15709_ (.A(_08781_),
    .B(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__xnor2_2 _15710_ (.A(_08778_),
    .B(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__nor2_1 _15711_ (.A(_08749_),
    .B(_08776_),
    .Y(_08786_));
 sky130_fd_sc_hd__a21oi_2 _15712_ (.A1(_08777_),
    .A2(_08785_),
    .B1(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__nor2_2 _15713_ (.A(_08746_),
    .B(_08787_),
    .Y(_08788_));
 sky130_fd_sc_hd__and2_4 _15714_ (.A(_08746_),
    .B(_08787_),
    .X(_08789_));
 sky130_fd_sc_hd__nor2_4 _15715_ (.A(_08788_),
    .B(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__or2b_1 _15716_ (.A(_08783_),
    .B_N(_08781_),
    .X(_08791_));
 sky130_fd_sc_hd__or2b_1 _15717_ (.A(_08778_),
    .B_N(_08784_),
    .X(_08792_));
 sky130_fd_sc_hd__nand2_4 _15718_ (.A(net6098),
    .B(_08299_),
    .Y(_08793_));
 sky130_fd_sc_hd__or2_1 _15719_ (.A(_08312_),
    .B(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__clkbuf_4 _15720_ (.A(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__or2_1 _15721_ (.A(_08325_),
    .B(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__nand2_1 _15722_ (.A(_08699_),
    .B(_08700_),
    .Y(_08797_));
 sky130_fd_sc_hd__a21oi_1 _15723_ (.A1(_08797_),
    .A2(_08709_),
    .B1(_08703_),
    .Y(_08798_));
 sky130_fd_sc_hd__nor2_1 _15724_ (.A(_08796_),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__and2_1 _15725_ (.A(_08796_),
    .B(_08798_),
    .X(_08800_));
 sky130_fd_sc_hd__or2_1 _15726_ (.A(_08799_),
    .B(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__a21oi_2 _15727_ (.A1(_08791_),
    .A2(_08792_),
    .B1(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__and3_1 _15728_ (.A(_08791_),
    .B(_08792_),
    .C(_08801_),
    .X(_08803_));
 sky130_fd_sc_hd__nor2_2 _15729_ (.A(_08802_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__xnor2_4 _15730_ (.A(_08790_),
    .B(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__xnor2_2 _15731_ (.A(_08777_),
    .B(_08785_),
    .Y(_08806_));
 sky130_fd_sc_hd__xnor2_2 _15732_ (.A(_08768_),
    .B(_08774_),
    .Y(_08807_));
 sky130_fd_sc_hd__xnor2_2 _15733_ (.A(_08760_),
    .B(_08765_),
    .Y(_08808_));
 sky130_fd_sc_hd__a21o_1 _15734_ (.A1(_08753_),
    .A2(_08756_),
    .B1(_08757_),
    .X(_08809_));
 sky130_fd_sc_hd__nor2_1 _15735_ (.A(_08548_),
    .B(net4954),
    .Y(_08810_));
 sky130_fd_sc_hd__nor2_2 _15736_ (.A(_08556_),
    .B(net7444),
    .Y(_08811_));
 sky130_fd_sc_hd__nor2_1 _15737_ (.A(_08353_),
    .B(_08625_),
    .Y(_08812_));
 sky130_fd_sc_hd__or2_1 _15738_ (.A(_08556_),
    .B(net4954),
    .X(_08813_));
 sky130_fd_sc_hd__or4_2 _15739_ (.A(net3722),
    .B(_08379_),
    .C(_08546_),
    .D(_08547_),
    .X(_08814_));
 sky130_fd_sc_hd__a32oi_4 _15740_ (.A1(_08754_),
    .A2(_08631_),
    .A3(_08811_),
    .B1(_08813_),
    .B2(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__a22o_1 _15741_ (.A1(_08810_),
    .A2(_08811_),
    .B1(_08812_),
    .B2(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__nand3_1 _15742_ (.A(_08758_),
    .B(_08809_),
    .C(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__a21o_1 _15743_ (.A1(_08758_),
    .A2(_08809_),
    .B1(_08816_),
    .X(_08818_));
 sky130_fd_sc_hd__and2_1 _15744_ (.A(_08396_),
    .B(_08374_),
    .X(_08819_));
 sky130_fd_sc_hd__xor2_1 _15745_ (.A(_08819_),
    .B(_08395_),
    .X(_08820_));
 sky130_fd_sc_hd__nand3_1 _15746_ (.A(_08817_),
    .B(_08818_),
    .C(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__and2_1 _15747_ (.A(_08817_),
    .B(_08821_),
    .X(_08822_));
 sky130_fd_sc_hd__xor2_2 _15748_ (.A(_08808_),
    .B(_08822_),
    .X(_08823_));
 sky130_fd_sc_hd__xnor2_2 _15749_ (.A(_08459_),
    .B(_08447_),
    .Y(_08824_));
 sky130_fd_sc_hd__nor2_1 _15750_ (.A(_08808_),
    .B(_08822_),
    .Y(_08825_));
 sky130_fd_sc_hd__a21oi_2 _15751_ (.A1(_08823_),
    .A2(_08824_),
    .B1(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__xor2_2 _15752_ (.A(_08807_),
    .B(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__xnor2_2 _15753_ (.A(_08524_),
    .B(_08511_),
    .Y(_08828_));
 sky130_fd_sc_hd__nor2_1 _15754_ (.A(_08807_),
    .B(_08826_),
    .Y(_08829_));
 sky130_fd_sc_hd__a21oi_2 _15755_ (.A1(_08827_),
    .A2(_08828_),
    .B1(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__xor2_1 _15756_ (.A(_08806_),
    .B(_08830_),
    .X(_08831_));
 sky130_fd_sc_hd__xor2_1 _15757_ (.A(_08332_),
    .B(_08526_),
    .X(_08832_));
 sky130_fd_sc_hd__nand2_2 _15758_ (.A(_08831_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__o21ai_4 _15759_ (.A1(_08806_),
    .A2(_08830_),
    .B1(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__xnor2_4 _15760_ (.A(_08805_),
    .B(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__xnor2_4 _15761_ (.A(_08528_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__xnor2_2 _15762_ (.A(_08827_),
    .B(_08828_),
    .Y(_08837_));
 sky130_fd_sc_hd__xnor2_2 _15763_ (.A(_08823_),
    .B(_08824_),
    .Y(_08838_));
 sky130_fd_sc_hd__a21o_1 _15764_ (.A1(_08817_),
    .A2(_08818_),
    .B1(_08820_),
    .X(_08839_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_08387_),
    .B(_08411_),
    .Y(_08840_));
 sky130_fd_sc_hd__or2_1 _15766_ (.A(_08347_),
    .B(_08373_),
    .X(_08841_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_08367_),
    .B(_08393_),
    .Y(_08842_));
 sky130_fd_sc_hd__xnor2_1 _15768_ (.A(_08841_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__xor2_1 _15769_ (.A(_08840_),
    .B(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__xor2_1 _15770_ (.A(_08812_),
    .B(_08815_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _15771_ (.A(_08373_),
    .B(_08625_),
    .Y(_08846_));
 sky130_fd_sc_hd__or4_1 _15772_ (.A(net3539),
    .B(_08311_),
    .C(_08305_),
    .D(_08351_),
    .X(_08847_));
 sky130_fd_sc_hd__xnor2_1 _15773_ (.A(_08811_),
    .B(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand2_8 _15774_ (.A(_08351_),
    .B(_08352_),
    .Y(_08849_));
 sky130_fd_sc_hd__and3_1 _15775_ (.A(_08849_),
    .B(_08665_),
    .C(_08811_),
    .X(_08850_));
 sky130_fd_sc_hd__a21o_1 _15776_ (.A1(_08846_),
    .A2(_08848_),
    .B1(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__xor2_1 _15777_ (.A(_08845_),
    .B(_08851_),
    .X(_08852_));
 sky130_fd_sc_hd__and2_1 _15778_ (.A(_08845_),
    .B(_08851_),
    .X(_08853_));
 sky130_fd_sc_hd__a21o_1 _15779_ (.A1(_08844_),
    .A2(_08852_),
    .B1(_08853_),
    .X(_08854_));
 sky130_fd_sc_hd__nand3_1 _15780_ (.A(_08821_),
    .B(_08839_),
    .C(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__a21o_1 _15781_ (.A1(_08821_),
    .A2(_08839_),
    .B1(_08854_),
    .X(_08856_));
 sky130_fd_sc_hd__or4_1 _15782_ (.A(_08405_),
    .B(_08422_),
    .C(_08432_),
    .D(_08455_),
    .X(_08857_));
 sky130_fd_sc_hd__nor2_1 _15783_ (.A(_08444_),
    .B(_08493_),
    .Y(_08858_));
 sky130_fd_sc_hd__o22ai_2 _15784_ (.A1(_08449_),
    .A2(_08433_),
    .B1(_08456_),
    .B2(_08424_),
    .Y(_08859_));
 sky130_fd_sc_hd__nand3_1 _15785_ (.A(_08857_),
    .B(_08858_),
    .C(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__nand2_1 _15786_ (.A(_08857_),
    .B(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__or3_1 _15787_ (.A(_08560_),
    .B(_08394_),
    .C(_08841_),
    .X(_08862_));
 sky130_fd_sc_hd__a21bo_1 _15788_ (.A1(_08840_),
    .A2(_08843_),
    .B1_N(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__a21o_1 _15789_ (.A1(_08448_),
    .A2(_08450_),
    .B1(_08457_),
    .X(_08864_));
 sky130_fd_sc_hd__nand3_1 _15790_ (.A(_08458_),
    .B(_08863_),
    .C(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__a21o_1 _15791_ (.A1(_08458_),
    .A2(_08864_),
    .B1(_08863_),
    .X(_08866_));
 sky130_fd_sc_hd__nand3_1 _15792_ (.A(_08861_),
    .B(_08865_),
    .C(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__a21o_1 _15793_ (.A1(_08865_),
    .A2(_08866_),
    .B1(_08861_),
    .X(_08868_));
 sky130_fd_sc_hd__nand4_1 _15794_ (.A(_08855_),
    .B(_08856_),
    .C(_08867_),
    .D(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__and2_1 _15795_ (.A(_08855_),
    .B(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__xor2_2 _15796_ (.A(_08838_),
    .B(_08870_),
    .X(_08871_));
 sky130_fd_sc_hd__buf_4 _15797_ (.A(_08471_),
    .X(_08872_));
 sky130_fd_sc_hd__buf_4 _15798_ (.A(_08516_),
    .X(_08873_));
 sky130_fd_sc_hd__clkbuf_4 _15799_ (.A(_08514_),
    .X(_08874_));
 sky130_fd_sc_hd__or4_2 _15800_ (.A(_08872_),
    .B(_08873_),
    .C(_08517_),
    .D(_08874_),
    .X(_08875_));
 sky130_fd_sc_hd__nor2_1 _15801_ (.A(_08516_),
    .B(_08517_),
    .Y(_08876_));
 sky130_fd_sc_hd__xnor2_1 _15802_ (.A(_08518_),
    .B(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__xnor2_1 _15803_ (.A(_08515_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__or2b_1 _15804_ (.A(_08875_),
    .B_N(_08878_),
    .X(_08879_));
 sky130_fd_sc_hd__nand2_1 _15805_ (.A(_08865_),
    .B(_08867_),
    .Y(_08880_));
 sky130_fd_sc_hd__xnor2_1 _15806_ (.A(_08512_),
    .B(_08522_),
    .Y(_08881_));
 sky130_fd_sc_hd__xnor2_2 _15807_ (.A(_08880_),
    .B(_08881_),
    .Y(_08882_));
 sky130_fd_sc_hd__xnor2_2 _15808_ (.A(_08879_),
    .B(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__nor2_1 _15809_ (.A(_08838_),
    .B(_08870_),
    .Y(_08884_));
 sky130_fd_sc_hd__a21oi_2 _15810_ (.A1(_08871_),
    .A2(_08883_),
    .B1(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__xnor2_2 _15811_ (.A(_08837_),
    .B(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__and2b_1 _15812_ (.A_N(_08881_),
    .B(_08880_),
    .X(_08887_));
 sky130_fd_sc_hd__and2b_1 _15813_ (.A_N(_08879_),
    .B(_08882_),
    .X(_08888_));
 sky130_fd_sc_hd__nor2_1 _15814_ (.A(_08887_),
    .B(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__xnor2_2 _15815_ (.A(_08886_),
    .B(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__nor2_1 _15816_ (.A(_08387_),
    .B(_08432_),
    .Y(_08891_));
 sky130_fd_sc_hd__nor2_1 _15817_ (.A(_08347_),
    .B(_08393_),
    .Y(_08892_));
 sky130_fd_sc_hd__nor2_1 _15818_ (.A(_08367_),
    .B(_08410_),
    .Y(_08893_));
 sky130_fd_sc_hd__xor2_2 _15819_ (.A(_08892_),
    .B(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__and2_1 _15820_ (.A(_08892_),
    .B(_08893_),
    .X(_08895_));
 sky130_fd_sc_hd__a21o_1 _15821_ (.A1(_08891_),
    .A2(_08894_),
    .B1(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__a21o_1 _15822_ (.A1(_08857_),
    .A2(_08859_),
    .B1(_08858_),
    .X(_08897_));
 sky130_fd_sc_hd__nand3_2 _15823_ (.A(_08860_),
    .B(_08896_),
    .C(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__inv_2 _15824_ (.A(_08422_),
    .Y(_08899_));
 sky130_fd_sc_hd__and3_1 _15825_ (.A(_08899_),
    .B(_08490_),
    .C(_08491_),
    .X(_08900_));
 sky130_fd_sc_hd__nor2_1 _15826_ (.A(_08405_),
    .B(_08455_),
    .Y(_08901_));
 sky130_fd_sc_hd__or2_1 _15827_ (.A(_08444_),
    .B(_08501_),
    .X(_08902_));
 sky130_fd_sc_hd__xor2_1 _15828_ (.A(_08900_),
    .B(_08901_),
    .X(_08903_));
 sky130_fd_sc_hd__or2b_1 _15829_ (.A(_08902_),
    .B_N(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__a21bo_1 _15830_ (.A1(_08900_),
    .A2(_08901_),
    .B1_N(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__a21o_1 _15831_ (.A1(_08860_),
    .A2(_08897_),
    .B1(_08896_),
    .X(_08906_));
 sky130_fd_sc_hd__nand3_2 _15832_ (.A(_08905_),
    .B(_08898_),
    .C(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__xor2_1 _15833_ (.A(_08875_),
    .B(_08878_),
    .X(_08908_));
 sky130_fd_sc_hd__a21oi_2 _15834_ (.A1(_08898_),
    .A2(_08907_),
    .B1(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__xnor2_2 _15835_ (.A(_08871_),
    .B(_08883_),
    .Y(_08910_));
 sky130_fd_sc_hd__a22o_1 _15836_ (.A1(_08855_),
    .A2(_08856_),
    .B1(_08867_),
    .B2(_08868_),
    .X(_08911_));
 sky130_fd_sc_hd__a21o_1 _15837_ (.A1(_08898_),
    .A2(_08906_),
    .B1(_08905_),
    .X(_08912_));
 sky130_fd_sc_hd__xnor2_1 _15838_ (.A(_08844_),
    .B(_08852_),
    .Y(_08913_));
 sky130_fd_sc_hd__xor2_2 _15839_ (.A(_08891_),
    .B(_08894_),
    .X(_08914_));
 sky130_fd_sc_hd__xnor2_1 _15840_ (.A(_08846_),
    .B(_08848_),
    .Y(_08915_));
 sky130_fd_sc_hd__nor2_1 _15841_ (.A(_08393_),
    .B(_08625_),
    .Y(_08916_));
 sky130_fd_sc_hd__nor2_2 _15842_ (.A(_08372_),
    .B(_08663_),
    .Y(_08917_));
 sky130_fd_sc_hd__or2_1 _15843_ (.A(_08372_),
    .B(_08632_),
    .X(_08918_));
 sky130_fd_sc_hd__or4_1 _15844_ (.A(net3722),
    .B(_08311_),
    .C(_08305_),
    .D(_08351_),
    .X(_08919_));
 sky130_fd_sc_hd__a32oi_4 _15845_ (.A1(_08849_),
    .A2(_08665_),
    .A3(_08917_),
    .B1(_08918_),
    .B2(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__and3_1 _15846_ (.A(_08849_),
    .B(_08665_),
    .C(_08917_),
    .X(_08921_));
 sky130_fd_sc_hd__a21o_1 _15847_ (.A1(_08916_),
    .A2(_08920_),
    .B1(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__xnor2_1 _15848_ (.A(_08915_),
    .B(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__or2b_1 _15849_ (.A(_08915_),
    .B_N(_08922_),
    .X(_08924_));
 sky130_fd_sc_hd__a21bo_1 _15850_ (.A1(_08914_),
    .A2(_08923_),
    .B1_N(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__xnor2_1 _15851_ (.A(_08913_),
    .B(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__and2b_1 _15852_ (.A_N(_08913_),
    .B(_08925_),
    .X(_08927_));
 sky130_fd_sc_hd__a31o_1 _15853_ (.A1(_08907_),
    .A2(_08912_),
    .A3(_08926_),
    .B1(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__nand3_1 _15854_ (.A(_08869_),
    .B(_08911_),
    .C(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__a21o_1 _15855_ (.A1(_08869_),
    .A2(_08911_),
    .B1(_08928_),
    .X(_08930_));
 sky130_fd_sc_hd__and3_1 _15856_ (.A(_08898_),
    .B(_08907_),
    .C(_08908_),
    .X(_08931_));
 sky130_fd_sc_hd__nor2_1 _15857_ (.A(_08909_),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand3_1 _15858_ (.A(_08929_),
    .B(_08930_),
    .C(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__and2_1 _15859_ (.A(_08929_),
    .B(_08933_),
    .X(_08934_));
 sky130_fd_sc_hd__xor2_2 _15860_ (.A(_08910_),
    .B(_08934_),
    .X(_08935_));
 sky130_fd_sc_hd__nor2_1 _15861_ (.A(_08910_),
    .B(_08934_),
    .Y(_08936_));
 sky130_fd_sc_hd__a21oi_2 _15862_ (.A1(_08909_),
    .A2(_08935_),
    .B1(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__nor2_1 _15863_ (.A(_08890_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__or2_4 _15864_ (.A(_08831_),
    .B(_08832_),
    .X(_08939_));
 sky130_fd_sc_hd__nand2_2 _15865_ (.A(_08833_),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__or2_1 _15866_ (.A(_08837_),
    .B(_08885_),
    .X(_08941_));
 sky130_fd_sc_hd__o21a_1 _15867_ (.A1(_08886_),
    .A2(_08889_),
    .B1(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__nor2_4 _15868_ (.A(_08940_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_2 _15869_ (.A(_08940_),
    .B(_08942_),
    .Y(_08944_));
 sky130_fd_sc_hd__nor2b_4 _15870_ (.A(_08943_),
    .B_N(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__nand2_1 _15871_ (.A(_08938_),
    .B(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__xnor2_2 _15872_ (.A(_08909_),
    .B(_08935_),
    .Y(_08947_));
 sky130_fd_sc_hd__a21o_1 _15873_ (.A1(_08929_),
    .A2(_08930_),
    .B1(_08932_),
    .X(_08948_));
 sky130_fd_sc_hd__nand3_1 _15874_ (.A(_08907_),
    .B(_08912_),
    .C(_08926_),
    .Y(_08949_));
 sky130_fd_sc_hd__a21o_1 _15875_ (.A1(_08907_),
    .A2(_08912_),
    .B1(_08926_),
    .X(_08950_));
 sky130_fd_sc_hd__xnor2_1 _15876_ (.A(_08914_),
    .B(_08923_),
    .Y(_08951_));
 sky130_fd_sc_hd__nor2_1 _15877_ (.A(_08387_),
    .B(_08456_),
    .Y(_08952_));
 sky130_fd_sc_hd__or4_1 _15878_ (.A(_08347_),
    .B(_08366_),
    .C(_08410_),
    .D(_08432_),
    .X(_08953_));
 sky130_fd_sc_hd__o22ai_2 _15879_ (.A1(_08559_),
    .A2(_08411_),
    .B1(_08432_),
    .B2(_08367_),
    .Y(_08954_));
 sky130_fd_sc_hd__and3_1 _15880_ (.A(_08952_),
    .B(_08953_),
    .C(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__a21oi_1 _15881_ (.A1(_08953_),
    .A2(_08954_),
    .B1(_08952_),
    .Y(_08956_));
 sky130_fd_sc_hd__xnor2_1 _15882_ (.A(_08916_),
    .B(_08920_),
    .Y(_08957_));
 sky130_fd_sc_hd__nor2_1 _15883_ (.A(_08410_),
    .B(_08625_),
    .Y(_08958_));
 sky130_fd_sc_hd__or4_1 _15884_ (.A(net3539),
    .B(_08311_),
    .C(_08379_),
    .D(_08391_),
    .X(_08959_));
 sky130_fd_sc_hd__xnor2_1 _15885_ (.A(_08917_),
    .B(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__nand2_1 _15886_ (.A(_08391_),
    .B(_08392_),
    .Y(_08961_));
 sky130_fd_sc_hd__clkbuf_4 _15887_ (.A(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__and3_1 _15888_ (.A(_08962_),
    .B(_08665_),
    .C(_08917_),
    .X(_08963_));
 sky130_fd_sc_hd__a21oi_1 _15889_ (.A1(_08958_),
    .A2(_08960_),
    .B1(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__xnor2_1 _15890_ (.A(_08957_),
    .B(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__o32a_1 _15891_ (.A1(_08955_),
    .A2(_08956_),
    .A3(_08965_),
    .B1(_08964_),
    .B2(_08957_),
    .X(_08966_));
 sky130_fd_sc_hd__nor2_1 _15892_ (.A(_08951_),
    .B(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__nor2_1 _15893_ (.A(_08444_),
    .B(_08514_),
    .Y(_08968_));
 sky130_fd_sc_hd__inv_2 _15894_ (.A(_08404_),
    .Y(_08969_));
 sky130_fd_sc_hd__and3_1 _15895_ (.A(_08969_),
    .B(_08490_),
    .C(_08491_),
    .X(_08970_));
 sky130_fd_sc_hd__nor2_1 _15896_ (.A(_08422_),
    .B(_08501_),
    .Y(_08971_));
 sky130_fd_sc_hd__xor2_1 _15897_ (.A(_08970_),
    .B(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__nand2_1 _15898_ (.A(_08970_),
    .B(_08971_),
    .Y(_08973_));
 sky130_fd_sc_hd__a21bo_1 _15899_ (.A1(_08968_),
    .A2(_08972_),
    .B1_N(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__a21bo_1 _15900_ (.A1(_08952_),
    .A2(_08954_),
    .B1_N(_08953_),
    .X(_08975_));
 sky130_fd_sc_hd__xnor2_1 _15901_ (.A(_08902_),
    .B(_08903_),
    .Y(_08976_));
 sky130_fd_sc_hd__xnor2_1 _15902_ (.A(_08975_),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__xnor2_1 _15903_ (.A(_08974_),
    .B(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__xor2_1 _15904_ (.A(_08951_),
    .B(_08966_),
    .X(_08979_));
 sky130_fd_sc_hd__and2_1 _15905_ (.A(_08978_),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__a211o_1 _15906_ (.A1(_08949_),
    .A2(_08950_),
    .B1(_08967_),
    .C1(_08980_),
    .X(_08981_));
 sky130_fd_sc_hd__or2b_1 _15907_ (.A(_08977_),
    .B_N(_08974_),
    .X(_08982_));
 sky130_fd_sc_hd__a21bo_1 _15908_ (.A1(_08975_),
    .A2(_08976_),
    .B1_N(_08982_),
    .X(_08983_));
 sky130_fd_sc_hd__o22ai_1 _15909_ (.A1(_08872_),
    .A2(_08517_),
    .B1(_08874_),
    .B2(_08873_),
    .Y(_08984_));
 sky130_fd_sc_hd__nand2_1 _15910_ (.A(_08875_),
    .B(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__xnor2_1 _15911_ (.A(_08983_),
    .B(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__o211ai_2 _15912_ (.A1(_08967_),
    .A2(_08980_),
    .B1(_08949_),
    .C1(_08950_),
    .Y(_08987_));
 sky130_fd_sc_hd__a21bo_1 _15913_ (.A1(_08981_),
    .A2(_08986_),
    .B1_N(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__nand3_1 _15914_ (.A(_08933_),
    .B(_08948_),
    .C(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__and3_1 _15915_ (.A(_08875_),
    .B(_08983_),
    .C(_08984_),
    .X(_08990_));
 sky130_fd_sc_hd__a21o_1 _15916_ (.A1(_08933_),
    .A2(_08948_),
    .B1(_08988_),
    .X(_08991_));
 sky130_fd_sc_hd__nand3_1 _15917_ (.A(_08990_),
    .B(_08989_),
    .C(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__and2_1 _15918_ (.A(_08989_),
    .B(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__nor2_1 _15919_ (.A(_08947_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__xor2_2 _15920_ (.A(_08890_),
    .B(_08937_),
    .X(_08995_));
 sky130_fd_sc_hd__and2_1 _15921_ (.A(_08994_),
    .B(_08995_),
    .X(_08996_));
 sky130_fd_sc_hd__xnor2_2 _15922_ (.A(_08947_),
    .B(_08993_),
    .Y(_08997_));
 sky130_fd_sc_hd__a21o_1 _15923_ (.A1(_08989_),
    .A2(_08991_),
    .B1(_08990_),
    .X(_08998_));
 sky130_fd_sc_hd__nor2_1 _15924_ (.A(_08387_),
    .B(_08493_),
    .Y(_08999_));
 sky130_fd_sc_hd__o22ai_2 _15925_ (.A1(_08559_),
    .A2(_08433_),
    .B1(_08456_),
    .B2(_08560_),
    .Y(_09000_));
 sky130_fd_sc_hd__or4_1 _15926_ (.A(_08347_),
    .B(_08367_),
    .C(_08432_),
    .D(_08455_),
    .X(_09001_));
 sky130_fd_sc_hd__a21boi_2 _15927_ (.A1(_08999_),
    .A2(_09000_),
    .B1_N(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__xnor2_1 _15928_ (.A(_08968_),
    .B(_08972_),
    .Y(_09003_));
 sky130_fd_sc_hd__xor2_1 _15929_ (.A(_09002_),
    .B(_09003_),
    .X(_09004_));
 sky130_fd_sc_hd__and4bb_1 _15930_ (.A_N(_08514_),
    .B_N(_08501_),
    .C(_08899_),
    .D(_08969_),
    .X(_09005_));
 sky130_fd_sc_hd__nor2_1 _15931_ (.A(_09002_),
    .B(_09003_),
    .Y(_09006_));
 sky130_fd_sc_hd__a21oi_1 _15932_ (.A1(_09004_),
    .A2(_09005_),
    .B1(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__nor2_1 _15933_ (.A(_08872_),
    .B(_08874_),
    .Y(_09008_));
 sky130_fd_sc_hd__and2b_1 _15934_ (.A_N(_09007_),
    .B(_09008_),
    .X(_09009_));
 sky130_fd_sc_hd__nand3_1 _15935_ (.A(_08987_),
    .B(_08981_),
    .C(_08986_),
    .Y(_09010_));
 sky130_fd_sc_hd__a21o_1 _15936_ (.A1(_08987_),
    .A2(_08981_),
    .B1(_08986_),
    .X(_09011_));
 sky130_fd_sc_hd__xnor2_1 _15937_ (.A(_09008_),
    .B(_09007_),
    .Y(_09012_));
 sky130_fd_sc_hd__xnor2_1 _15938_ (.A(_08978_),
    .B(_08979_),
    .Y(_09013_));
 sky130_fd_sc_hd__xor2_1 _15939_ (.A(_09004_),
    .B(_09005_),
    .X(_09014_));
 sky130_fd_sc_hd__or3_1 _15940_ (.A(_08955_),
    .B(_08956_),
    .C(_08965_),
    .X(_09015_));
 sky130_fd_sc_hd__o21ai_1 _15941_ (.A1(_08955_),
    .A2(_08956_),
    .B1(_08965_),
    .Y(_09016_));
 sky130_fd_sc_hd__nand3_1 _15942_ (.A(_08999_),
    .B(_09000_),
    .C(_09001_),
    .Y(_09017_));
 sky130_fd_sc_hd__a21o_1 _15943_ (.A1(_09000_),
    .A2(_09001_),
    .B1(_08999_),
    .X(_09018_));
 sky130_fd_sc_hd__xnor2_1 _15944_ (.A(_08958_),
    .B(_08960_),
    .Y(_09019_));
 sky130_fd_sc_hd__or2_1 _15945_ (.A(_08409_),
    .B(_08632_),
    .X(_09020_));
 sky130_fd_sc_hd__a21boi_1 _15946_ (.A1(_08962_),
    .A2(_08755_),
    .B1_N(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__or3b_1 _15947_ (.A(_08664_),
    .B(_09020_),
    .C_N(_08961_),
    .X(_09022_));
 sky130_fd_sc_hd__o31a_1 _15948_ (.A1(_08432_),
    .A2(_08626_),
    .A3(_09021_),
    .B1(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__xor2_1 _15949_ (.A(_09019_),
    .B(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__nor2_1 _15950_ (.A(_09019_),
    .B(_09023_),
    .Y(_09025_));
 sky130_fd_sc_hd__a31o_1 _15951_ (.A1(_09017_),
    .A2(_09018_),
    .A3(_09024_),
    .B1(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__a21o_1 _15952_ (.A1(_09015_),
    .A2(_09016_),
    .B1(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__and3_1 _15953_ (.A(_09015_),
    .B(_09016_),
    .C(_09026_),
    .X(_09028_));
 sky130_fd_sc_hd__a21oi_1 _15954_ (.A1(_09014_),
    .A2(_09027_),
    .B1(_09028_),
    .Y(_09029_));
 sky130_fd_sc_hd__xor2_1 _15955_ (.A(_09013_),
    .B(_09029_),
    .X(_09030_));
 sky130_fd_sc_hd__nor2_1 _15956_ (.A(_09013_),
    .B(_09029_),
    .Y(_09031_));
 sky130_fd_sc_hd__a21o_1 _15957_ (.A1(_09012_),
    .A2(_09030_),
    .B1(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__a21o_1 _15958_ (.A1(_09010_),
    .A2(_09011_),
    .B1(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__and3_1 _15959_ (.A(_09010_),
    .B(_09011_),
    .C(_09032_),
    .X(_09034_));
 sky130_fd_sc_hd__a21o_1 _15960_ (.A1(_09009_),
    .A2(_09033_),
    .B1(_09034_),
    .X(_09035_));
 sky130_fd_sc_hd__nand3_2 _15961_ (.A(_08992_),
    .B(_08998_),
    .C(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__a21o_1 _15962_ (.A1(_08992_),
    .A2(_08998_),
    .B1(_09035_),
    .X(_09037_));
 sky130_fd_sc_hd__or2b_1 _15963_ (.A(_09034_),
    .B_N(_09033_),
    .X(_09038_));
 sky130_fd_sc_hd__xnor2_2 _15964_ (.A(_09009_),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__and2b_1 _15965_ (.A_N(_09028_),
    .B(_09027_),
    .X(_09040_));
 sky130_fd_sc_hd__xnor2_1 _15966_ (.A(_09014_),
    .B(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__and3_1 _15967_ (.A(_09017_),
    .B(_09018_),
    .C(_09024_),
    .X(_09042_));
 sky130_fd_sc_hd__a21oi_1 _15968_ (.A1(_09017_),
    .A2(_09018_),
    .B1(_09024_),
    .Y(_09043_));
 sky130_fd_sc_hd__or4b_1 _15969_ (.A(_08432_),
    .B(_09021_),
    .C(_08625_),
    .D_N(_09022_),
    .X(_09044_));
 sky130_fd_sc_hd__a21bo_1 _15970_ (.A1(_08962_),
    .A2(_08755_),
    .B1_N(_09020_),
    .X(_09045_));
 sky130_fd_sc_hd__a2bb2o_1 _15971_ (.A1_N(_08432_),
    .A2_N(_08626_),
    .B1(_09022_),
    .B2(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__nand2_1 _15972_ (.A(_09044_),
    .B(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__nor2_1 _15973_ (.A(_08456_),
    .B(_08626_),
    .Y(_09048_));
 sky130_fd_sc_hd__or2_1 _15974_ (.A(_08409_),
    .B(_08664_),
    .X(_09049_));
 sky130_fd_sc_hd__o41ai_2 _15975_ (.A1(net3539),
    .A2(_08313_),
    .A3(_08628_),
    .A4(_08430_),
    .B1(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__nand2_4 _15976_ (.A(_08430_),
    .B(_08431_),
    .Y(_09051_));
 sky130_fd_sc_hd__nand2_1 _15977_ (.A(_09051_),
    .B(_08755_),
    .Y(_09052_));
 sky130_fd_sc_hd__o2bb2a_1 _15978_ (.A1_N(_09048_),
    .A2_N(_09050_),
    .B1(_09020_),
    .B2(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__xor2_1 _15979_ (.A(_09047_),
    .B(_09053_),
    .X(_09054_));
 sky130_fd_sc_hd__or2_1 _15980_ (.A(_08587_),
    .B(_08501_),
    .X(_09055_));
 sky130_fd_sc_hd__o22a_1 _15981_ (.A1(_08559_),
    .A2(_08456_),
    .B1(_08493_),
    .B2(_08560_),
    .X(_09056_));
 sky130_fd_sc_hd__or4_1 _15982_ (.A(_08347_),
    .B(_08367_),
    .C(_08455_),
    .D(_08492_),
    .X(_09057_));
 sky130_fd_sc_hd__and2b_1 _15983_ (.A_N(_09056_),
    .B(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__xnor2_1 _15984_ (.A(_09055_),
    .B(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__nor2_1 _15985_ (.A(_09047_),
    .B(_09053_),
    .Y(_09060_));
 sky130_fd_sc_hd__a21oi_1 _15986_ (.A1(_09054_),
    .A2(_09059_),
    .B1(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__o21ai_1 _15987_ (.A1(_09042_),
    .A2(_09043_),
    .B1(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__o21a_1 _15988_ (.A1(_09055_),
    .A2(_09056_),
    .B1(_09057_),
    .X(_09063_));
 sky130_fd_sc_hd__clkbuf_4 _15989_ (.A(_08424_),
    .X(_09064_));
 sky130_fd_sc_hd__o22a_1 _15990_ (.A1(_08449_),
    .A2(_08501_),
    .B1(_08514_),
    .B2(_09064_),
    .X(_09065_));
 sky130_fd_sc_hd__or2_1 _15991_ (.A(_09005_),
    .B(_09065_),
    .X(_09066_));
 sky130_fd_sc_hd__or2_1 _15992_ (.A(_09063_),
    .B(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__nand2_1 _15993_ (.A(_09063_),
    .B(_09066_),
    .Y(_09068_));
 sky130_fd_sc_hd__and2_1 _15994_ (.A(_09067_),
    .B(_09068_),
    .X(_09069_));
 sky130_fd_sc_hd__or3_1 _15995_ (.A(_09042_),
    .B(_09043_),
    .C(_09061_),
    .X(_09070_));
 sky130_fd_sc_hd__a21boi_1 _15996_ (.A1(_09062_),
    .A2(_09069_),
    .B1_N(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__or2_1 _15997_ (.A(_09041_),
    .B(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__xnor2_1 _15998_ (.A(_09041_),
    .B(_09071_),
    .Y(_09073_));
 sky130_fd_sc_hd__or2_1 _15999_ (.A(_09067_),
    .B(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__xnor2_1 _16000_ (.A(_09012_),
    .B(_09030_),
    .Y(_09075_));
 sky130_fd_sc_hd__a21o_1 _16001_ (.A1(_09072_),
    .A2(_09074_),
    .B1(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__inv_2 _16002_ (.A(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__nand4_2 _16003_ (.A(_09036_),
    .B(_09037_),
    .C(_09039_),
    .D(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__a22o_1 _16004_ (.A1(_09036_),
    .A2(_09037_),
    .B1(_09039_),
    .B2(_09077_),
    .X(_09079_));
 sky130_fd_sc_hd__and3_1 _16005_ (.A(_09070_),
    .B(_09062_),
    .C(_09069_),
    .X(_09080_));
 sky130_fd_sc_hd__a21oi_1 _16006_ (.A1(_09070_),
    .A2(_09062_),
    .B1(_09069_),
    .Y(_09081_));
 sky130_fd_sc_hd__or2_1 _16007_ (.A(_09080_),
    .B(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_09054_),
    .B(_09059_),
    .Y(_09083_));
 sky130_fd_sc_hd__or2_1 _16009_ (.A(_08587_),
    .B(_08874_),
    .X(_09084_));
 sky130_fd_sc_hd__or2_1 _16010_ (.A(_08559_),
    .B(_08493_),
    .X(_09085_));
 sky130_fd_sc_hd__clkbuf_4 _16011_ (.A(_08560_),
    .X(_09086_));
 sky130_fd_sc_hd__nor2_1 _16012_ (.A(_09086_),
    .B(_08517_),
    .Y(_09087_));
 sky130_fd_sc_hd__xnor2_1 _16013_ (.A(_09085_),
    .B(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__xnor2_1 _16014_ (.A(_09084_),
    .B(_09088_),
    .Y(_09089_));
 sky130_fd_sc_hd__and2_1 _16015_ (.A(_08430_),
    .B(_08431_),
    .X(_09090_));
 sky130_fd_sc_hd__clkbuf_4 _16016_ (.A(_09090_),
    .X(_09091_));
 sky130_fd_sc_hd__o31a_1 _16017_ (.A1(_09091_),
    .A2(_08664_),
    .A3(_09020_),
    .B1(_09050_),
    .X(_09092_));
 sky130_fd_sc_hd__xnor2_1 _16018_ (.A(_09048_),
    .B(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__nor2_1 _16019_ (.A(_08454_),
    .B(_08632_),
    .Y(_09094_));
 sky130_fd_sc_hd__or3b_2 _16020_ (.A(_09090_),
    .B(_08664_),
    .C_N(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__clkbuf_4 _16021_ (.A(_08626_),
    .X(_09096_));
 sky130_fd_sc_hd__a21o_1 _16022_ (.A1(_09051_),
    .A2(_08755_),
    .B1(_09094_),
    .X(_09097_));
 sky130_fd_sc_hd__or4bb_1 _16023_ (.A(_08493_),
    .B(_09096_),
    .C_N(_09095_),
    .D_N(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__nand3_1 _16024_ (.A(_09093_),
    .B(_09095_),
    .C(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__a21oi_1 _16025_ (.A1(_09095_),
    .A2(_09098_),
    .B1(_09093_),
    .Y(_09100_));
 sky130_fd_sc_hd__a21oi_1 _16026_ (.A1(_09089_),
    .A2(_09099_),
    .B1(_09100_),
    .Y(_09101_));
 sky130_fd_sc_hd__xor2_1 _16027_ (.A(_09083_),
    .B(_09101_),
    .X(_09102_));
 sky130_fd_sc_hd__clkbuf_4 _16028_ (.A(_08449_),
    .X(_09103_));
 sky130_fd_sc_hd__o21a_1 _16029_ (.A1(_09086_),
    .A2(_08517_),
    .B1(_09085_),
    .X(_09104_));
 sky130_fd_sc_hd__or3_1 _16030_ (.A(_09086_),
    .B(_08517_),
    .C(_09085_),
    .X(_09105_));
 sky130_fd_sc_hd__o21a_1 _16031_ (.A1(_09084_),
    .A2(_09104_),
    .B1(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__or3_2 _16032_ (.A(_09103_),
    .B(_08874_),
    .C(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__buf_4 _16033_ (.A(_09103_),
    .X(_09108_));
 sky130_fd_sc_hd__o21ai_1 _16034_ (.A1(_09108_),
    .A2(_08874_),
    .B1(_09106_),
    .Y(_09109_));
 sky130_fd_sc_hd__and2_1 _16035_ (.A(_09107_),
    .B(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__nand2_1 _16036_ (.A(_09102_),
    .B(_09110_),
    .Y(_09111_));
 sky130_fd_sc_hd__o21ai_2 _16037_ (.A1(_09083_),
    .A2(_09101_),
    .B1(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__and2b_1 _16038_ (.A_N(_09082_),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__xnor2_1 _16039_ (.A(_09082_),
    .B(_09112_),
    .Y(_09114_));
 sky130_fd_sc_hd__and2b_1 _16040_ (.A_N(_09107_),
    .B(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__nand2_1 _16041_ (.A(_09075_),
    .B(_09072_),
    .Y(_09116_));
 sky130_fd_sc_hd__nand2_1 _16042_ (.A(_09067_),
    .B(_09073_),
    .Y(_09117_));
 sky130_fd_sc_hd__and2_1 _16043_ (.A(_09074_),
    .B(_09117_),
    .X(_09118_));
 sky130_fd_sc_hd__o211a_1 _16044_ (.A1(_09113_),
    .A2(_09115_),
    .B1(_09116_),
    .C1(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__and3_1 _16045_ (.A(_09039_),
    .B(_09076_),
    .C(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__a21o_1 _16046_ (.A1(_09078_),
    .A2(_09079_),
    .B1(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__a21bo_1 _16047_ (.A1(_09117_),
    .A2(_09113_),
    .B1_N(_09116_),
    .X(_09122_));
 sky130_fd_sc_hd__nand2_1 _16048_ (.A(_09074_),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__or2_1 _16049_ (.A(_09102_),
    .B(_09110_),
    .X(_09124_));
 sky130_fd_sc_hd__nand2_1 _16050_ (.A(_09111_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__and2b_1 _16051_ (.A_N(_09100_),
    .B(_09099_),
    .X(_09126_));
 sky130_fd_sc_hd__xnor2_1 _16052_ (.A(_09089_),
    .B(_09126_),
    .Y(_09127_));
 sky130_fd_sc_hd__a2bb2o_1 _16053_ (.A1_N(_08493_),
    .A2_N(_09096_),
    .B1(_09095_),
    .B2(_09097_),
    .X(_09128_));
 sky130_fd_sc_hd__nand2_1 _16054_ (.A(_09098_),
    .B(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__or2_1 _16055_ (.A(_08517_),
    .B(_09096_),
    .X(_09130_));
 sky130_fd_sc_hd__and2_1 _16056_ (.A(_08490_),
    .B(_08755_),
    .X(_09131_));
 sky130_fd_sc_hd__nand2_1 _16057_ (.A(_09094_),
    .B(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__clkbuf_4 _16058_ (.A(_08490_),
    .X(_09133_));
 sky130_fd_sc_hd__a2bb2o_1 _16059_ (.A1_N(_08724_),
    .A2_N(_08664_),
    .B1(_09133_),
    .B2(_08665_),
    .X(_09134_));
 sky130_fd_sc_hd__nand2_1 _16060_ (.A(_09132_),
    .B(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__o21a_1 _16061_ (.A1(_09130_),
    .A2(_09135_),
    .B1(_09132_),
    .X(_09136_));
 sky130_fd_sc_hd__xor2_1 _16062_ (.A(_09129_),
    .B(_09136_),
    .X(_09137_));
 sky130_fd_sc_hd__clkbuf_4 _16063_ (.A(_08584_),
    .X(_09138_));
 sky130_fd_sc_hd__clkbuf_4 _16064_ (.A(_09086_),
    .X(_09139_));
 sky130_fd_sc_hd__or4_1 _16065_ (.A(_09138_),
    .B(_09139_),
    .C(_08517_),
    .D(_08874_),
    .X(_09140_));
 sky130_fd_sc_hd__o22ai_1 _16066_ (.A1(_09138_),
    .A2(_08517_),
    .B1(_08874_),
    .B2(_09139_),
    .Y(_09141_));
 sky130_fd_sc_hd__and2_1 _16067_ (.A(_09140_),
    .B(_09141_),
    .X(_09142_));
 sky130_fd_sc_hd__nor2_1 _16068_ (.A(_09129_),
    .B(_09136_),
    .Y(_09143_));
 sky130_fd_sc_hd__a21oi_1 _16069_ (.A1(_09137_),
    .A2(_09142_),
    .B1(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__xnor2_1 _16070_ (.A(_09127_),
    .B(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__nor2_1 _16071_ (.A(_09140_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__o21ba_1 _16072_ (.A1(_09127_),
    .A2(_09144_),
    .B1_N(_09146_),
    .X(_09147_));
 sky130_fd_sc_hd__and2_1 _16073_ (.A(_09140_),
    .B(_09145_),
    .X(_09148_));
 sky130_fd_sc_hd__and2_1 _16074_ (.A(_09137_),
    .B(_09142_),
    .X(_09149_));
 sky130_fd_sc_hd__xor2_1 _16075_ (.A(_09130_),
    .B(_09135_),
    .X(_09150_));
 sky130_fd_sc_hd__nor2_1 _16076_ (.A(_08309_),
    .B(_08632_),
    .Y(_09151_));
 sky130_fd_sc_hd__or2_1 _16077_ (.A(_08514_),
    .B(_08626_),
    .X(_09152_));
 sky130_fd_sc_hd__xnor2_1 _16078_ (.A(_09131_),
    .B(_09151_),
    .Y(_09153_));
 sky130_fd_sc_hd__nor2_1 _16079_ (.A(_09152_),
    .B(_09153_),
    .Y(_09154_));
 sky130_fd_sc_hd__a21o_1 _16080_ (.A1(_09131_),
    .A2(_09151_),
    .B1(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__nor2_1 _16081_ (.A(_09150_),
    .B(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__or4b_1 _16082_ (.A(_08325_),
    .B(net7444),
    .C(_09154_),
    .D_N(_09151_),
    .X(_09157_));
 sky130_fd_sc_hd__a21o_1 _16083_ (.A1(_09152_),
    .A2(_09153_),
    .B1(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__o21a_1 _16084_ (.A1(_09138_),
    .A2(_08874_),
    .B1(_09158_),
    .X(_09159_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(_09150_),
    .B(_09155_),
    .Y(_09160_));
 sky130_fd_sc_hd__or3_1 _16086_ (.A(_09138_),
    .B(_08874_),
    .C(_09158_),
    .X(_09161_));
 sky130_fd_sc_hd__o211a_1 _16087_ (.A1(_09156_),
    .A2(_09159_),
    .B1(_09160_),
    .C1(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__nor2_1 _16088_ (.A(_09137_),
    .B(_09142_),
    .Y(_09163_));
 sky130_fd_sc_hd__o32a_1 _16089_ (.A1(_09149_),
    .A2(_09162_),
    .A3(_09163_),
    .B1(_09160_),
    .B2(_09161_),
    .X(_09164_));
 sky130_fd_sc_hd__a2111o_1 _16090_ (.A1(_09125_),
    .A2(_09147_),
    .B1(_09148_),
    .C1(_09164_),
    .D1(_09146_),
    .X(_09165_));
 sky130_fd_sc_hd__o21ai_1 _16091_ (.A1(_09125_),
    .A2(_09147_),
    .B1(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__xnor2_1 _16092_ (.A(_09107_),
    .B(_09114_),
    .Y(_09167_));
 sky130_fd_sc_hd__o2111a_1 _16093_ (.A1(_09118_),
    .A2(_09113_),
    .B1(_09166_),
    .C1(_09167_),
    .D1(_09076_),
    .X(_09168_));
 sky130_fd_sc_hd__and3_1 _16094_ (.A(_09039_),
    .B(_09123_),
    .C(_09168_),
    .X(_09169_));
 sky130_fd_sc_hd__and3_1 _16095_ (.A(_09078_),
    .B(_09079_),
    .C(_09120_),
    .X(_09170_));
 sky130_fd_sc_hd__a21oi_1 _16096_ (.A1(_09121_),
    .A2(_09169_),
    .B1(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__and2_1 _16097_ (.A(_09036_),
    .B(_09078_),
    .X(_09172_));
 sky130_fd_sc_hd__xnor2_1 _16098_ (.A(_08997_),
    .B(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__o22a_2 _16099_ (.A1(_08997_),
    .A2(_09078_),
    .B1(_09171_),
    .B2(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__nor2_1 _16100_ (.A(_09036_),
    .B(_08997_),
    .Y(_09175_));
 sky130_fd_sc_hd__or2_1 _16101_ (.A(_08994_),
    .B(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__xnor2_2 _16102_ (.A(_08995_),
    .B(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__a2bb2o_2 _16103_ (.A1_N(_09174_),
    .A2_N(_09177_),
    .B1(_08995_),
    .B2(_09175_),
    .X(_09178_));
 sky130_fd_sc_hd__nor2_2 _16104_ (.A(_08938_),
    .B(_08996_),
    .Y(_09179_));
 sky130_fd_sc_hd__xnor2_4 _16105_ (.A(_08945_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__a22o_4 _16106_ (.A1(_08945_),
    .A2(_08996_),
    .B1(_09178_),
    .B2(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__a21o_1 _16107_ (.A1(_08938_),
    .A2(_08944_),
    .B1(_08943_),
    .X(_09182_));
 sky130_fd_sc_hd__xnor2_4 _16108_ (.A(_08836_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__a2bb2o_4 _16109_ (.A1_N(_08836_),
    .A2_N(_08946_),
    .B1(_09181_),
    .B2(_09183_),
    .X(_09184_));
 sky130_fd_sc_hd__a21o_1 _16110_ (.A1(_08730_),
    .A2(_08740_),
    .B1(_08738_),
    .X(_09185_));
 sky130_fd_sc_hd__or2b_1 _16111_ (.A(_08572_),
    .B_N(_08533_),
    .X(_09186_));
 sky130_fd_sc_hd__nand2_1 _16112_ (.A(_08698_),
    .B(_08701_),
    .Y(_09187_));
 sky130_fd_sc_hd__or3_1 _16113_ (.A(_09091_),
    .B(_08454_),
    .C(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__a2bb2o_1 _16114_ (.A1_N(_08724_),
    .A2_N(_08331_),
    .B1(_08698_),
    .B2(_09051_),
    .X(_09189_));
 sky130_fd_sc_hd__nand2_1 _16115_ (.A(_09188_),
    .B(_09189_),
    .Y(_09190_));
 sky130_fd_sc_hd__and2b_1 _16116_ (.A_N(_08707_),
    .B(_09133_),
    .X(_09191_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_09190_),
    .B(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__or2_1 _16118_ (.A(_08394_),
    .B(_08484_),
    .X(_09193_));
 sky130_fd_sc_hd__nor2_1 _16119_ (.A(_08529_),
    .B(_08470_),
    .Y(_09194_));
 sky130_fd_sc_hd__xnor2_1 _16120_ (.A(_09193_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__nor2_1 _16121_ (.A(_08411_),
    .B(_08498_),
    .Y(_09196_));
 sky130_fd_sc_hd__xnor2_1 _16122_ (.A(_09195_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__o31a_1 _16123_ (.A1(_08433_),
    .A2(_08498_),
    .A3(_08733_),
    .B1(_08731_),
    .X(_09198_));
 sky130_fd_sc_hd__nor2_1 _16124_ (.A(_09197_),
    .B(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__and2_1 _16125_ (.A(_09197_),
    .B(_09198_),
    .X(_09200_));
 sky130_fd_sc_hd__nor2_1 _16126_ (.A(_09199_),
    .B(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__xnor2_1 _16127_ (.A(_09192_),
    .B(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__a21o_1 _16128_ (.A1(_08570_),
    .A2(_09186_),
    .B1(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__nand3_1 _16129_ (.A(_08570_),
    .B(_09186_),
    .C(_09202_),
    .Y(_09204_));
 sky130_fd_sc_hd__nand2_1 _16130_ (.A(_09203_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__xnor2_1 _16131_ (.A(_09185_),
    .B(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__a21bo_1 _16132_ (.A1(_08566_),
    .A2(_08568_),
    .B1_N(_08563_),
    .X(_09207_));
 sky130_fd_sc_hd__a21bo_1 _16133_ (.A1(_08585_),
    .A2(_08589_),
    .B1_N(_08583_),
    .X(_09208_));
 sky130_fd_sc_hd__or4_1 _16134_ (.A(_08449_),
    .B(_08424_),
    .C(_08550_),
    .D(_08565_),
    .X(_09209_));
 sky130_fd_sc_hd__o22ai_1 _16135_ (.A1(_08449_),
    .A2(_08588_),
    .B1(_08565_),
    .B2(_09064_),
    .Y(_09210_));
 sky130_fd_sc_hd__nand2_1 _16136_ (.A(_09209_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nor2_1 _16137_ (.A(_08564_),
    .B(_08684_),
    .Y(_09212_));
 sky130_fd_sc_hd__xnor2_2 _16138_ (.A(_09211_),
    .B(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__xnor2_2 _16139_ (.A(_09208_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__xnor2_2 _16140_ (.A(_09207_),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__a21oi_4 _16141_ (.A1(_08596_),
    .A2(_08597_),
    .B1(_08598_),
    .Y(_09216_));
 sky130_fd_sc_hd__or4_1 _16142_ (.A(_08559_),
    .B(_08560_),
    .C(_08581_),
    .D(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__o22ai_1 _16143_ (.A1(_09086_),
    .A2(_08582_),
    .B1(_09216_),
    .B2(_08584_),
    .Y(_09218_));
 sky130_fd_sc_hd__nand2_1 _16144_ (.A(_09217_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__nor2_1 _16145_ (.A(_08587_),
    .B(_08574_),
    .Y(_09220_));
 sky130_fd_sc_hd__xnor2_2 _16146_ (.A(_09219_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__a21boi_2 _16147_ (.A1(net3170),
    .A2(_08313_),
    .B1_N(_08630_),
    .Y(_09222_));
 sky130_fd_sc_hd__nor2_1 _16148_ (.A(_08626_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__o21ai_1 _16149_ (.A1(_08615_),
    .A2(_08607_),
    .B1(_08173_),
    .Y(_09224_));
 sky130_fd_sc_hd__or3_1 _16150_ (.A(_08615_),
    .B(_08173_),
    .C(_08607_),
    .X(_09225_));
 sky130_fd_sc_hd__a31o_1 _16151_ (.A1(_08633_),
    .A2(_09224_),
    .A3(_09225_),
    .B1(_08610_),
    .X(_09226_));
 sky130_fd_sc_hd__or4_4 _16152_ (.A(net3722),
    .B(_08328_),
    .C(_08628_),
    .D(_09226_),
    .X(_09227_));
 sky130_fd_sc_hd__nand2_1 _16153_ (.A(_08618_),
    .B(_08665_),
    .Y(_09228_));
 sky130_fd_sc_hd__xor2_2 _16154_ (.A(_09227_),
    .B(_09228_),
    .X(_09229_));
 sky130_fd_sc_hd__xnor2_2 _16155_ (.A(_09223_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_4 _16156_ (.A(_06211_),
    .B(_08618_),
    .Y(_09231_));
 sky130_fd_sc_hd__o32a_1 _16157_ (.A1(_08612_),
    .A2(net7444),
    .A3(_09231_),
    .B1(_08620_),
    .B2(_08603_),
    .X(_09232_));
 sky130_fd_sc_hd__xor2_2 _16158_ (.A(_09230_),
    .B(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__xnor2_2 _16159_ (.A(_09221_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_1 _16160_ (.A(_08621_),
    .B(_08637_),
    .Y(_09235_));
 sky130_fd_sc_hd__a21bo_1 _16161_ (.A1(_08590_),
    .A2(_08638_),
    .B1_N(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__xnor2_2 _16162_ (.A(_09234_),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__xnor2_2 _16163_ (.A(_09215_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__and2b_1 _16164_ (.A_N(_08639_),
    .B(_08653_),
    .X(_09239_));
 sky130_fd_sc_hd__a21oi_1 _16165_ (.A1(_08573_),
    .A2(_08654_),
    .B1(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__xor2_1 _16166_ (.A(_09238_),
    .B(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__xnor2_1 _16167_ (.A(_09206_),
    .B(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__nor2_1 _16168_ (.A(_08655_),
    .B(_08696_),
    .Y(_09243_));
 sky130_fd_sc_hd__a21oi_1 _16169_ (.A1(_08697_),
    .A2(_08745_),
    .B1(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__nor2_1 _16170_ (.A(_09242_),
    .B(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__and2_1 _16171_ (.A(_09242_),
    .B(_09244_),
    .X(_09246_));
 sky130_fd_sc_hd__nor2_1 _16172_ (.A(_09245_),
    .B(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__or2b_1 _16173_ (.A(_08744_),
    .B_N(_08722_),
    .X(_09248_));
 sky130_fd_sc_hd__nand2_4 _16174_ (.A(net6148),
    .B(_08299_),
    .Y(_09249_));
 sky130_fd_sc_hd__or2_2 _16175_ (.A(_08312_),
    .B(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__clkbuf_4 _16176_ (.A(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__or2_1 _16177_ (.A(_08310_),
    .B(_09251_),
    .X(_09252_));
 sky130_fd_sc_hd__nor2_1 _16178_ (.A(_08796_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__o22a_1 _16179_ (.A1(_08310_),
    .A2(_08795_),
    .B1(_09251_),
    .B2(_08326_),
    .X(_09254_));
 sky130_fd_sc_hd__or2_1 _16180_ (.A(_09253_),
    .B(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__a21oi_1 _16181_ (.A1(_08726_),
    .A2(_08728_),
    .B1(_09255_),
    .Y(_09256_));
 sky130_fd_sc_hd__and3_1 _16182_ (.A(_08726_),
    .B(_08728_),
    .C(_09255_),
    .X(_09257_));
 sky130_fd_sc_hd__nor2_1 _16183_ (.A(_09256_),
    .B(_09257_),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_1 _16184_ (.A(_08799_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__or2_1 _16185_ (.A(_08799_),
    .B(_09258_),
    .X(_09260_));
 sky130_fd_sc_hd__nand2_1 _16186_ (.A(_09259_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__a21oi_4 _16187_ (.A1(_08742_),
    .A2(_09248_),
    .B1(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__and3_1 _16188_ (.A(_08742_),
    .B(_09248_),
    .C(_09261_),
    .X(_09263_));
 sky130_fd_sc_hd__nor2_1 _16189_ (.A(_09262_),
    .B(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__xnor2_2 _16190_ (.A(_09247_),
    .B(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__a21oi_2 _16191_ (.A1(_08790_),
    .A2(_08804_),
    .B1(_08788_),
    .Y(_09266_));
 sky130_fd_sc_hd__xor2_2 _16192_ (.A(_09265_),
    .B(_09266_),
    .X(_09267_));
 sky130_fd_sc_hd__xnor2_1 _16193_ (.A(_08802_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__or2b_1 _16194_ (.A(_08805_),
    .B_N(_08834_),
    .X(_09269_));
 sky130_fd_sc_hd__a21boi_2 _16195_ (.A1(_08528_),
    .A2(_08835_),
    .B1_N(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__xor2_1 _16196_ (.A(_09268_),
    .B(_09270_),
    .X(_09271_));
 sky130_fd_sc_hd__and2b_1 _16197_ (.A_N(_08943_),
    .B(_08836_),
    .X(_09272_));
 sky130_fd_sc_hd__nand2_1 _16198_ (.A(_09271_),
    .B(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__or2_1 _16199_ (.A(_09271_),
    .B(_09272_),
    .X(_09274_));
 sky130_fd_sc_hd__and2_4 _16200_ (.A(_09273_),
    .B(_09274_),
    .X(_09275_));
 sky130_fd_sc_hd__xor2_4 _16201_ (.A(_09184_),
    .B(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__mux2_1 _16202_ (.A0(net2942),
    .A1(net7732),
    .S(net4087),
    .X(_09277_));
 sky130_fd_sc_hd__nand2_1 _16203_ (.A(_09276_),
    .B(net2943),
    .Y(_09278_));
 sky130_fd_sc_hd__or2_1 _16204_ (.A(_09276_),
    .B(net2943),
    .X(_09279_));
 sky130_fd_sc_hd__and2_1 _16205_ (.A(_09278_),
    .B(_09279_),
    .X(_09280_));
 sky130_fd_sc_hd__xor2_4 _16206_ (.A(_09181_),
    .B(_09183_),
    .X(_09281_));
 sky130_fd_sc_hd__mux2_2 _16207_ (.A0(net4893),
    .A1(net5463),
    .S(net4088),
    .X(_09282_));
 sky130_fd_sc_hd__nor2_1 _16208_ (.A(_09281_),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__xor2_4 _16209_ (.A(_09178_),
    .B(_09180_),
    .X(_09284_));
 sky130_fd_sc_hd__mux2_1 _16210_ (.A0(net3024),
    .A1(net4306),
    .S(net4087),
    .X(_09285_));
 sky130_fd_sc_hd__xor2_4 _16211_ (.A(_09174_),
    .B(_09177_),
    .X(_09286_));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(net4355),
    .A1(net7370),
    .S(_08293_),
    .X(_09287_));
 sky130_fd_sc_hd__o211a_1 _16213_ (.A1(_09284_),
    .A2(net3025),
    .B1(_09286_),
    .C1(net7371),
    .X(_09288_));
 sky130_fd_sc_hd__a21oi_1 _16214_ (.A1(_09284_),
    .A2(net3025),
    .B1(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_1 _16215_ (.A(_09281_),
    .B(net8010),
    .Y(_09290_));
 sky130_fd_sc_hd__o21ai_1 _16216_ (.A1(_09283_),
    .A2(_09289_),
    .B1(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__nand2_1 _16217_ (.A(_09280_),
    .B(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__or2_1 _16218_ (.A(_09280_),
    .B(_09291_),
    .X(_09293_));
 sky130_fd_sc_hd__buf_4 _16219_ (.A(net7405),
    .X(_09294_));
 sky130_fd_sc_hd__inv_2 _16220_ (.A(_09294_),
    .Y(_09295_));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(_09295_),
    .A1(_06396_),
    .S(net4088),
    .X(_09296_));
 sky130_fd_sc_hd__buf_1 _16222_ (.A(net7406),
    .X(_09297_));
 sky130_fd_sc_hd__a21oi_1 _16223_ (.A1(_09292_),
    .A2(_09293_),
    .B1(net7407),
    .Y(_09298_));
 sky130_fd_sc_hd__a31o_1 _16224_ (.A1(_09292_),
    .A2(_09293_),
    .A3(net7407),
    .B1(_08633_),
    .X(_09299_));
 sky130_fd_sc_hd__o221a_1 _16225_ (.A1(net4376),
    .A2(_08296_),
    .B1(_09298_),
    .B2(_09299_),
    .C1(_08239_),
    .X(_00466_));
 sky130_fd_sc_hd__a21boi_2 _16226_ (.A1(_09184_),
    .A2(_09275_),
    .B1_N(_09273_),
    .Y(_09300_));
 sky130_fd_sc_hd__or2_4 _16227_ (.A(_09268_),
    .B(_09270_),
    .X(_09301_));
 sky130_fd_sc_hd__or2b_1 _16228_ (.A(_09205_),
    .B_N(_09185_),
    .X(_09302_));
 sky130_fd_sc_hd__or2b_1 _16229_ (.A(_09190_),
    .B_N(_09191_),
    .X(_09303_));
 sky130_fd_sc_hd__clkbuf_4 _16230_ (.A(_08328_),
    .X(_09304_));
 sky130_fd_sc_hd__clkbuf_4 _16231_ (.A(_09304_),
    .X(_09305_));
 sky130_fd_sc_hd__nor2_2 _16232_ (.A(_09305_),
    .B(_08793_),
    .Y(_09306_));
 sky130_fd_sc_hd__and3b_1 _16233_ (.A_N(_09252_),
    .B(_09133_),
    .C(_09306_),
    .X(_09307_));
 sky130_fd_sc_hd__a21boi_1 _16234_ (.A1(_09133_),
    .A2(_09306_),
    .B1_N(_09252_),
    .Y(_09308_));
 sky130_fd_sc_hd__nor2_1 _16235_ (.A(_09307_),
    .B(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand2_2 _16236_ (.A(net6150),
    .B(_08314_),
    .Y(_09310_));
 sky130_fd_sc_hd__or2_2 _16237_ (.A(_08313_),
    .B(_09310_),
    .X(_09311_));
 sky130_fd_sc_hd__clkbuf_4 _16238_ (.A(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__nor2_1 _16239_ (.A(_08325_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__xnor2_1 _16240_ (.A(_09309_),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__and3_1 _16241_ (.A(_09188_),
    .B(_09303_),
    .C(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__a21o_1 _16242_ (.A1(_09188_),
    .A2(_09303_),
    .B1(_09314_),
    .X(_09316_));
 sky130_fd_sc_hd__or2b_1 _16243_ (.A(_09315_),
    .B_N(_09316_),
    .X(_09317_));
 sky130_fd_sc_hd__nor2_1 _16244_ (.A(_09253_),
    .B(_09256_),
    .Y(_09318_));
 sky130_fd_sc_hd__xnor2_1 _16245_ (.A(_09317_),
    .B(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__a21oi_1 _16246_ (.A1(_09203_),
    .A2(_09302_),
    .B1(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__and3_1 _16247_ (.A(_09203_),
    .B(_09302_),
    .C(_09319_),
    .X(_09321_));
 sky130_fd_sc_hd__nor2_1 _16248_ (.A(_09320_),
    .B(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__xnor2_1 _16249_ (.A(_09259_),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__a21o_1 _16250_ (.A1(_09192_),
    .A2(_09201_),
    .B1(_09199_),
    .X(_09324_));
 sky130_fd_sc_hd__nand2_1 _16251_ (.A(_09208_),
    .B(_09213_),
    .Y(_09325_));
 sky130_fd_sc_hd__or2b_1 _16252_ (.A(_09214_),
    .B_N(_09207_),
    .X(_09326_));
 sky130_fd_sc_hd__or3_1 _16253_ (.A(_08409_),
    .B(_09091_),
    .C(_09187_),
    .X(_09327_));
 sky130_fd_sc_hd__buf_2 _16254_ (.A(_08409_),
    .X(_09328_));
 sky130_fd_sc_hd__a2bb2o_1 _16255_ (.A1_N(_08316_),
    .A2_N(_09328_),
    .B1(_09051_),
    .B2(_08701_),
    .X(_09329_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(_09327_),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__or3_1 _16257_ (.A(_08724_),
    .B(_08707_),
    .C(_09330_),
    .X(_09331_));
 sky130_fd_sc_hd__o21ai_1 _16258_ (.A1(_08724_),
    .A2(_08708_),
    .B1(_09330_),
    .Y(_09332_));
 sky130_fd_sc_hd__and2_1 _16259_ (.A(_09331_),
    .B(_09332_),
    .X(_09333_));
 sky130_fd_sc_hd__or4_1 _16260_ (.A(_08564_),
    .B(_08529_),
    .C(_08471_),
    .D(_08484_),
    .X(_09334_));
 sky130_fd_sc_hd__o22ai_1 _16261_ (.A1(_08564_),
    .A2(_08471_),
    .B1(_08516_),
    .B2(_08529_),
    .Y(_09335_));
 sky130_fd_sc_hd__nand2_1 _16262_ (.A(_09334_),
    .B(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__or2_1 _16263_ (.A(_08394_),
    .B(_08498_),
    .X(_09337_));
 sky130_fd_sc_hd__xnor2_1 _16264_ (.A(_09336_),
    .B(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__or3_1 _16265_ (.A(_08529_),
    .B(_08471_),
    .C(_09193_),
    .X(_09339_));
 sky130_fd_sc_hd__a21boi_1 _16266_ (.A1(_09195_),
    .A2(_09196_),
    .B1_N(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__nor2_1 _16267_ (.A(_09338_),
    .B(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__and2_1 _16268_ (.A(_09338_),
    .B(_09340_),
    .X(_09342_));
 sky130_fd_sc_hd__nor2_1 _16269_ (.A(_09341_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__xnor2_1 _16270_ (.A(_09333_),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__a21o_1 _16271_ (.A1(_09325_),
    .A2(_09326_),
    .B1(_09344_),
    .X(_09345_));
 sky130_fd_sc_hd__nand3_1 _16272_ (.A(_09325_),
    .B(_09326_),
    .C(_09344_),
    .Y(_09346_));
 sky130_fd_sc_hd__nand2_1 _16273_ (.A(_09345_),
    .B(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__xnor2_1 _16274_ (.A(_09324_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__a21bo_1 _16275_ (.A1(_09210_),
    .A2(_09212_),
    .B1_N(_09209_),
    .X(_09349_));
 sky130_fd_sc_hd__a21bo_1 _16276_ (.A1(_09218_),
    .A2(_09220_),
    .B1_N(_09217_),
    .X(_09350_));
 sky130_fd_sc_hd__or4_1 _16277_ (.A(_08449_),
    .B(_09064_),
    .C(_08574_),
    .D(_08588_),
    .X(_09351_));
 sky130_fd_sc_hd__a2bb2o_1 _16278_ (.A1_N(_08588_),
    .A2_N(_09064_),
    .B1(_08969_),
    .B2(_08642_),
    .X(_09352_));
 sky130_fd_sc_hd__nand2_1 _16279_ (.A(_09351_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__nor2_1 _16280_ (.A(_08684_),
    .B(_08565_),
    .Y(_09354_));
 sky130_fd_sc_hd__xnor2_2 _16281_ (.A(_09353_),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__xnor2_2 _16282_ (.A(_09350_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__xnor2_2 _16283_ (.A(_09349_),
    .B(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__nor2_1 _16284_ (.A(_08587_),
    .B(_08582_),
    .Y(_09358_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(_08560_),
    .B(_09216_),
    .Y(_09359_));
 sky130_fd_sc_hd__nor2_1 _16286_ (.A(_08559_),
    .B(_09222_),
    .Y(_09360_));
 sky130_fd_sc_hd__xor2_2 _16287_ (.A(_09359_),
    .B(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__xor2_2 _16288_ (.A(_09358_),
    .B(_09361_),
    .X(_09362_));
 sky130_fd_sc_hd__nor2_1 _16289_ (.A(net3273),
    .B(_06211_),
    .Y(_09363_));
 sky130_fd_sc_hd__a21oi_2 _16290_ (.A1(_06211_),
    .A2(_08618_),
    .B1(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__or2_1 _16291_ (.A(_08626_),
    .B(_09364_),
    .X(_09365_));
 sky130_fd_sc_hd__nor4_4 _16292_ (.A(_08615_),
    .B(_08173_),
    .C(_08177_),
    .D(_08607_),
    .Y(_09366_));
 sky130_fd_sc_hd__o31a_1 _16293_ (.A1(_08615_),
    .A2(_08173_),
    .A3(_08607_),
    .B1(_08177_),
    .X(_09367_));
 sky130_fd_sc_hd__o31ai_4 _16294_ (.A1(_08296_),
    .A2(_09366_),
    .A3(_09367_),
    .B1(_08609_),
    .Y(_09368_));
 sky130_fd_sc_hd__or4_1 _16295_ (.A(net3722),
    .B(_08328_),
    .C(_08628_),
    .D(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__or4_1 _16296_ (.A(net3539),
    .B(_08328_),
    .C(_08628_),
    .D(_09226_),
    .X(_09370_));
 sky130_fd_sc_hd__or4_2 _16297_ (.A(net3539),
    .B(_08313_),
    .C(_08628_),
    .D(_09368_),
    .X(_09371_));
 sky130_fd_sc_hd__o2bb2a_1 _16298_ (.A1_N(_09369_),
    .A2_N(_09370_),
    .B1(_09227_),
    .B2(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__xor2_1 _16299_ (.A(_09365_),
    .B(_09372_),
    .X(_09373_));
 sky130_fd_sc_hd__nand2_1 _16300_ (.A(net3103),
    .B(_08628_),
    .Y(_09374_));
 sky130_fd_sc_hd__a21o_2 _16301_ (.A1(_09374_),
    .A2(_09226_),
    .B1(_08328_),
    .X(_09375_));
 sky130_fd_sc_hd__nor2_1 _16302_ (.A(net7444),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__a32o_1 _16303_ (.A1(_08618_),
    .A2(_08665_),
    .A3(_09376_),
    .B1(_09229_),
    .B2(_09223_),
    .X(_09377_));
 sky130_fd_sc_hd__xnor2_2 _16304_ (.A(_09373_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__xnor2_2 _16305_ (.A(_09362_),
    .B(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__nor2_1 _16306_ (.A(_09230_),
    .B(_09232_),
    .Y(_09380_));
 sky130_fd_sc_hd__a21oi_2 _16307_ (.A1(_09221_),
    .A2(_09233_),
    .B1(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__xor2_2 _16308_ (.A(_09379_),
    .B(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__xnor2_2 _16309_ (.A(_09357_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__and2b_1 _16310_ (.A_N(_09234_),
    .B(_09236_),
    .X(_09384_));
 sky130_fd_sc_hd__a21oi_2 _16311_ (.A1(_09215_),
    .A2(_09237_),
    .B1(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__nor2_1 _16312_ (.A(_09383_),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand2_1 _16313_ (.A(_09383_),
    .B(_09385_),
    .Y(_09387_));
 sky130_fd_sc_hd__and2b_1 _16314_ (.A_N(_09386_),
    .B(_09387_),
    .X(_09388_));
 sky130_fd_sc_hd__xnor2_1 _16315_ (.A(_09348_),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__nor2_1 _16316_ (.A(_09238_),
    .B(_09240_),
    .Y(_09390_));
 sky130_fd_sc_hd__a21oi_1 _16317_ (.A1(_09206_),
    .A2(_09241_),
    .B1(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__xor2_1 _16318_ (.A(_09389_),
    .B(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__xnor2_1 _16319_ (.A(_09323_),
    .B(_09392_),
    .Y(_09393_));
 sky130_fd_sc_hd__a21oi_1 _16320_ (.A1(_09247_),
    .A2(_09264_),
    .B1(_09245_),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_1 _16321_ (.A(_09393_),
    .B(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(_09393_),
    .B(_09394_),
    .Y(_09396_));
 sky130_fd_sc_hd__and2b_1 _16323_ (.A_N(_09395_),
    .B(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__xnor2_4 _16324_ (.A(_09262_),
    .B(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__nor2_1 _16325_ (.A(_09265_),
    .B(_09266_),
    .Y(_09399_));
 sky130_fd_sc_hd__a21oi_2 _16326_ (.A1(_08802_),
    .A2(_09267_),
    .B1(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__xnor2_4 _16327_ (.A(_09398_),
    .B(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__xor2_4 _16328_ (.A(_09301_),
    .B(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__xnor2_4 _16329_ (.A(_09300_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__mux2_1 _16330_ (.A0(net7380),
    .A1(net2935),
    .S(_08293_),
    .X(_09404_));
 sky130_fd_sc_hd__and2_1 _16331_ (.A(_09403_),
    .B(net7381),
    .X(_09405_));
 sky130_fd_sc_hd__nor2_1 _16332_ (.A(_09403_),
    .B(net7381),
    .Y(_09406_));
 sky130_fd_sc_hd__or2_1 _16333_ (.A(_09405_),
    .B(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__a21oi_1 _16334_ (.A1(_09278_),
    .A2(_09292_),
    .B1(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__and3_1 _16335_ (.A(_09278_),
    .B(_09292_),
    .C(_09407_),
    .X(_09409_));
 sky130_fd_sc_hd__nor2_1 _16336_ (.A(_09408_),
    .B(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__nor2_1 _16337_ (.A(net7407),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__a21o_1 _16338_ (.A1(net7407),
    .A2(_09410_),
    .B1(_08633_),
    .X(_09412_));
 sky130_fd_sc_hd__o221a_1 _16339_ (.A1(net4351),
    .A2(_08296_),
    .B1(_09411_),
    .B2(_09412_),
    .C1(_08239_),
    .X(_00467_));
 sky130_fd_sc_hd__nor2_1 _16340_ (.A(_09398_),
    .B(_09400_),
    .Y(_09413_));
 sky130_fd_sc_hd__a31o_1 _16341_ (.A1(_08799_),
    .A2(_09258_),
    .A3(_09322_),
    .B1(_09320_),
    .X(_09414_));
 sky130_fd_sc_hd__or2_1 _16342_ (.A(_09389_),
    .B(_09391_),
    .X(_09415_));
 sky130_fd_sc_hd__nand2_1 _16343_ (.A(_09323_),
    .B(_09392_),
    .Y(_09416_));
 sky130_fd_sc_hd__or2b_1 _16344_ (.A(_09347_),
    .B_N(_09324_),
    .X(_09417_));
 sky130_fd_sc_hd__nand2_2 _16345_ (.A(net7951),
    .B(_08314_),
    .Y(_09418_));
 sky130_fd_sc_hd__or2_1 _16346_ (.A(_09305_),
    .B(_09418_),
    .X(_09419_));
 sky130_fd_sc_hd__clkbuf_4 _16347_ (.A(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__or2_2 _16348_ (.A(_08326_),
    .B(_09420_),
    .X(_09421_));
 sky130_fd_sc_hd__a21o_1 _16349_ (.A1(_09309_),
    .A2(_09313_),
    .B1(_09307_),
    .X(_09422_));
 sky130_fd_sc_hd__inv_2 _16350_ (.A(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__nand2_1 _16351_ (.A(_09327_),
    .B(_09331_),
    .Y(_09424_));
 sky130_fd_sc_hd__nor2_1 _16352_ (.A(_08454_),
    .B(_08795_),
    .Y(_09425_));
 sky130_fd_sc_hd__and2b_1 _16353_ (.A_N(_09250_),
    .B(_08490_),
    .X(_09426_));
 sky130_fd_sc_hd__or2_1 _16354_ (.A(_09425_),
    .B(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__nand2_1 _16355_ (.A(_09425_),
    .B(_09426_),
    .Y(_09428_));
 sky130_fd_sc_hd__and2_1 _16356_ (.A(_09427_),
    .B(_09428_),
    .X(_09429_));
 sky130_fd_sc_hd__nor2_1 _16357_ (.A(_08310_),
    .B(_09311_),
    .Y(_09430_));
 sky130_fd_sc_hd__xnor2_1 _16358_ (.A(_09429_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__xor2_1 _16359_ (.A(_09424_),
    .B(_09431_),
    .X(_09432_));
 sky130_fd_sc_hd__xnor2_1 _16360_ (.A(_09423_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__inv_2 _16361_ (.A(_09253_),
    .Y(_09434_));
 sky130_fd_sc_hd__a21o_1 _16362_ (.A1(_09434_),
    .A2(_09316_),
    .B1(_09315_),
    .X(_09435_));
 sky130_fd_sc_hd__xor2_1 _16363_ (.A(_09433_),
    .B(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__xor2_1 _16364_ (.A(_09421_),
    .B(_09436_),
    .X(_09437_));
 sky130_fd_sc_hd__a21oi_1 _16365_ (.A1(_09345_),
    .A2(_09417_),
    .B1(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__nand3_1 _16366_ (.A(_09345_),
    .B(_09417_),
    .C(_09437_),
    .Y(_09439_));
 sky130_fd_sc_hd__or2b_1 _16367_ (.A(_09438_),
    .B_N(_09439_),
    .X(_09440_));
 sky130_fd_sc_hd__and3b_1 _16368_ (.A_N(_09315_),
    .B(_09316_),
    .C(_09256_),
    .X(_09441_));
 sky130_fd_sc_hd__xnor2_1 _16369_ (.A(_09440_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__a21o_1 _16370_ (.A1(_09333_),
    .A2(_09343_),
    .B1(_09341_),
    .X(_09443_));
 sky130_fd_sc_hd__or2b_1 _16371_ (.A(_09356_),
    .B_N(_09349_),
    .X(_09444_));
 sky130_fd_sc_hd__a21bo_1 _16372_ (.A1(_09350_),
    .A2(_09355_),
    .B1_N(_09444_),
    .X(_09445_));
 sky130_fd_sc_hd__or3b_1 _16373_ (.A(_09187_),
    .B(_09328_),
    .C_N(_08962_),
    .X(_09446_));
 sky130_fd_sc_hd__buf_2 _16374_ (.A(_08962_),
    .X(_09447_));
 sky130_fd_sc_hd__a2bb2o_1 _16375_ (.A1_N(_09328_),
    .A2_N(_08331_),
    .B1(_08698_),
    .B2(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__nand2_1 _16376_ (.A(_09446_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nor2_1 _16377_ (.A(_09091_),
    .B(_08707_),
    .Y(_09450_));
 sky130_fd_sc_hd__xnor2_2 _16378_ (.A(_09449_),
    .B(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__or4_1 _16379_ (.A(_08564_),
    .B(_08471_),
    .C(_08516_),
    .D(_08565_),
    .X(_09452_));
 sky130_fd_sc_hd__o22ai_1 _16380_ (.A1(_08564_),
    .A2(_08873_),
    .B1(_08565_),
    .B2(_08471_),
    .Y(_09453_));
 sky130_fd_sc_hd__and2_1 _16381_ (.A(_09452_),
    .B(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__nor2_1 _16382_ (.A(_08529_),
    .B(_08498_),
    .Y(_09455_));
 sky130_fd_sc_hd__xnor2_1 _16383_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__o31a_1 _16384_ (.A1(_08394_),
    .A2(_08717_),
    .A3(_09336_),
    .B1(_09334_),
    .X(_09457_));
 sky130_fd_sc_hd__nor2_1 _16385_ (.A(_09456_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__and2_1 _16386_ (.A(_09456_),
    .B(_09457_),
    .X(_09459_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(_09458_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__xor2_2 _16388_ (.A(_09451_),
    .B(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__xnor2_1 _16389_ (.A(_09445_),
    .B(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__xnor2_1 _16390_ (.A(_09443_),
    .B(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__a21bo_1 _16391_ (.A1(_09352_),
    .A2(_09354_),
    .B1_N(_09351_),
    .X(_09464_));
 sky130_fd_sc_hd__nand2_1 _16392_ (.A(_09359_),
    .B(_09360_),
    .Y(_09465_));
 sky130_fd_sc_hd__a21bo_1 _16393_ (.A1(_09358_),
    .A2(_09361_),
    .B1_N(_09465_),
    .X(_09466_));
 sky130_fd_sc_hd__or2_1 _16394_ (.A(_08424_),
    .B(_08574_),
    .X(_09467_));
 sky130_fd_sc_hd__or2_1 _16395_ (.A(_08449_),
    .B(_08582_),
    .X(_09468_));
 sky130_fd_sc_hd__xnor2_1 _16396_ (.A(_09467_),
    .B(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__nor2_1 _16397_ (.A(_08684_),
    .B(_08588_),
    .Y(_09470_));
 sky130_fd_sc_hd__xnor2_1 _16398_ (.A(_09469_),
    .B(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__and2_1 _16399_ (.A(_09466_),
    .B(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__or2_1 _16400_ (.A(_09466_),
    .B(_09471_),
    .X(_09473_));
 sky130_fd_sc_hd__or2b_1 _16401_ (.A(_09472_),
    .B_N(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__xnor2_2 _16402_ (.A(_09464_),
    .B(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__nor2_1 _16403_ (.A(_08587_),
    .B(_09216_),
    .Y(_09476_));
 sky130_fd_sc_hd__clkbuf_4 _16404_ (.A(_09222_),
    .X(_09477_));
 sky130_fd_sc_hd__nor2_1 _16405_ (.A(_09086_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__nor2_1 _16406_ (.A(_08584_),
    .B(_09364_),
    .Y(_09479_));
 sky130_fd_sc_hd__xor2_2 _16407_ (.A(_09478_),
    .B(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__xor2_2 _16408_ (.A(_09476_),
    .B(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__nand2_1 _16409_ (.A(net3537),
    .B(_08313_),
    .Y(_09482_));
 sky130_fd_sc_hd__and2_1 _16410_ (.A(_09375_),
    .B(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__clkbuf_4 _16411_ (.A(_09483_),
    .X(_09484_));
 sky130_fd_sc_hd__nor2_1 _16412_ (.A(_09096_),
    .B(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__clkbuf_4 _16413_ (.A(_08628_),
    .X(_09486_));
 sky130_fd_sc_hd__or2_1 _16414_ (.A(_08180_),
    .B(net77),
    .X(_09487_));
 sky130_fd_sc_hd__nand2_1 _16415_ (.A(_08180_),
    .B(net77),
    .Y(_09488_));
 sky130_fd_sc_hd__a31o_2 _16416_ (.A1(_08633_),
    .A2(_09487_),
    .A3(_09488_),
    .B1(_08610_),
    .X(_09489_));
 sky130_fd_sc_hd__or4_2 _16417_ (.A(net3722),
    .B(_08313_),
    .C(_09486_),
    .D(_09489_),
    .X(_09490_));
 sky130_fd_sc_hd__xor2_2 _16418_ (.A(_09371_),
    .B(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__xor2_2 _16419_ (.A(_09485_),
    .B(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__nor2_1 _16420_ (.A(_09227_),
    .B(_09371_),
    .Y(_09493_));
 sky130_fd_sc_hd__and2_1 _16421_ (.A(_09369_),
    .B(_09370_),
    .X(_09494_));
 sky130_fd_sc_hd__or3_1 _16422_ (.A(_09365_),
    .B(_09493_),
    .C(_09494_),
    .X(_09495_));
 sky130_fd_sc_hd__and2b_1 _16423_ (.A_N(_09493_),
    .B(_09495_),
    .X(_09496_));
 sky130_fd_sc_hd__xnor2_2 _16424_ (.A(_09492_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__xnor2_2 _16425_ (.A(_09481_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__o21ai_1 _16426_ (.A1(_09493_),
    .A2(_09494_),
    .B1(_09365_),
    .Y(_09499_));
 sky130_fd_sc_hd__a32o_1 _16427_ (.A1(_09495_),
    .A2(_09499_),
    .A3(_09377_),
    .B1(_09378_),
    .B2(_09362_),
    .X(_09500_));
 sky130_fd_sc_hd__xnor2_2 _16428_ (.A(_09498_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__xnor2_2 _16429_ (.A(_09475_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__nor2_1 _16430_ (.A(_09379_),
    .B(_09381_),
    .Y(_09503_));
 sky130_fd_sc_hd__a21oi_2 _16431_ (.A1(_09357_),
    .A2(_09382_),
    .B1(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__xor2_2 _16432_ (.A(_09502_),
    .B(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__xnor2_1 _16433_ (.A(_09463_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__a21oi_1 _16434_ (.A1(_09348_),
    .A2(_09387_),
    .B1(_09386_),
    .Y(_09507_));
 sky130_fd_sc_hd__xor2_1 _16435_ (.A(_09506_),
    .B(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__xnor2_1 _16436_ (.A(_09442_),
    .B(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__a21oi_2 _16437_ (.A1(_09415_),
    .A2(_09416_),
    .B1(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__and3_1 _16438_ (.A(_09415_),
    .B(_09416_),
    .C(_09509_),
    .X(_09511_));
 sky130_fd_sc_hd__nor2_2 _16439_ (.A(_09510_),
    .B(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__xnor2_1 _16440_ (.A(_09414_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__a21oi_1 _16441_ (.A1(_09262_),
    .A2(_09396_),
    .B1(_09395_),
    .Y(_09514_));
 sky130_fd_sc_hd__xor2_1 _16442_ (.A(_09513_),
    .B(_09514_),
    .X(_09515_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(_09413_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__or2_1 _16444_ (.A(_09413_),
    .B(_09515_),
    .X(_09517_));
 sky130_fd_sc_hd__nand2_2 _16445_ (.A(_09516_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__a21oi_1 _16446_ (.A1(_09301_),
    .A2(_09273_),
    .B1(_09401_),
    .Y(_09519_));
 sky130_fd_sc_hd__a31oi_4 _16447_ (.A1(_09184_),
    .A2(_09275_),
    .A3(_09402_),
    .B1(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__xor2_4 _16448_ (.A(_09518_),
    .B(_09520_),
    .X(_09521_));
 sky130_fd_sc_hd__mux2_1 _16449_ (.A0(net3003),
    .A1(net7428),
    .S(_08293_),
    .X(_09522_));
 sky130_fd_sc_hd__xor2_1 _16450_ (.A(_09521_),
    .B(net3004),
    .X(_09523_));
 sky130_fd_sc_hd__o21a_1 _16451_ (.A1(_09405_),
    .A2(_09408_),
    .B1(_09523_),
    .X(_09524_));
 sky130_fd_sc_hd__nor3_1 _16452_ (.A(_09405_),
    .B(_09408_),
    .C(_09523_),
    .Y(_09525_));
 sky130_fd_sc_hd__nor2_1 _16453_ (.A(_09524_),
    .B(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__nor2_1 _16454_ (.A(net7407),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__a21o_1 _16455_ (.A1(net7407),
    .A2(_09526_),
    .B1(_08633_),
    .X(_09528_));
 sky130_fd_sc_hd__o221a_1 _16456_ (.A1(net4313),
    .A2(_08296_),
    .B1(_09527_),
    .B2(_09528_),
    .C1(_08239_),
    .X(_00468_));
 sky130_fd_sc_hd__o21a_1 _16457_ (.A1(_09518_),
    .A2(_09520_),
    .B1(_09516_),
    .X(_09529_));
 sky130_fd_sc_hd__or2_2 _16458_ (.A(_09513_),
    .B(_09514_),
    .X(_09530_));
 sky130_fd_sc_hd__a21o_2 _16459_ (.A1(_09439_),
    .A2(_09441_),
    .B1(_09438_),
    .X(_09531_));
 sky130_fd_sc_hd__or2b_1 _16460_ (.A(_09421_),
    .B_N(_09436_),
    .X(_09532_));
 sky130_fd_sc_hd__o21ai_1 _16461_ (.A1(_09433_),
    .A2(_09435_),
    .B1(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__or2b_1 _16462_ (.A(_09462_),
    .B_N(_09443_),
    .X(_09534_));
 sky130_fd_sc_hd__a21bo_1 _16463_ (.A1(_09445_),
    .A2(_09461_),
    .B1_N(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__nand2_2 _16464_ (.A(net7442),
    .B(_08314_),
    .Y(_09536_));
 sky130_fd_sc_hd__or2_2 _16465_ (.A(_09304_),
    .B(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__clkbuf_4 _16466_ (.A(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__o22a_1 _16467_ (.A1(_08310_),
    .A2(_09420_),
    .B1(_09538_),
    .B2(_08326_),
    .X(_09539_));
 sky130_fd_sc_hd__or2_1 _16468_ (.A(_08310_),
    .B(_09537_),
    .X(_09540_));
 sky130_fd_sc_hd__nor2_1 _16469_ (.A(_09421_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__or2_1 _16470_ (.A(_09539_),
    .B(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__a21bo_1 _16471_ (.A1(_09429_),
    .A2(_09430_),
    .B1_N(_09428_),
    .X(_09543_));
 sky130_fd_sc_hd__a21bo_1 _16472_ (.A1(_09448_),
    .A2(_09450_),
    .B1_N(_09446_),
    .X(_09544_));
 sky130_fd_sc_hd__nor2_1 _16473_ (.A(_09091_),
    .B(_08795_),
    .Y(_09545_));
 sky130_fd_sc_hd__nor2_1 _16474_ (.A(_08724_),
    .B(_09251_),
    .Y(_09546_));
 sky130_fd_sc_hd__nor2_1 _16475_ (.A(_09091_),
    .B(_09251_),
    .Y(_09547_));
 sky130_fd_sc_hd__nand2_1 _16476_ (.A(_09425_),
    .B(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__o21a_1 _16477_ (.A1(_09545_),
    .A2(_09546_),
    .B1(_09548_),
    .X(_09549_));
 sky130_fd_sc_hd__and2b_1 _16478_ (.A_N(_09311_),
    .B(_09133_),
    .X(_09550_));
 sky130_fd_sc_hd__xnor2_2 _16479_ (.A(_09549_),
    .B(_09550_),
    .Y(_09551_));
 sky130_fd_sc_hd__xnor2_2 _16480_ (.A(_09544_),
    .B(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__xnor2_2 _16481_ (.A(_09543_),
    .B(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__a21o_1 _16482_ (.A1(_09327_),
    .A2(_09331_),
    .B1(_09431_),
    .X(_09554_));
 sky130_fd_sc_hd__o21a_1 _16483_ (.A1(_09423_),
    .A2(_09432_),
    .B1(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__xor2_1 _16484_ (.A(_09553_),
    .B(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__xnor2_1 _16485_ (.A(_09542_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__xnor2_1 _16486_ (.A(_09535_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__xnor2_1 _16487_ (.A(_09533_),
    .B(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__a21o_1 _16488_ (.A1(_09451_),
    .A2(_09460_),
    .B1(_09458_),
    .X(_09560_));
 sky130_fd_sc_hd__a21o_1 _16489_ (.A1(_09464_),
    .A2(_09473_),
    .B1(_09472_),
    .X(_09561_));
 sky130_fd_sc_hd__clkbuf_4 _16490_ (.A(_08372_),
    .X(_09562_));
 sky130_fd_sc_hd__nor2_1 _16491_ (.A(_08316_),
    .B(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__a21o_1 _16492_ (.A1(_08701_),
    .A2(_08962_),
    .B1(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__and4b_1 _16493_ (.A_N(_09562_),
    .B(_08962_),
    .C(_08698_),
    .D(_08701_),
    .X(_09565_));
 sky130_fd_sc_hd__inv_2 _16494_ (.A(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand2_1 _16495_ (.A(_09564_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nor2_1 _16496_ (.A(_09328_),
    .B(_08707_),
    .Y(_09568_));
 sky130_fd_sc_hd__xnor2_2 _16497_ (.A(_09567_),
    .B(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__or4_1 _16498_ (.A(_08470_),
    .B(_08484_),
    .C(_08550_),
    .D(_08565_),
    .X(_09570_));
 sky130_fd_sc_hd__o22ai_1 _16499_ (.A1(_08471_),
    .A2(_08588_),
    .B1(_08565_),
    .B2(_08516_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand2_1 _16500_ (.A(_09570_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__or2_1 _16501_ (.A(_08564_),
    .B(_08497_),
    .X(_09573_));
 sky130_fd_sc_hd__xnor2_1 _16502_ (.A(_09572_),
    .B(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__a21boi_1 _16503_ (.A1(_09453_),
    .A2(_09455_),
    .B1_N(_09452_),
    .Y(_09575_));
 sky130_fd_sc_hd__nor2_1 _16504_ (.A(_09574_),
    .B(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__and2_1 _16505_ (.A(_09574_),
    .B(_09575_),
    .X(_09577_));
 sky130_fd_sc_hd__nor2_1 _16506_ (.A(_09576_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__xor2_2 _16507_ (.A(_09569_),
    .B(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__xnor2_2 _16508_ (.A(_09561_),
    .B(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__xnor2_2 _16509_ (.A(_09560_),
    .B(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__clkbuf_4 _16510_ (.A(_08684_),
    .X(_09582_));
 sky130_fd_sc_hd__o32a_1 _16511_ (.A1(_09582_),
    .A2(_08588_),
    .A3(_09469_),
    .B1(_09468_),
    .B2(_09467_),
    .X(_09583_));
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(_09478_),
    .B(_09479_),
    .Y(_09584_));
 sky130_fd_sc_hd__a21bo_1 _16513_ (.A1(_09476_),
    .A2(_09480_),
    .B1_N(_09584_),
    .X(_09585_));
 sky130_fd_sc_hd__nor2_1 _16514_ (.A(_09064_),
    .B(_08582_),
    .Y(_09586_));
 sky130_fd_sc_hd__nor2_1 _16515_ (.A(_09103_),
    .B(_09216_),
    .Y(_09587_));
 sky130_fd_sc_hd__xnor2_1 _16516_ (.A(_09586_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__or2_1 _16517_ (.A(_08684_),
    .B(_08574_),
    .X(_09589_));
 sky130_fd_sc_hd__xor2_1 _16518_ (.A(_09588_),
    .B(_09589_),
    .X(_09590_));
 sky130_fd_sc_hd__xor2_1 _16519_ (.A(_09585_),
    .B(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__xnor2_1 _16520_ (.A(_09583_),
    .B(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__clkbuf_4 _16521_ (.A(_08587_),
    .X(_09593_));
 sky130_fd_sc_hd__nor2_1 _16522_ (.A(_09593_),
    .B(_09477_),
    .Y(_09594_));
 sky130_fd_sc_hd__clkbuf_4 _16523_ (.A(_09364_),
    .X(_09595_));
 sky130_fd_sc_hd__a21o_1 _16524_ (.A1(_09375_),
    .A2(_09482_),
    .B1(_08584_),
    .X(_09596_));
 sky130_fd_sc_hd__or3_1 _16525_ (.A(_09086_),
    .B(_09595_),
    .C(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__o21ai_1 _16526_ (.A1(_09139_),
    .A2(_09595_),
    .B1(_09596_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(_09597_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__xnor2_1 _16528_ (.A(_09594_),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__nand2_1 _16529_ (.A(net3143),
    .B(_08628_),
    .Y(_09601_));
 sky130_fd_sc_hd__a21o_2 _16530_ (.A1(_09601_),
    .A2(_09368_),
    .B1(_08313_),
    .X(_09602_));
 sky130_fd_sc_hd__a21boi_4 _16531_ (.A1(net3793),
    .A2(_09304_),
    .B1_N(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__nor2_1 _16532_ (.A(_09096_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__a221oi_4 _16533_ (.A1(_08150_),
    .A2(_08142_),
    .B1(_08183_),
    .B2(_08176_),
    .C1(_08047_),
    .Y(_09605_));
 sky130_fd_sc_hd__a21oi_2 _16534_ (.A1(_08180_),
    .A2(net77),
    .B1(_09605_),
    .Y(_09606_));
 sky130_fd_sc_hd__a31o_1 _16535_ (.A1(_08180_),
    .A2(_09605_),
    .A3(net77),
    .B1(_08296_),
    .X(_09607_));
 sky130_fd_sc_hd__o21ai_4 _16536_ (.A1(_09606_),
    .A2(_09607_),
    .B1(_08609_),
    .Y(_09608_));
 sky130_fd_sc_hd__or4_1 _16537_ (.A(net3722),
    .B(_09304_),
    .C(_09486_),
    .D(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__nand2_1 _16538_ (.A(net3185),
    .B(_08628_),
    .Y(_09610_));
 sky130_fd_sc_hd__a21oi_1 _16539_ (.A1(_09610_),
    .A2(_09489_),
    .B1(_08632_),
    .Y(_09611_));
 sky130_fd_sc_hd__xnor2_1 _16540_ (.A(_09609_),
    .B(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__xnor2_1 _16541_ (.A(_09604_),
    .B(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__nor2_1 _16542_ (.A(_09371_),
    .B(_09490_),
    .Y(_09614_));
 sky130_fd_sc_hd__a21o_1 _16543_ (.A1(_09485_),
    .A2(_09491_),
    .B1(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__xnor2_1 _16544_ (.A(_09613_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__xnor2_1 _16545_ (.A(_09600_),
    .B(_09616_),
    .Y(_09617_));
 sky130_fd_sc_hd__or2b_1 _16546_ (.A(_09496_),
    .B_N(_09492_),
    .X(_09618_));
 sky130_fd_sc_hd__a21bo_1 _16547_ (.A1(_09481_),
    .A2(_09497_),
    .B1_N(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__xnor2_1 _16548_ (.A(_09617_),
    .B(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__xnor2_1 _16549_ (.A(_09592_),
    .B(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__or2b_1 _16550_ (.A(_09498_),
    .B_N(_09500_),
    .X(_09622_));
 sky130_fd_sc_hd__a21boi_1 _16551_ (.A1(_09475_),
    .A2(_09501_),
    .B1_N(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__nor2_1 _16552_ (.A(_09621_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand2_1 _16553_ (.A(_09621_),
    .B(_09623_),
    .Y(_09625_));
 sky130_fd_sc_hd__and2b_1 _16554_ (.A_N(_09624_),
    .B(_09625_),
    .X(_09626_));
 sky130_fd_sc_hd__xnor2_2 _16555_ (.A(_09581_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__nor2_1 _16556_ (.A(_09502_),
    .B(_09504_),
    .Y(_09628_));
 sky130_fd_sc_hd__a21oi_2 _16557_ (.A1(_09463_),
    .A2(_09505_),
    .B1(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__xor2_2 _16558_ (.A(_09627_),
    .B(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__xnor2_1 _16559_ (.A(_09559_),
    .B(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__nor2_1 _16560_ (.A(_09506_),
    .B(_09507_),
    .Y(_09632_));
 sky130_fd_sc_hd__a21oi_1 _16561_ (.A1(_09442_),
    .A2(_09508_),
    .B1(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__nor2_1 _16562_ (.A(_09631_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__nand2_1 _16563_ (.A(_09631_),
    .B(_09633_),
    .Y(_09635_));
 sky130_fd_sc_hd__and2b_1 _16564_ (.A_N(_09634_),
    .B(_09635_),
    .X(_09636_));
 sky130_fd_sc_hd__xnor2_4 _16565_ (.A(_09531_),
    .B(_09636_),
    .Y(_09637_));
 sky130_fd_sc_hd__a21oi_4 _16566_ (.A1(_09414_),
    .A2(_09512_),
    .B1(_09510_),
    .Y(_09638_));
 sky130_fd_sc_hd__xnor2_4 _16567_ (.A(_09637_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__xnor2_4 _16568_ (.A(_09530_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__xnor2_4 _16569_ (.A(_09529_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__inv_2 _16570_ (.A(_09641_),
    .Y(_09642_));
 sky130_fd_sc_hd__mux2_1 _16571_ (.A0(net4063),
    .A1(net3008),
    .S(_08293_),
    .X(_09643_));
 sky130_fd_sc_hd__and2_1 _16572_ (.A(_09642_),
    .B(net3009),
    .X(_09644_));
 sky130_fd_sc_hd__or2_1 _16573_ (.A(_09642_),
    .B(net3009),
    .X(_09645_));
 sky130_fd_sc_hd__or2b_1 _16574_ (.A(_09644_),
    .B_N(_09645_),
    .X(_09646_));
 sky130_fd_sc_hd__a21o_1 _16575_ (.A1(_09521_),
    .A2(net3004),
    .B1(_09524_),
    .X(_09647_));
 sky130_fd_sc_hd__xnor2_1 _16576_ (.A(_09646_),
    .B(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__nor2_1 _16577_ (.A(net7407),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21o_1 _16578_ (.A1(net7407),
    .A2(_09648_),
    .B1(_08633_),
    .X(_09650_));
 sky130_fd_sc_hd__o221a_1 _16579_ (.A1(net4384),
    .A2(_08296_),
    .B1(_09649_),
    .B2(_09650_),
    .C1(_08239_),
    .X(_00469_));
 sky130_fd_sc_hd__a21o_1 _16580_ (.A1(_09530_),
    .A2(_09516_),
    .B1(_09639_),
    .X(_09651_));
 sky130_fd_sc_hd__o31a_4 _16581_ (.A1(_09518_),
    .A2(_09520_),
    .A3(_09640_),
    .B1(_09651_),
    .X(_09652_));
 sky130_fd_sc_hd__nor2_2 _16582_ (.A(_09637_),
    .B(_09638_),
    .Y(_09653_));
 sky130_fd_sc_hd__a21o_2 _16583_ (.A1(_09531_),
    .A2(_09635_),
    .B1(_09634_),
    .X(_09654_));
 sky130_fd_sc_hd__or2b_1 _16584_ (.A(_09558_),
    .B_N(_09533_),
    .X(_09655_));
 sky130_fd_sc_hd__a21bo_2 _16585_ (.A1(_09535_),
    .A2(_09557_),
    .B1_N(_09655_),
    .X(_09656_));
 sky130_fd_sc_hd__or2b_1 _16586_ (.A(_09542_),
    .B_N(_09556_),
    .X(_09657_));
 sky130_fd_sc_hd__o21ai_4 _16587_ (.A1(_09553_),
    .A2(_09555_),
    .B1(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__or2b_1 _16588_ (.A(_09580_),
    .B_N(_09560_),
    .X(_09659_));
 sky130_fd_sc_hd__a21bo_2 _16589_ (.A1(_09561_),
    .A2(_09579_),
    .B1_N(_09659_),
    .X(_09660_));
 sky130_fd_sc_hd__or3b_1 _16590_ (.A(_09419_),
    .B(_09540_),
    .C_N(_09133_),
    .X(_09661_));
 sky130_fd_sc_hd__nor2_2 _16591_ (.A(_09305_),
    .B(_09418_),
    .Y(_09662_));
 sky130_fd_sc_hd__a21bo_1 _16592_ (.A1(_09133_),
    .A2(_09662_),
    .B1_N(_09540_),
    .X(_09663_));
 sky130_fd_sc_hd__nand2_1 _16593_ (.A(_09661_),
    .B(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__or3b_1 _16594_ (.A(_09305_),
    .B(_09486_),
    .C_N(net7440),
    .X(_09665_));
 sky130_fd_sc_hd__buf_2 _16595_ (.A(net7441),
    .X(_09666_));
 sky130_fd_sc_hd__nor2_1 _16596_ (.A(_08326_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__xnor2_1 _16597_ (.A(_09664_),
    .B(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand2_2 _16598_ (.A(_09541_),
    .B(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__or2_1 _16599_ (.A(_09541_),
    .B(_09668_),
    .X(_09670_));
 sky130_fd_sc_hd__and2_1 _16600_ (.A(_09669_),
    .B(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__a21bo_1 _16601_ (.A1(_09549_),
    .A2(_09550_),
    .B1_N(_09548_),
    .X(_09672_));
 sky130_fd_sc_hd__a21o_1 _16602_ (.A1(_09564_),
    .A2(_09568_),
    .B1(_09565_),
    .X(_09673_));
 sky130_fd_sc_hd__or2_1 _16603_ (.A(_08454_),
    .B(_09311_),
    .X(_09674_));
 sky130_fd_sc_hd__nor2_1 _16604_ (.A(_08409_),
    .B(_08795_),
    .Y(_09675_));
 sky130_fd_sc_hd__or2_1 _16605_ (.A(_08409_),
    .B(_09250_),
    .X(_09676_));
 sky130_fd_sc_hd__or3_1 _16606_ (.A(_09091_),
    .B(_08795_),
    .C(_09676_),
    .X(_09677_));
 sky130_fd_sc_hd__o21a_1 _16607_ (.A1(_09547_),
    .A2(_09675_),
    .B1(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__xnor2_1 _16608_ (.A(_09674_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__and2_1 _16609_ (.A(_09673_),
    .B(_09679_),
    .X(_09680_));
 sky130_fd_sc_hd__nor2_1 _16610_ (.A(_09673_),
    .B(_09679_),
    .Y(_09681_));
 sky130_fd_sc_hd__nor2_1 _16611_ (.A(_09680_),
    .B(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__xnor2_1 _16612_ (.A(_09672_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__and2b_1 _16613_ (.A_N(_09551_),
    .B(_09544_),
    .X(_09684_));
 sky130_fd_sc_hd__a21oi_1 _16614_ (.A1(_09543_),
    .A2(_09552_),
    .B1(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__nor2_1 _16615_ (.A(_09683_),
    .B(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__and2_1 _16616_ (.A(_09683_),
    .B(_09685_),
    .X(_09687_));
 sky130_fd_sc_hd__nor2_1 _16617_ (.A(_09686_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__xor2_2 _16618_ (.A(_09671_),
    .B(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__xnor2_2 _16619_ (.A(_09660_),
    .B(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__xnor2_4 _16620_ (.A(_09658_),
    .B(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__a21o_1 _16621_ (.A1(_09569_),
    .A2(_09578_),
    .B1(_09576_),
    .X(_09692_));
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(_09585_),
    .B(_09590_),
    .Y(_09693_));
 sky130_fd_sc_hd__or2b_1 _16623_ (.A(_09583_),
    .B_N(_09591_),
    .X(_09694_));
 sky130_fd_sc_hd__and2_1 _16624_ (.A(_08351_),
    .B(_08352_),
    .X(_09695_));
 sky130_fd_sc_hd__o22a_1 _16625_ (.A1(_08317_),
    .A2(_09695_),
    .B1(_09562_),
    .B2(_08331_),
    .X(_09696_));
 sky130_fd_sc_hd__and3_1 _16626_ (.A(_08701_),
    .B(_08849_),
    .C(_09563_),
    .X(_09697_));
 sky130_fd_sc_hd__or2_1 _16627_ (.A(_09696_),
    .B(_09697_),
    .X(_09698_));
 sky130_fd_sc_hd__and2b_1 _16628_ (.A_N(_08707_),
    .B(_09447_),
    .X(_09699_));
 sky130_fd_sc_hd__xnor2_1 _16629_ (.A(_09698_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__or4_1 _16630_ (.A(_08470_),
    .B(_08484_),
    .C(_08574_),
    .D(_08550_),
    .X(_09701_));
 sky130_fd_sc_hd__o22ai_2 _16631_ (.A1(_08471_),
    .A2(_08574_),
    .B1(_08588_),
    .B2(_08516_),
    .Y(_09702_));
 sky130_fd_sc_hd__and2_1 _16632_ (.A(_09701_),
    .B(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__nor2_1 _16633_ (.A(_08498_),
    .B(_08565_),
    .Y(_09704_));
 sky130_fd_sc_hd__xnor2_1 _16634_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__o31a_1 _16635_ (.A1(_08564_),
    .A2(_08717_),
    .A3(_09572_),
    .B1(_09570_),
    .X(_09706_));
 sky130_fd_sc_hd__nor2_1 _16636_ (.A(_09705_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__and2_1 _16637_ (.A(_09705_),
    .B(_09706_),
    .X(_09708_));
 sky130_fd_sc_hd__nor2_1 _16638_ (.A(_09707_),
    .B(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__xnor2_1 _16639_ (.A(_09700_),
    .B(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__a21o_1 _16640_ (.A1(_09693_),
    .A2(_09694_),
    .B1(_09710_),
    .X(_09711_));
 sky130_fd_sc_hd__nand3_1 _16641_ (.A(_09693_),
    .B(_09694_),
    .C(_09710_),
    .Y(_09712_));
 sky130_fd_sc_hd__and2_1 _16642_ (.A(_09711_),
    .B(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__nand2_1 _16643_ (.A(_09692_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__or2_1 _16644_ (.A(_09692_),
    .B(_09713_),
    .X(_09715_));
 sky130_fd_sc_hd__and2_1 _16645_ (.A(_09714_),
    .B(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__nor2_1 _16646_ (.A(_09588_),
    .B(_09589_),
    .Y(_09717_));
 sky130_fd_sc_hd__a21o_1 _16647_ (.A1(_09586_),
    .A2(_09587_),
    .B1(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__a21boi_1 _16648_ (.A1(_09594_),
    .A2(_09598_),
    .B1_N(_09597_),
    .Y(_09719_));
 sky130_fd_sc_hd__nand2_1 _16649_ (.A(_08899_),
    .B(_08599_),
    .Y(_09720_));
 sky130_fd_sc_hd__nor2_1 _16650_ (.A(_09103_),
    .B(_09477_),
    .Y(_09721_));
 sky130_fd_sc_hd__xnor2_1 _16651_ (.A(_09720_),
    .B(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__nor2_1 _16652_ (.A(_08684_),
    .B(_08582_),
    .Y(_09723_));
 sky130_fd_sc_hd__xnor2_1 _16653_ (.A(_09722_),
    .B(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__xnor2_1 _16654_ (.A(_09719_),
    .B(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__xnor2_1 _16655_ (.A(_09718_),
    .B(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__or4_1 _16656_ (.A(_08584_),
    .B(_09086_),
    .C(_09483_),
    .D(_09603_),
    .X(_09727_));
 sky130_fd_sc_hd__o22ai_1 _16657_ (.A1(_09139_),
    .A2(_09484_),
    .B1(_09603_),
    .B2(_09138_),
    .Y(_09728_));
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(_09727_),
    .B(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__nor2_1 _16659_ (.A(_09593_),
    .B(_09595_),
    .Y(_09730_));
 sky130_fd_sc_hd__xnor2_1 _16660_ (.A(_09729_),
    .B(_09730_),
    .Y(_09731_));
 sky130_fd_sc_hd__a21o_2 _16661_ (.A1(_09610_),
    .A2(_09489_),
    .B1(_09304_),
    .X(_09732_));
 sky130_fd_sc_hd__nand2_1 _16662_ (.A(net3420),
    .B(_09304_),
    .Y(_09733_));
 sky130_fd_sc_hd__a21oi_1 _16663_ (.A1(_09732_),
    .A2(_09733_),
    .B1(_09096_),
    .Y(_09734_));
 sky130_fd_sc_hd__inv_2 _16664_ (.A(_08186_),
    .Y(_09735_));
 sky130_fd_sc_hd__a31o_1 _16665_ (.A1(_08180_),
    .A2(_09605_),
    .A3(net77),
    .B1(_09735_),
    .X(_09736_));
 sky130_fd_sc_hd__or4b_4 _16666_ (.A(_08181_),
    .B(_08184_),
    .C(_08186_),
    .D_N(net77),
    .X(_09737_));
 sky130_fd_sc_hd__a31o_4 _16667_ (.A1(_08633_),
    .A2(_09736_),
    .A3(_09737_),
    .B1(_08610_),
    .X(_09738_));
 sky130_fd_sc_hd__or4_4 _16668_ (.A(net3722),
    .B(_09304_),
    .C(_09486_),
    .D(_09738_),
    .X(_09739_));
 sky130_fd_sc_hd__nand2_1 _16669_ (.A(net3127),
    .B(_09486_),
    .Y(_09740_));
 sky130_fd_sc_hd__a21oi_1 _16670_ (.A1(_09740_),
    .A2(_09608_),
    .B1(_08632_),
    .Y(_09741_));
 sky130_fd_sc_hd__xnor2_2 _16671_ (.A(_09739_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__xor2_1 _16672_ (.A(_09734_),
    .B(_09742_),
    .X(_09743_));
 sky130_fd_sc_hd__a21oi_1 _16673_ (.A1(_09740_),
    .A2(_09608_),
    .B1(_09305_),
    .Y(_09744_));
 sky130_fd_sc_hd__a32o_1 _16674_ (.A1(_08613_),
    .A2(_09744_),
    .A3(_09611_),
    .B1(_09612_),
    .B2(_09604_),
    .X(_09745_));
 sky130_fd_sc_hd__xor2_1 _16675_ (.A(_09743_),
    .B(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__xnor2_1 _16676_ (.A(_09731_),
    .B(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__and2b_1 _16677_ (.A_N(_09613_),
    .B(_09615_),
    .X(_09748_));
 sky130_fd_sc_hd__a21oi_1 _16678_ (.A1(_09600_),
    .A2(_09616_),
    .B1(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__xor2_1 _16679_ (.A(_09747_),
    .B(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__xnor2_1 _16680_ (.A(_09726_),
    .B(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__and2b_1 _16681_ (.A_N(_09617_),
    .B(_09619_),
    .X(_09752_));
 sky130_fd_sc_hd__a21oi_1 _16682_ (.A1(_09592_),
    .A2(_09620_),
    .B1(_09752_),
    .Y(_09753_));
 sky130_fd_sc_hd__nor2_1 _16683_ (.A(_09751_),
    .B(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_1 _16684_ (.A(_09751_),
    .B(_09753_),
    .Y(_09755_));
 sky130_fd_sc_hd__and2b_1 _16685_ (.A_N(_09754_),
    .B(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__xnor2_1 _16686_ (.A(_09716_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__a21oi_1 _16687_ (.A1(_09581_),
    .A2(_09625_),
    .B1(_09624_),
    .Y(_09758_));
 sky130_fd_sc_hd__nor2_1 _16688_ (.A(_09757_),
    .B(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__and2_1 _16689_ (.A(_09757_),
    .B(_09758_),
    .X(_09760_));
 sky130_fd_sc_hd__nor2_2 _16690_ (.A(_09759_),
    .B(_09760_),
    .Y(_09761_));
 sky130_fd_sc_hd__xnor2_4 _16691_ (.A(_09691_),
    .B(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__nor2_1 _16692_ (.A(_09627_),
    .B(_09629_),
    .Y(_09763_));
 sky130_fd_sc_hd__a21oi_2 _16693_ (.A1(_09559_),
    .A2(_09630_),
    .B1(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__xor2_4 _16694_ (.A(_09762_),
    .B(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__xnor2_4 _16695_ (.A(_09656_),
    .B(_09765_),
    .Y(_09766_));
 sky130_fd_sc_hd__xnor2_4 _16696_ (.A(_09654_),
    .B(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__xor2_4 _16697_ (.A(_09653_),
    .B(_09767_),
    .X(_09768_));
 sky130_fd_sc_hd__xnor2_4 _16698_ (.A(_09652_),
    .B(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__mux2_1 _16699_ (.A0(net7446),
    .A1(net3028),
    .S(_08293_),
    .X(_09770_));
 sky130_fd_sc_hd__nor2_1 _16700_ (.A(_09769_),
    .B(net3029),
    .Y(_09771_));
 sky130_fd_sc_hd__and2_1 _16701_ (.A(_09769_),
    .B(net3029),
    .X(_09772_));
 sky130_fd_sc_hd__nor2_1 _16702_ (.A(_09771_),
    .B(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__a21oi_1 _16703_ (.A1(_09645_),
    .A2(_09647_),
    .B1(_09644_),
    .Y(_09774_));
 sky130_fd_sc_hd__xnor2_1 _16704_ (.A(net7407),
    .B(_09774_),
    .Y(_09775_));
 sky130_fd_sc_hd__nor2_1 _16705_ (.A(_09773_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__a21o_1 _16706_ (.A1(_09773_),
    .A2(_09775_),
    .B1(_08633_),
    .X(_09777_));
 sky130_fd_sc_hd__o221a_1 _16707_ (.A1(net4519),
    .A2(_08296_),
    .B1(_09776_),
    .B2(_09777_),
    .C1(_08239_),
    .X(_00470_));
 sky130_fd_sc_hd__o21ba_1 _16708_ (.A1(_09771_),
    .A2(_09774_),
    .B1_N(_09772_),
    .X(_09778_));
 sky130_fd_sc_hd__inv_2 _16709_ (.A(_09768_),
    .Y(_09779_));
 sky130_fd_sc_hd__nand2_1 _16710_ (.A(_09653_),
    .B(_09767_),
    .Y(_09780_));
 sky130_fd_sc_hd__o21ai_2 _16711_ (.A1(_09652_),
    .A2(_09779_),
    .B1(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__or2b_2 _16712_ (.A(_09766_),
    .B_N(_09654_),
    .X(_09782_));
 sky130_fd_sc_hd__or3_1 _16713_ (.A(net4828),
    .B(_09305_),
    .C(_09486_),
    .X(_09783_));
 sky130_fd_sc_hd__buf_4 _16714_ (.A(_09783_),
    .X(_09784_));
 sky130_fd_sc_hd__or2b_1 _16715_ (.A(_09690_),
    .B_N(_09658_),
    .X(_09785_));
 sky130_fd_sc_hd__a21boi_2 _16716_ (.A1(_09660_),
    .A2(_09689_),
    .B1_N(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__or3b_2 _16717_ (.A(_09784_),
    .B(_09786_),
    .C_N(_08326_),
    .X(_09787_));
 sky130_fd_sc_hd__or2_1 _16718_ (.A(_09669_),
    .B(_09786_),
    .X(_09788_));
 sky130_fd_sc_hd__nand2_1 _16719_ (.A(_09669_),
    .B(_09786_),
    .Y(_09789_));
 sky130_fd_sc_hd__and3_1 _16720_ (.A(net7554),
    .B(_06211_),
    .C(_08314_),
    .X(_09790_));
 sky130_fd_sc_hd__a22o_1 _16721_ (.A1(_09788_),
    .A2(_09789_),
    .B1(net7378),
    .B2(_08326_),
    .X(_09791_));
 sky130_fd_sc_hd__and2_1 _16722_ (.A(_09787_),
    .B(_09791_),
    .X(_09792_));
 sky130_fd_sc_hd__a21o_1 _16723_ (.A1(_09671_),
    .A2(_09688_),
    .B1(_09686_),
    .X(_09793_));
 sky130_fd_sc_hd__nor2_1 _16724_ (.A(_09305_),
    .B(_09536_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_1 _16725_ (.A(_09133_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__o22a_1 _16726_ (.A1(_09091_),
    .A2(_09312_),
    .B1(_09419_),
    .B2(_08724_),
    .X(_09796_));
 sky130_fd_sc_hd__nand2_1 _16727_ (.A(_09051_),
    .B(_09662_),
    .Y(_09797_));
 sky130_fd_sc_hd__or2_1 _16728_ (.A(_09674_),
    .B(_09797_),
    .X(_09798_));
 sky130_fd_sc_hd__and2b_1 _16729_ (.A_N(_09796_),
    .B(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__xor2_1 _16730_ (.A(_09795_),
    .B(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__o31a_1 _16731_ (.A1(_08326_),
    .A2(_09664_),
    .A3(_09666_),
    .B1(_09661_),
    .X(_09801_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_09800_),
    .B(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__and2_1 _16733_ (.A(_09800_),
    .B(_09801_),
    .X(_09803_));
 sky130_fd_sc_hd__nor2_1 _16734_ (.A(_09802_),
    .B(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__clkbuf_4 _16735_ (.A(_09666_),
    .X(_09805_));
 sky130_fd_sc_hd__nor2_1 _16736_ (.A(_08310_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__xor2_1 _16737_ (.A(_09804_),
    .B(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__or2b_1 _16738_ (.A(_09674_),
    .B_N(_09678_),
    .X(_09808_));
 sky130_fd_sc_hd__nand2_1 _16739_ (.A(_09677_),
    .B(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__inv_2 _16740_ (.A(_09696_),
    .Y(_09810_));
 sky130_fd_sc_hd__a21o_1 _16741_ (.A1(_09810_),
    .A2(_09699_),
    .B1(_09697_),
    .X(_09811_));
 sky130_fd_sc_hd__a2bb2o_1 _16742_ (.A1_N(_09562_),
    .A2_N(_08707_),
    .B1(_09306_),
    .B2(_08962_),
    .X(_09812_));
 sky130_fd_sc_hd__or2_2 _16743_ (.A(_08372_),
    .B(_08795_),
    .X(_09813_));
 sky130_fd_sc_hd__or3b_1 _16744_ (.A(_08707_),
    .B(_09813_),
    .C_N(_08962_),
    .X(_09814_));
 sky130_fd_sc_hd__nand2_1 _16745_ (.A(_09812_),
    .B(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__xor2_1 _16746_ (.A(_09676_),
    .B(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__and2_1 _16747_ (.A(_09811_),
    .B(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__or2_1 _16748_ (.A(_09811_),
    .B(_09816_),
    .X(_09818_));
 sky130_fd_sc_hd__and2b_1 _16749_ (.A_N(_09817_),
    .B(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__xnor2_1 _16750_ (.A(_09809_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__a21oi_1 _16751_ (.A1(_09672_),
    .A2(_09682_),
    .B1(_09680_),
    .Y(_09821_));
 sky130_fd_sc_hd__nor2_1 _16752_ (.A(_09820_),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__and2_1 _16753_ (.A(_09820_),
    .B(_09821_),
    .X(_09823_));
 sky130_fd_sc_hd__nor2_1 _16754_ (.A(_09822_),
    .B(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__xnor2_1 _16755_ (.A(_09807_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__a21o_1 _16756_ (.A1(_09711_),
    .A2(_09714_),
    .B1(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__nand3_1 _16757_ (.A(_09711_),
    .B(_09714_),
    .C(_09825_),
    .Y(_09827_));
 sky130_fd_sc_hd__nand2_1 _16758_ (.A(_09826_),
    .B(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__xnor2_1 _16759_ (.A(_09793_),
    .B(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__a21o_1 _16760_ (.A1(_09700_),
    .A2(_09709_),
    .B1(_09707_),
    .X(_09830_));
 sky130_fd_sc_hd__or2_1 _16761_ (.A(_09719_),
    .B(_09724_),
    .X(_09831_));
 sky130_fd_sc_hd__or2b_1 _16762_ (.A(_09725_),
    .B_N(_09718_),
    .X(_09832_));
 sky130_fd_sc_hd__nand2_2 _16763_ (.A(_08701_),
    .B(_08849_),
    .Y(_09833_));
 sky130_fd_sc_hd__or4_2 _16764_ (.A(_08317_),
    .B(_08498_),
    .C(_08588_),
    .D(_08556_),
    .X(_09834_));
 sky130_fd_sc_hd__inv_2 _16765_ (.A(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__o22a_1 _16766_ (.A1(_08717_),
    .A2(_08588_),
    .B1(_08556_),
    .B2(_08317_),
    .X(_09836_));
 sky130_fd_sc_hd__nor2_1 _16767_ (.A(_09835_),
    .B(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__xnor2_1 _16768_ (.A(_09833_),
    .B(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__or2_1 _16769_ (.A(_08873_),
    .B(_08574_),
    .X(_09839_));
 sky130_fd_sc_hd__nor2_1 _16770_ (.A(_08684_),
    .B(_09216_),
    .Y(_09840_));
 sky130_fd_sc_hd__nor2_1 _16771_ (.A(_08872_),
    .B(_08582_),
    .Y(_09841_));
 sky130_fd_sc_hd__xor2_1 _16772_ (.A(_09840_),
    .B(_09841_),
    .X(_09842_));
 sky130_fd_sc_hd__xor2_1 _16773_ (.A(_09839_),
    .B(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__a21boi_2 _16774_ (.A1(_09702_),
    .A2(_09704_),
    .B1_N(_09701_),
    .Y(_09844_));
 sky130_fd_sc_hd__xor2_1 _16775_ (.A(_09843_),
    .B(_09844_),
    .X(_09845_));
 sky130_fd_sc_hd__xnor2_1 _16776_ (.A(_09838_),
    .B(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__a21o_1 _16777_ (.A1(_09831_),
    .A2(_09832_),
    .B1(_09846_),
    .X(_09847_));
 sky130_fd_sc_hd__nand3_1 _16778_ (.A(_09831_),
    .B(_09832_),
    .C(_09846_),
    .Y(_09848_));
 sky130_fd_sc_hd__nand2_1 _16779_ (.A(_09847_),
    .B(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__xnor2_1 _16780_ (.A(_09830_),
    .B(_09849_),
    .Y(_09850_));
 sky130_fd_sc_hd__and2_1 _16781_ (.A(_09722_),
    .B(_09723_),
    .X(_09851_));
 sky130_fd_sc_hd__a31o_1 _16782_ (.A1(_08899_),
    .A2(_08599_),
    .A3(_09721_),
    .B1(_09851_),
    .X(_09852_));
 sky130_fd_sc_hd__o31a_1 _16783_ (.A1(_09593_),
    .A2(_09595_),
    .A3(_09729_),
    .B1(_09727_),
    .X(_09853_));
 sky130_fd_sc_hd__or2_1 _16784_ (.A(_09064_),
    .B(_09477_),
    .X(_09854_));
 sky130_fd_sc_hd__or2_2 _16785_ (.A(_08587_),
    .B(_09483_),
    .X(_09855_));
 sky130_fd_sc_hd__nor2_1 _16786_ (.A(_09103_),
    .B(_09595_),
    .Y(_09856_));
 sky130_fd_sc_hd__xnor2_1 _16787_ (.A(_09855_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__xnor2_1 _16788_ (.A(_09854_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__xnor2_1 _16789_ (.A(_09853_),
    .B(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__xor2_1 _16790_ (.A(_09852_),
    .B(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__clkbuf_4 _16791_ (.A(_09603_),
    .X(_09861_));
 sky130_fd_sc_hd__nor2_1 _16792_ (.A(_09139_),
    .B(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__a21o_2 _16793_ (.A1(_09740_),
    .A2(_09608_),
    .B1(_09304_),
    .X(_09863_));
 sky130_fd_sc_hd__nand2_1 _16794_ (.A(net3717),
    .B(_09304_),
    .Y(_09864_));
 sky130_fd_sc_hd__a21o_1 _16795_ (.A1(_09863_),
    .A2(_09864_),
    .B1(_08626_),
    .X(_09865_));
 sky130_fd_sc_hd__a21oi_1 _16796_ (.A1(_09732_),
    .A2(_09733_),
    .B1(_08584_),
    .Y(_09866_));
 sky130_fd_sc_hd__xnor2_1 _16797_ (.A(_09865_),
    .B(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__xor2_1 _16798_ (.A(_09862_),
    .B(_09867_),
    .X(_09868_));
 sky130_fd_sc_hd__o21ai_1 _16799_ (.A1(_08188_),
    .A2(_09737_),
    .B1(_08633_),
    .Y(_09869_));
 sky130_fd_sc_hd__a22o_2 _16800_ (.A1(net3042),
    .A2(_09486_),
    .B1(_08609_),
    .B2(_09869_),
    .X(_09870_));
 sky130_fd_sc_hd__a21o_1 _16801_ (.A1(_08755_),
    .A2(_09870_),
    .B1(_09790_),
    .X(_09871_));
 sky130_fd_sc_hd__or3b_1 _16802_ (.A(net4828),
    .B(_08664_),
    .C_N(_09870_),
    .X(_09872_));
 sky130_fd_sc_hd__nand2_1 _16803_ (.A(net3528),
    .B(_09486_),
    .Y(_09873_));
 sky130_fd_sc_hd__a21oi_1 _16804_ (.A1(_09873_),
    .A2(_09738_),
    .B1(_08632_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand3_1 _16805_ (.A(_09871_),
    .B(_09872_),
    .C(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__a21o_1 _16806_ (.A1(_09871_),
    .A2(_09872_),
    .B1(_09874_),
    .X(_09876_));
 sky130_fd_sc_hd__a21oi_1 _16807_ (.A1(_09873_),
    .A2(_09738_),
    .B1(_09305_),
    .Y(_09877_));
 sky130_fd_sc_hd__a32o_1 _16808_ (.A1(_08613_),
    .A2(_09877_),
    .A3(_09741_),
    .B1(_09742_),
    .B2(_09734_),
    .X(_09878_));
 sky130_fd_sc_hd__nand3_1 _16809_ (.A(_09875_),
    .B(_09876_),
    .C(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__a21o_1 _16810_ (.A1(_09875_),
    .A2(_09876_),
    .B1(_09878_),
    .X(_09880_));
 sky130_fd_sc_hd__nand3_1 _16811_ (.A(_09868_),
    .B(_09879_),
    .C(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__a21o_1 _16812_ (.A1(_09879_),
    .A2(_09880_),
    .B1(_09868_),
    .X(_09882_));
 sky130_fd_sc_hd__nand2_1 _16813_ (.A(_09743_),
    .B(_09745_),
    .Y(_09883_));
 sky130_fd_sc_hd__a21bo_1 _16814_ (.A1(_09731_),
    .A2(_09746_),
    .B1_N(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__nand3_1 _16815_ (.A(_09881_),
    .B(_09882_),
    .C(_09884_),
    .Y(_09885_));
 sky130_fd_sc_hd__a21o_1 _16816_ (.A1(_09881_),
    .A2(_09882_),
    .B1(_09884_),
    .X(_09886_));
 sky130_fd_sc_hd__nand3_1 _16817_ (.A(_09860_),
    .B(_09885_),
    .C(_09886_),
    .Y(_09887_));
 sky130_fd_sc_hd__a21o_1 _16818_ (.A1(_09885_),
    .A2(_09886_),
    .B1(_09860_),
    .X(_09888_));
 sky130_fd_sc_hd__nor2_1 _16819_ (.A(_09747_),
    .B(_09749_),
    .Y(_09889_));
 sky130_fd_sc_hd__a21o_1 _16820_ (.A1(_09726_),
    .A2(_09750_),
    .B1(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__nand3_1 _16821_ (.A(_09887_),
    .B(_09888_),
    .C(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__a21o_1 _16822_ (.A1(_09887_),
    .A2(_09888_),
    .B1(_09890_),
    .X(_09892_));
 sky130_fd_sc_hd__and3_1 _16823_ (.A(_09850_),
    .B(_09891_),
    .C(_09892_),
    .X(_09893_));
 sky130_fd_sc_hd__a21oi_1 _16824_ (.A1(_09891_),
    .A2(_09892_),
    .B1(_09850_),
    .Y(_09894_));
 sky130_fd_sc_hd__or2_4 _16825_ (.A(_09893_),
    .B(_09894_),
    .X(_09895_));
 sky130_fd_sc_hd__a21oi_2 _16826_ (.A1(_09716_),
    .A2(_09755_),
    .B1(_09754_),
    .Y(_09896_));
 sky130_fd_sc_hd__xor2_2 _16827_ (.A(_09895_),
    .B(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__xnor2_2 _16828_ (.A(_09829_),
    .B(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__a21oi_1 _16829_ (.A1(_09691_),
    .A2(_09761_),
    .B1(_09759_),
    .Y(_09899_));
 sky130_fd_sc_hd__xor2_2 _16830_ (.A(_09898_),
    .B(_09899_),
    .X(_09900_));
 sky130_fd_sc_hd__xnor2_2 _16831_ (.A(_09792_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__nor2_1 _16832_ (.A(_09762_),
    .B(_09764_),
    .Y(_09902_));
 sky130_fd_sc_hd__a21oi_1 _16833_ (.A1(_09656_),
    .A2(_09765_),
    .B1(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__nor2_2 _16834_ (.A(_09901_),
    .B(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__and2_1 _16835_ (.A(_09901_),
    .B(_09903_),
    .X(_09905_));
 sky130_fd_sc_hd__or2_2 _16836_ (.A(_09904_),
    .B(_09905_),
    .X(_09906_));
 sky130_fd_sc_hd__xnor2_4 _16837_ (.A(_09782_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__xnor2_4 _16838_ (.A(_09781_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__mux2_1 _16839_ (.A0(net4288),
    .A1(net4105),
    .S(net4088),
    .X(_09909_));
 sky130_fd_sc_hd__xor2_1 _16840_ (.A(_09297_),
    .B(net4106),
    .X(_09910_));
 sky130_fd_sc_hd__xnor2_1 _16841_ (.A(_09908_),
    .B(net4107),
    .Y(_09911_));
 sky130_fd_sc_hd__and2_1 _16842_ (.A(_09778_),
    .B(_09911_),
    .X(_09912_));
 sky130_fd_sc_hd__o21ai_1 _16843_ (.A1(_09778_),
    .A2(_09911_),
    .B1(_08296_),
    .Y(_09913_));
 sky130_fd_sc_hd__o221a_1 _16844_ (.A1(net7368),
    .A2(_08296_),
    .B1(_09912_),
    .B2(_09913_),
    .C1(_08195_),
    .X(_00471_));
 sky130_fd_sc_hd__o21ai_1 _16845_ (.A1(_04164_),
    .A2(_04161_),
    .B1(net3975),
    .Y(_09914_));
 sky130_fd_sc_hd__nor2_1 _16846_ (.A(_04165_),
    .B(net3976),
    .Y(_09915_));
 sky130_fd_sc_hd__and4_1 _16847_ (.A(_04760_),
    .B(_04812_),
    .C(_04852_),
    .D(net3977),
    .X(_09916_));
 sky130_fd_sc_hd__clkbuf_1 _16848_ (.A(net3978),
    .X(_09917_));
 sky130_fd_sc_hd__or2_1 _16849_ (.A(_04241_),
    .B(net3979),
    .X(_09918_));
 sky130_fd_sc_hd__clkbuf_4 _16850_ (.A(_09918_),
    .X(_09919_));
 sky130_fd_sc_hd__nor2_1 _16851_ (.A(_04160_),
    .B(_09919_),
    .Y(_00472_));
 sky130_fd_sc_hd__a21oi_1 _16852_ (.A1(net3870),
    .A2(_04795_),
    .B1(_09919_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2_4 _16853_ (.A(_04241_),
    .B(net3979),
    .Y(_09920_));
 sky130_fd_sc_hd__o21ai_1 _16854_ (.A1(_04727_),
    .A2(_04725_),
    .B1(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__nor2_1 _16855_ (.A(net3989),
    .B(_09921_),
    .Y(_00474_));
 sky130_fd_sc_hd__nor2_1 _16856_ (.A(net3910),
    .B(_09919_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _16857_ (.A(net3762),
    .B(_09919_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _16858_ (.A(net4011),
    .B(_09919_),
    .Y(_00477_));
 sky130_fd_sc_hd__and2_1 _16859_ (.A(net4038),
    .B(_09920_),
    .X(_09922_));
 sky130_fd_sc_hd__clkbuf_1 _16860_ (.A(net4039),
    .X(_00478_));
 sky130_fd_sc_hd__and2_1 _16861_ (.A(net4074),
    .B(_09920_),
    .X(_09923_));
 sky130_fd_sc_hd__clkbuf_1 _16862_ (.A(net4075),
    .X(_00479_));
 sky130_fd_sc_hd__and4_1 _16863_ (.A(_04165_),
    .B(_04637_),
    .C(_04603_),
    .D(_04760_),
    .X(_09924_));
 sky130_fd_sc_hd__and3_1 _16864_ (.A(_04162_),
    .B(_04812_),
    .C(net4054),
    .X(_09925_));
 sky130_fd_sc_hd__a31o_1 _16865_ (.A1(_04777_),
    .A2(net3989),
    .A3(net4054),
    .B1(_04162_),
    .X(_09926_));
 sky130_fd_sc_hd__and3b_1 _16866_ (.A_N(_09925_),
    .B(_09920_),
    .C(net4055),
    .X(_09927_));
 sky130_fd_sc_hd__clkbuf_1 _16867_ (.A(net4056),
    .X(_00480_));
 sky130_fd_sc_hd__a21oi_1 _16868_ (.A1(net3993),
    .A2(_09925_),
    .B1(_09919_),
    .Y(_09928_));
 sky130_fd_sc_hd__o21a_1 _16869_ (.A1(net3993),
    .A2(_09925_),
    .B1(_09928_),
    .X(_00481_));
 sky130_fd_sc_hd__inv_2 _16870_ (.A(net3979),
    .Y(_09929_));
 sky130_fd_sc_hd__or3_4 _16871_ (.A(_04818_),
    .B(net3535),
    .C(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__and2_1 _16872_ (.A(_04622_),
    .B(_09930_),
    .X(_09931_));
 sky130_fd_sc_hd__clkbuf_4 _16873_ (.A(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__clkbuf_8 _16874_ (.A(_09932_),
    .X(_09933_));
 sky130_fd_sc_hd__clkbuf_4 _16875_ (.A(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__nor2_4 _16876_ (.A(_04632_),
    .B(_09930_),
    .Y(_09935_));
 sky130_fd_sc_hd__clkbuf_4 _16877_ (.A(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__a22o_1 _16878_ (.A1(net4532),
    .A2(_09934_),
    .B1(_09936_),
    .B2(net4088),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _16879_ (.A1(net4275),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08074_),
    .X(_00483_));
 sky130_fd_sc_hd__a22o_1 _16880_ (.A1(net4317),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08086_),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _16881_ (.A1(net4278),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08096_),
    .X(_00485_));
 sky130_fd_sc_hd__a22o_1 _16882_ (.A1(net4265),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08106_),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _16883_ (.A1(net6023),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08117_),
    .X(_00487_));
 sky130_fd_sc_hd__a22o_1 _16884_ (.A1(net4284),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08125_),
    .X(_00488_));
 sky130_fd_sc_hd__a22o_1 _16885_ (.A1(net4611),
    .A2(_09934_),
    .B1(_09936_),
    .B2(net7437),
    .X(_00489_));
 sky130_fd_sc_hd__a22o_1 _16886_ (.A1(net4344),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08137_),
    .X(_00490_));
 sky130_fd_sc_hd__a22o_1 _16887_ (.A1(net4391),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_08144_),
    .X(_00491_));
 sky130_fd_sc_hd__clkbuf_4 _16888_ (.A(_09933_),
    .X(_09937_));
 sky130_fd_sc_hd__buf_4 _16889_ (.A(_09935_),
    .X(_09938_));
 sky130_fd_sc_hd__a22o_1 _16890_ (.A1(net4509),
    .A2(_09937_),
    .B1(_09938_),
    .B2(_08152_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _16891_ (.A1(net4109),
    .A2(_09937_),
    .B1(_09938_),
    .B2(_08155_),
    .X(_00493_));
 sky130_fd_sc_hd__a22o_1 _16892_ (.A1(net4239),
    .A2(_09937_),
    .B1(_09938_),
    .B2(net1422),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _16893_ (.A1(net4271),
    .A2(_09937_),
    .B1(_09938_),
    .B2(net1189),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _16894_ (.A1(net4303),
    .A2(_09937_),
    .B1(_09938_),
    .B2(net1304),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _16895_ (.A1(net4280),
    .A2(_09937_),
    .B1(_09938_),
    .B2(net1393),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _16896_ (.A1(net4254),
    .A2(_09937_),
    .B1(_09938_),
    .B2(net1495),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _16897_ (.A1(net773),
    .A2(_09937_),
    .B1(_09938_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _16898_ (.A1(net839),
    .A2(_09937_),
    .B1(_09938_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _16899_ (.A1(net1011),
    .A2(_09937_),
    .B1(_09938_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00501_));
 sky130_fd_sc_hd__clkbuf_4 _16900_ (.A(_09933_),
    .X(_09939_));
 sky130_fd_sc_hd__clkbuf_4 _16901_ (.A(_09935_),
    .X(_09940_));
 sky130_fd_sc_hd__a22o_1 _16902_ (.A1(net890),
    .A2(_09939_),
    .B1(_09940_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16903_ (.A1(net5379),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net3206),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _16904_ (.A1(net5471),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net3356),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _16905_ (.A1(net5310),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net3262),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16906_ (.A1(net4152),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net645),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _16907_ (.A1(net4146),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net6253),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _16908_ (.A1(net4130),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net6278),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _16909_ (.A1(net4173),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net6281),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_1 _16910_ (.A1(net4167),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net6259),
    .X(_00510_));
 sky130_fd_sc_hd__a22o_1 _16911_ (.A1(net4179),
    .A2(_09939_),
    .B1(_09940_),
    .B2(net7552),
    .X(_00511_));
 sky130_fd_sc_hd__clkbuf_4 _16912_ (.A(_09933_),
    .X(_09941_));
 sky130_fd_sc_hd__clkbuf_4 _16913_ (.A(_09935_),
    .X(_09942_));
 sky130_fd_sc_hd__a22o_1 _16914_ (.A1(net1100),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net7476),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16915_ (.A1(net1144),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net6123),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _16916_ (.A1(net4186),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net6098),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _16917_ (.A1(net4143),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net6148),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16918_ (.A1(net4160),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net6150),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _16919_ (.A1(net4176),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net6146),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16920_ (.A1(net4133),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net7442),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _16921_ (.A1(net4136),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net7440),
    .X(_00519_));
 sky130_fd_sc_hd__a22o_1 _16922_ (.A1(net4155),
    .A2(_09941_),
    .B1(_09942_),
    .B2(net7554),
    .X(_00520_));
 sky130_fd_sc_hd__or2_4 _16923_ (.A(_08246_),
    .B(_09930_),
    .X(_09943_));
 sky130_fd_sc_hd__mux2_1 _16924_ (.A0(_04693_),
    .A1(net3378),
    .S(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__clkbuf_1 _16925_ (.A(net3379),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _16926_ (.A0(_04692_),
    .A1(net3218),
    .S(_09943_),
    .X(_09945_));
 sky130_fd_sc_hd__clkbuf_1 _16927_ (.A(net3219),
    .X(_00522_));
 sky130_fd_sc_hd__xor2_1 _16928_ (.A(net2807),
    .B(_09294_),
    .X(_09946_));
 sky130_fd_sc_hd__xor2_2 _16929_ (.A(net3265),
    .B(_09294_),
    .X(_09947_));
 sky130_fd_sc_hd__xnor2_2 _16930_ (.A(_06229_),
    .B(_09294_),
    .Y(_09948_));
 sky130_fd_sc_hd__or2_1 _16931_ (.A(_06222_),
    .B(_09294_),
    .X(_09949_));
 sky130_fd_sc_hd__xnor2_1 _16932_ (.A(_06221_),
    .B(_08381_),
    .Y(_09950_));
 sky130_fd_sc_hd__nand2_1 _16933_ (.A(_06217_),
    .B(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__o21ai_1 _16934_ (.A1(_06221_),
    .A2(_09295_),
    .B1(_09951_),
    .Y(_09952_));
 sky130_fd_sc_hd__xnor2_1 _16935_ (.A(_06213_),
    .B(_09294_),
    .Y(_09953_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(_09952_),
    .B(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__o21ai_1 _16937_ (.A1(_06213_),
    .A2(_09295_),
    .B1(_09954_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(_06222_),
    .B(_09294_),
    .Y(_09956_));
 sky130_fd_sc_hd__a21bo_1 _16939_ (.A1(_09949_),
    .A2(_09955_),
    .B1_N(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__o21a_1 _16940_ (.A1(net4874),
    .A2(net3265),
    .B1(_09294_),
    .X(_09958_));
 sky130_fd_sc_hd__a31o_1 _16941_ (.A1(_09947_),
    .A2(_09948_),
    .A3(_09957_),
    .B1(net4875),
    .X(_09959_));
 sky130_fd_sc_hd__or2_1 _16942_ (.A(_09946_),
    .B(net4876),
    .X(_09960_));
 sky130_fd_sc_hd__nand2_1 _16943_ (.A(_09946_),
    .B(net4876),
    .Y(_09961_));
 sky130_fd_sc_hd__nand2_1 _16944_ (.A(_06383_),
    .B(_06344_),
    .Y(_09962_));
 sky130_fd_sc_hd__a21oi_1 _16945_ (.A1(net4900),
    .A2(_09962_),
    .B1(_06203_),
    .Y(_09963_));
 sky130_fd_sc_hd__a211o_1 _16946_ (.A1(_06204_),
    .A2(_06211_),
    .B1(net4901),
    .C1(_06391_),
    .X(_09964_));
 sky130_fd_sc_hd__nor2_2 _16947_ (.A(_06206_),
    .B(net4902),
    .Y(_09965_));
 sky130_fd_sc_hd__buf_4 _16948_ (.A(net4902),
    .X(_09966_));
 sky130_fd_sc_hd__a32o_1 _16949_ (.A1(_09960_),
    .A2(net4877),
    .A3(_09965_),
    .B1(_09966_),
    .B2(net2807),
    .X(_00523_));
 sky130_fd_sc_hd__xor2_1 _16950_ (.A(net5969),
    .B(_09294_),
    .X(_09967_));
 sky130_fd_sc_hd__buf_2 _16951_ (.A(_09294_),
    .X(_09968_));
 sky130_fd_sc_hd__a21bo_1 _16952_ (.A1(net2807),
    .A2(_09968_),
    .B1_N(net4877),
    .X(_09969_));
 sky130_fd_sc_hd__xor2_1 _16953_ (.A(_09967_),
    .B(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__a22o_1 _16954_ (.A1(net5969),
    .A2(_09966_),
    .B1(_09965_),
    .B2(_09970_),
    .X(_00524_));
 sky130_fd_sc_hd__and2_1 _16955_ (.A(net4922),
    .B(_09968_),
    .X(_09971_));
 sky130_fd_sc_hd__nor2_1 _16956_ (.A(net4922),
    .B(_09968_),
    .Y(_09972_));
 sky130_fd_sc_hd__nor2_1 _16957_ (.A(_09971_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__and2_1 _16958_ (.A(_09948_),
    .B(_09957_),
    .X(_09974_));
 sky130_fd_sc_hd__and4_1 _16959_ (.A(_09946_),
    .B(_09947_),
    .C(_09974_),
    .D(_09967_),
    .X(_09975_));
 sky130_fd_sc_hd__o21a_1 _16960_ (.A1(net2611),
    .A2(net2807),
    .B1(_09968_),
    .X(_09976_));
 sky130_fd_sc_hd__or3_1 _16961_ (.A(net4875),
    .B(_09975_),
    .C(_09976_),
    .X(_09977_));
 sky130_fd_sc_hd__xor2_1 _16962_ (.A(_09973_),
    .B(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__a22o_1 _16963_ (.A1(net4922),
    .A2(_09966_),
    .B1(_09965_),
    .B2(_09978_),
    .X(_00525_));
 sky130_fd_sc_hd__xnor2_1 _16964_ (.A(net5746),
    .B(_09968_),
    .Y(_09979_));
 sky130_fd_sc_hd__a21o_1 _16965_ (.A1(_09973_),
    .A2(_09977_),
    .B1(_09971_),
    .X(_09980_));
 sky130_fd_sc_hd__xnor2_1 _16966_ (.A(_09979_),
    .B(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__a22o_1 _16967_ (.A1(net5746),
    .A2(_09966_),
    .B1(_09965_),
    .B2(_09981_),
    .X(_00526_));
 sky130_fd_sc_hd__o21a_1 _16968_ (.A1(net2787),
    .A2(_09968_),
    .B1(_09980_),
    .X(_09982_));
 sky130_fd_sc_hd__a21oi_1 _16969_ (.A1(net2787),
    .A2(_09968_),
    .B1(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__xnor2_1 _16970_ (.A(net5420),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__or2_1 _16971_ (.A(_09968_),
    .B(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__nand2_1 _16972_ (.A(_09968_),
    .B(_09984_),
    .Y(_09986_));
 sky130_fd_sc_hd__a32o_1 _16973_ (.A1(_09965_),
    .A2(_09985_),
    .A3(_09986_),
    .B1(_09966_),
    .B2(net5420),
    .X(_00527_));
 sky130_fd_sc_hd__buf_4 _16974_ (.A(net3508),
    .X(_09987_));
 sky130_fd_sc_hd__nand2_1 _16975_ (.A(net4568),
    .B(net4566),
    .Y(_09988_));
 sky130_fd_sc_hd__or2_1 _16976_ (.A(net4568),
    .B(net4566),
    .X(_09989_));
 sky130_fd_sc_hd__and2b_1 _16977_ (.A_N(_09170_),
    .B(_09121_),
    .X(_09990_));
 sky130_fd_sc_hd__a21oi_1 _16978_ (.A1(_09990_),
    .A2(_09169_),
    .B1(net3508),
    .Y(_09991_));
 sky130_fd_sc_hd__o21a_1 _16979_ (.A1(_09990_),
    .A2(_09169_),
    .B1(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__a31o_1 _16980_ (.A1(_09987_),
    .A2(_09988_),
    .A3(_09989_),
    .B1(_09992_),
    .X(_09993_));
 sky130_fd_sc_hd__mux2_1 _16981_ (.A0(_09993_),
    .A1(net4568),
    .S(_09966_),
    .X(_09994_));
 sky130_fd_sc_hd__clkbuf_1 _16982_ (.A(_09994_),
    .X(_00528_));
 sky130_fd_sc_hd__nand2_1 _16983_ (.A(net4507),
    .B(net4579),
    .Y(_09995_));
 sky130_fd_sc_hd__or2_1 _16984_ (.A(net4507),
    .B(net4579),
    .X(_09996_));
 sky130_fd_sc_hd__nand2_1 _16985_ (.A(_09995_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__xnor2_1 _16986_ (.A(_09988_),
    .B(_09997_),
    .Y(_09998_));
 sky130_fd_sc_hd__buf_6 _16987_ (.A(net3508),
    .X(_09999_));
 sky130_fd_sc_hd__nor2_1 _16988_ (.A(_09171_),
    .B(_09173_),
    .Y(_10000_));
 sky130_fd_sc_hd__and2_1 _16989_ (.A(_09171_),
    .B(_09173_),
    .X(_10001_));
 sky130_fd_sc_hd__or3_2 _16990_ (.A(_09999_),
    .B(_10000_),
    .C(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__o21ai_1 _16991_ (.A1(_06206_),
    .A2(_09998_),
    .B1(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__mux2_1 _16992_ (.A0(_10003_),
    .A1(net4507),
    .S(_09966_),
    .X(_10004_));
 sky130_fd_sc_hd__clkbuf_1 _16993_ (.A(_10004_),
    .X(_00529_));
 sky130_fd_sc_hd__o21a_1 _16994_ (.A1(_09988_),
    .A2(_09997_),
    .B1(_09995_),
    .X(_10005_));
 sky130_fd_sc_hd__nor2_1 _16995_ (.A(net4689),
    .B(net4570),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_1 _16996_ (.A(net4689),
    .B(net4570),
    .Y(_10007_));
 sky130_fd_sc_hd__or2b_1 _16997_ (.A(_10006_),
    .B_N(_10007_),
    .X(_10008_));
 sky130_fd_sc_hd__xnor2_1 _16998_ (.A(_10005_),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__buf_4 _16999_ (.A(_06205_),
    .X(_10010_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_10010_),
    .B(_09286_),
    .Y(_10011_));
 sky130_fd_sc_hd__o21ai_1 _17001_ (.A1(_06206_),
    .A2(_10009_),
    .B1(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__mux2_1 _17002_ (.A0(_10012_),
    .A1(net4689),
    .S(_09966_),
    .X(_10013_));
 sky130_fd_sc_hd__clkbuf_1 _17003_ (.A(_10013_),
    .X(_00530_));
 sky130_fd_sc_hd__o21a_1 _17004_ (.A1(_10005_),
    .A2(_10006_),
    .B1(_10007_),
    .X(_10014_));
 sky130_fd_sc_hd__nor2_1 _17005_ (.A(net4528),
    .B(net4727),
    .Y(_10015_));
 sky130_fd_sc_hd__nand2_1 _17006_ (.A(net4528),
    .B(net4727),
    .Y(_10016_));
 sky130_fd_sc_hd__or2b_1 _17007_ (.A(_10015_),
    .B_N(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__nor2_1 _17008_ (.A(_10014_),
    .B(_10017_),
    .Y(_10018_));
 sky130_fd_sc_hd__buf_4 _17009_ (.A(_06204_),
    .X(_10019_));
 sky130_fd_sc_hd__a21o_1 _17010_ (.A1(_10014_),
    .A2(_10017_),
    .B1(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__nand2_1 _17011_ (.A(_10010_),
    .B(_09284_),
    .Y(_10021_));
 sky130_fd_sc_hd__o21ai_1 _17012_ (.A1(_10018_),
    .A2(_10020_),
    .B1(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__mux2_1 _17013_ (.A0(_10022_),
    .A1(net4528),
    .S(_09966_),
    .X(_10023_));
 sky130_fd_sc_hd__clkbuf_1 _17014_ (.A(_10023_),
    .X(_00531_));
 sky130_fd_sc_hd__or2_1 _17015_ (.A(net4597),
    .B(net4370),
    .X(_10024_));
 sky130_fd_sc_hd__nand2_1 _17016_ (.A(net4597),
    .B(net4370),
    .Y(_10025_));
 sky130_fd_sc_hd__o21ai_2 _17017_ (.A1(_10014_),
    .A2(_10015_),
    .B1(_10016_),
    .Y(_10026_));
 sky130_fd_sc_hd__a21oi_1 _17018_ (.A1(_10024_),
    .A2(_10025_),
    .B1(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__a31o_1 _17019_ (.A1(_10026_),
    .A2(_10024_),
    .A3(_10025_),
    .B1(_06205_),
    .X(_10028_));
 sky130_fd_sc_hd__nand2_1 _17020_ (.A(_10019_),
    .B(_09281_),
    .Y(_10029_));
 sky130_fd_sc_hd__o21ai_1 _17021_ (.A1(net7796),
    .A2(_10028_),
    .B1(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__mux2_1 _17022_ (.A0(_10030_),
    .A1(net4597),
    .S(_09966_),
    .X(_10031_));
 sky130_fd_sc_hd__clkbuf_1 _17023_ (.A(_10031_),
    .X(_00532_));
 sky130_fd_sc_hd__a21boi_2 _17024_ (.A1(_10026_),
    .A2(_10024_),
    .B1_N(_10025_),
    .Y(_10032_));
 sky130_fd_sc_hd__nor2_1 _17025_ (.A(net4556),
    .B(net4719),
    .Y(_10033_));
 sky130_fd_sc_hd__nand2_1 _17026_ (.A(net4556),
    .B(net4719),
    .Y(_10034_));
 sky130_fd_sc_hd__or2b_1 _17027_ (.A(_10033_),
    .B_N(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__xnor2_1 _17028_ (.A(_10032_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__nand2_1 _17029_ (.A(_10019_),
    .B(_09276_),
    .Y(_10037_));
 sky130_fd_sc_hd__o21ai_1 _17030_ (.A1(_06206_),
    .A2(_10036_),
    .B1(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__clkbuf_1 _17031_ (.A(net4902),
    .X(_10039_));
 sky130_fd_sc_hd__mux2_1 _17032_ (.A0(_10038_),
    .A1(net4556),
    .S(net4903),
    .X(_10040_));
 sky130_fd_sc_hd__clkbuf_1 _17033_ (.A(_10040_),
    .X(_00533_));
 sky130_fd_sc_hd__o21a_1 _17034_ (.A1(_10032_),
    .A2(_10033_),
    .B1(_10034_),
    .X(_10041_));
 sky130_fd_sc_hd__nor2_1 _17035_ (.A(net4560),
    .B(net4399),
    .Y(_10042_));
 sky130_fd_sc_hd__nand2_1 _17036_ (.A(net4560),
    .B(net4399),
    .Y(_10043_));
 sky130_fd_sc_hd__or2b_1 _17037_ (.A(_10042_),
    .B_N(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__nor2_1 _17038_ (.A(_10041_),
    .B(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__a21o_1 _17039_ (.A1(_10041_),
    .A2(_10044_),
    .B1(_10019_),
    .X(_10046_));
 sky130_fd_sc_hd__nand2_1 _17040_ (.A(_10019_),
    .B(_09403_),
    .Y(_10047_));
 sky130_fd_sc_hd__o21ai_1 _17041_ (.A1(_10045_),
    .A2(_10046_),
    .B1(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__mux2_1 _17042_ (.A0(_10048_),
    .A1(net4560),
    .S(net4903),
    .X(_10049_));
 sky130_fd_sc_hd__clkbuf_1 _17043_ (.A(_10049_),
    .X(_00534_));
 sky130_fd_sc_hd__o21a_1 _17044_ (.A1(_10041_),
    .A2(_10042_),
    .B1(_10043_),
    .X(_10050_));
 sky130_fd_sc_hd__nor2_1 _17045_ (.A(net3462),
    .B(net4716),
    .Y(_10051_));
 sky130_fd_sc_hd__nand2_1 _17046_ (.A(net3462),
    .B(net4716),
    .Y(_10052_));
 sky130_fd_sc_hd__or2b_1 _17047_ (.A(_10051_),
    .B_N(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__xnor2_1 _17048_ (.A(_10050_),
    .B(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__nand2_1 _17049_ (.A(_10019_),
    .B(_09521_),
    .Y(_10055_));
 sky130_fd_sc_hd__o21ai_1 _17050_ (.A1(_06206_),
    .A2(net7596),
    .B1(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__mux2_1 _17051_ (.A0(_10056_),
    .A1(net3462),
    .S(net4903),
    .X(_10057_));
 sky130_fd_sc_hd__clkbuf_1 _17052_ (.A(_10057_),
    .X(_00535_));
 sky130_fd_sc_hd__o21a_1 _17053_ (.A1(_10050_),
    .A2(_10051_),
    .B1(_10052_),
    .X(_10058_));
 sky130_fd_sc_hd__nor2_1 _17054_ (.A(net3795),
    .B(net3419),
    .Y(_10059_));
 sky130_fd_sc_hd__nand2_1 _17055_ (.A(net3795),
    .B(net3419),
    .Y(_10060_));
 sky130_fd_sc_hd__or2b_1 _17056_ (.A(_10059_),
    .B_N(net3398),
    .X(_10061_));
 sky130_fd_sc_hd__nor2_1 _17057_ (.A(_10058_),
    .B(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__a21o_1 _17058_ (.A1(_10058_),
    .A2(_10061_),
    .B1(_10019_),
    .X(_10063_));
 sky130_fd_sc_hd__or2_1 _17059_ (.A(_09999_),
    .B(_09641_),
    .X(_10064_));
 sky130_fd_sc_hd__o21ai_1 _17060_ (.A1(_10062_),
    .A2(_10063_),
    .B1(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__mux2_1 _17061_ (.A0(_10065_),
    .A1(net3795),
    .S(net4903),
    .X(_10066_));
 sky130_fd_sc_hd__clkbuf_1 _17062_ (.A(_10066_),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _17063_ (.A(net3417),
    .B(net4714),
    .X(_10067_));
 sky130_fd_sc_hd__nand2_1 _17064_ (.A(net3417),
    .B(net4714),
    .Y(_10068_));
 sky130_fd_sc_hd__o21ai_1 _17065_ (.A1(_10058_),
    .A2(_10059_),
    .B1(net3398),
    .Y(_10069_));
 sky130_fd_sc_hd__a21oi_1 _17066_ (.A1(_10067_),
    .A2(_10068_),
    .B1(net3399),
    .Y(_10070_));
 sky130_fd_sc_hd__a31o_1 _17067_ (.A1(net3399),
    .A2(_10067_),
    .A3(_10068_),
    .B1(_06205_),
    .X(_10071_));
 sky130_fd_sc_hd__nand2_1 _17068_ (.A(_10019_),
    .B(_09769_),
    .Y(_10072_));
 sky130_fd_sc_hd__o21ai_1 _17069_ (.A1(_10070_),
    .A2(_10071_),
    .B1(_10072_),
    .Y(_10073_));
 sky130_fd_sc_hd__mux2_1 _17070_ (.A0(_10073_),
    .A1(net3417),
    .S(net4903),
    .X(_10074_));
 sky130_fd_sc_hd__clkbuf_1 _17071_ (.A(_10074_),
    .X(_00537_));
 sky130_fd_sc_hd__nand2_1 _17072_ (.A(net3399),
    .B(_10067_),
    .Y(_10075_));
 sky130_fd_sc_hd__and2_1 _17073_ (.A(net4595),
    .B(net4362),
    .X(_10076_));
 sky130_fd_sc_hd__nor2_1 _17074_ (.A(net4595),
    .B(net4362),
    .Y(_10077_));
 sky130_fd_sc_hd__a211oi_1 _17075_ (.A1(_10068_),
    .A2(net3400),
    .B1(_10076_),
    .C1(_10077_),
    .Y(_10078_));
 sky130_fd_sc_hd__o211a_1 _17076_ (.A1(_10077_),
    .A2(_10076_),
    .B1(net3400),
    .C1(_10068_),
    .X(_10079_));
 sky130_fd_sc_hd__nand2_1 _17077_ (.A(_10019_),
    .B(_09908_),
    .Y(_10080_));
 sky130_fd_sc_hd__o31ai_1 _17078_ (.A1(_10010_),
    .A2(net3401),
    .A3(_10079_),
    .B1(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__mux2_1 _17079_ (.A0(_10081_),
    .A1(net4595),
    .S(net4903),
    .X(_10082_));
 sky130_fd_sc_hd__clkbuf_1 _17080_ (.A(_10082_),
    .X(_00538_));
 sky130_fd_sc_hd__or2_1 _17081_ (.A(net3578),
    .B(net4334),
    .X(_10083_));
 sky130_fd_sc_hd__nand2_1 _17082_ (.A(net3578),
    .B(net4334),
    .Y(_10084_));
 sky130_fd_sc_hd__a211o_1 _17083_ (.A1(_10083_),
    .A2(_10084_),
    .B1(_10076_),
    .C1(net3401),
    .X(_10085_));
 sky130_fd_sc_hd__o211ai_1 _17084_ (.A1(_10076_),
    .A2(net3401),
    .B1(_10083_),
    .C1(_10084_),
    .Y(_10086_));
 sky130_fd_sc_hd__o21ai_4 _17085_ (.A1(_09669_),
    .A2(_09786_),
    .B1(_09787_),
    .Y(_10087_));
 sky130_fd_sc_hd__or2b_1 _17086_ (.A(_09828_),
    .B_N(_09793_),
    .X(_10088_));
 sky130_fd_sc_hd__a21oi_1 _17087_ (.A1(_09804_),
    .A2(_09806_),
    .B1(_09802_),
    .Y(_10089_));
 sky130_fd_sc_hd__a21oi_2 _17088_ (.A1(_09826_),
    .A2(_10088_),
    .B1(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__and3_1 _17089_ (.A(_09826_),
    .B(_10088_),
    .C(_10089_),
    .X(_10091_));
 sky130_fd_sc_hd__nor2_2 _17090_ (.A(_10090_),
    .B(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__a21o_1 _17091_ (.A1(_09807_),
    .A2(_09824_),
    .B1(_09822_),
    .X(_10093_));
 sky130_fd_sc_hd__or2b_1 _17092_ (.A(_09849_),
    .B_N(_09830_),
    .X(_10094_));
 sky130_fd_sc_hd__nor2_1 _17093_ (.A(_08724_),
    .B(_09537_),
    .Y(_10095_));
 sky130_fd_sc_hd__and3_1 _17094_ (.A(_09051_),
    .B(_09662_),
    .C(_10095_),
    .X(_10096_));
 sky130_fd_sc_hd__a21oi_1 _17095_ (.A1(_09051_),
    .A2(_09662_),
    .B1(_10095_),
    .Y(_10097_));
 sky130_fd_sc_hd__nor2_1 _17096_ (.A(_10096_),
    .B(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__and2b_1 _17097_ (.A_N(_09666_),
    .B(_09133_),
    .X(_10099_));
 sky130_fd_sc_hd__xnor2_1 _17098_ (.A(_10098_),
    .B(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__o21a_1 _17099_ (.A1(_09795_),
    .A2(_09796_),
    .B1(_09798_),
    .X(_10101_));
 sky130_fd_sc_hd__nor2_1 _17100_ (.A(_10100_),
    .B(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__and2_1 _17101_ (.A(_10100_),
    .B(_10101_),
    .X(_10103_));
 sky130_fd_sc_hd__nor2_1 _17102_ (.A(_10102_),
    .B(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__and2_1 _17103_ (.A(_08310_),
    .B(net7378),
    .X(_10105_));
 sky130_fd_sc_hd__xor2_1 _17104_ (.A(_10104_),
    .B(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__o21ai_2 _17105_ (.A1(_09676_),
    .A2(_09815_),
    .B1(_09814_),
    .Y(_10107_));
 sky130_fd_sc_hd__o21ai_4 _17106_ (.A1(_09833_),
    .A2(_09836_),
    .B1(_09834_),
    .Y(_10108_));
 sky130_fd_sc_hd__or2b_1 _17107_ (.A(_09251_),
    .B_N(_08962_),
    .X(_10109_));
 sky130_fd_sc_hd__xor2_1 _17108_ (.A(_09813_),
    .B(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__nor2_1 _17109_ (.A(_09328_),
    .B(_09312_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand2_1 _17110_ (.A(_10110_),
    .B(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__or2_1 _17111_ (.A(_10110_),
    .B(_10111_),
    .X(_10113_));
 sky130_fd_sc_hd__nand2_1 _17112_ (.A(_10112_),
    .B(_10113_),
    .Y(_10114_));
 sky130_fd_sc_hd__xnor2_2 _17113_ (.A(_10108_),
    .B(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__xnor2_1 _17114_ (.A(_10107_),
    .B(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__a21oi_1 _17115_ (.A1(_09809_),
    .A2(_09819_),
    .B1(_09817_),
    .Y(_10117_));
 sky130_fd_sc_hd__nor2_1 _17116_ (.A(_10116_),
    .B(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__and2_1 _17117_ (.A(_10116_),
    .B(_10117_),
    .X(_10119_));
 sky130_fd_sc_hd__nor2_1 _17118_ (.A(_10118_),
    .B(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__xnor2_1 _17119_ (.A(_10106_),
    .B(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__a21o_1 _17120_ (.A1(_09847_),
    .A2(_10094_),
    .B1(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__nand3_1 _17121_ (.A(_09847_),
    .B(_10094_),
    .C(_10121_),
    .Y(_10123_));
 sky130_fd_sc_hd__nand2_1 _17122_ (.A(_10122_),
    .B(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__xnor2_1 _17123_ (.A(_10093_),
    .B(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__nor2_1 _17124_ (.A(_09843_),
    .B(_09844_),
    .Y(_10126_));
 sky130_fd_sc_hd__a21o_1 _17125_ (.A1(_09838_),
    .A2(_09845_),
    .B1(_10126_),
    .X(_10127_));
 sky130_fd_sc_hd__or2b_1 _17126_ (.A(_09853_),
    .B_N(_09858_),
    .X(_10128_));
 sky130_fd_sc_hd__a21bo_1 _17127_ (.A1(_09852_),
    .A2(_09859_),
    .B1_N(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__buf_2 _17128_ (.A(_09695_),
    .X(_10130_));
 sky130_fd_sc_hd__o22ai_1 _17129_ (.A1(_08317_),
    .A2(_08548_),
    .B1(_08556_),
    .B2(_08331_),
    .Y(_10131_));
 sky130_fd_sc_hd__or4_1 _17130_ (.A(_08317_),
    .B(_08331_),
    .C(_08548_),
    .D(_08556_),
    .X(_10132_));
 sky130_fd_sc_hd__nand2_1 _17131_ (.A(_10131_),
    .B(_10132_),
    .Y(_10133_));
 sky130_fd_sc_hd__or3_1 _17132_ (.A(_10130_),
    .B(_08708_),
    .C(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__o21ai_1 _17133_ (.A1(_10130_),
    .A2(_08708_),
    .B1(_10133_),
    .Y(_10135_));
 sky130_fd_sc_hd__and2_1 _17134_ (.A(_10134_),
    .B(_10135_),
    .X(_10136_));
 sky130_fd_sc_hd__nand2_1 _17135_ (.A(_09840_),
    .B(_09841_),
    .Y(_10137_));
 sky130_fd_sc_hd__or2b_1 _17136_ (.A(_09839_),
    .B_N(_09842_),
    .X(_10138_));
 sky130_fd_sc_hd__nor2_1 _17137_ (.A(_08872_),
    .B(_09216_),
    .Y(_10139_));
 sky130_fd_sc_hd__nor2_1 _17138_ (.A(_08873_),
    .B(_08582_),
    .Y(_10140_));
 sky130_fd_sc_hd__xor2_2 _17139_ (.A(_10139_),
    .B(_10140_),
    .X(_10141_));
 sky130_fd_sc_hd__nor2_1 _17140_ (.A(_08717_),
    .B(_08574_),
    .Y(_10142_));
 sky130_fd_sc_hd__xnor2_1 _17141_ (.A(_10141_),
    .B(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__a21oi_1 _17142_ (.A1(_10137_),
    .A2(_10138_),
    .B1(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__and3_1 _17143_ (.A(_10137_),
    .B(_10138_),
    .C(_10143_),
    .X(_10145_));
 sky130_fd_sc_hd__nor2_1 _17144_ (.A(_10144_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__xnor2_2 _17145_ (.A(_10136_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__xor2_2 _17146_ (.A(_10129_),
    .B(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__xnor2_2 _17147_ (.A(_10127_),
    .B(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__or2b_1 _17148_ (.A(_09854_),
    .B_N(_09857_),
    .X(_10150_));
 sky130_fd_sc_hd__o31ai_4 _17149_ (.A1(_09108_),
    .A2(_09595_),
    .A3(_09855_),
    .B1(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__and2_1 _17150_ (.A(_09732_),
    .B(_09733_),
    .X(_10152_));
 sky130_fd_sc_hd__or3_1 _17151_ (.A(_08584_),
    .B(_10152_),
    .C(_09865_),
    .X(_10153_));
 sky130_fd_sc_hd__a21bo_1 _17152_ (.A1(_09862_),
    .A2(_09867_),
    .B1_N(_10153_),
    .X(_10154_));
 sky130_fd_sc_hd__nor2_1 _17153_ (.A(_09103_),
    .B(_09483_),
    .Y(_10155_));
 sky130_fd_sc_hd__nor2_1 _17154_ (.A(_09064_),
    .B(_09364_),
    .Y(_10156_));
 sky130_fd_sc_hd__xnor2_2 _17155_ (.A(_10155_),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__nor2_1 _17156_ (.A(_08684_),
    .B(_09477_),
    .Y(_10158_));
 sky130_fd_sc_hd__xnor2_2 _17157_ (.A(_10157_),
    .B(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__xor2_2 _17158_ (.A(_10154_),
    .B(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__xor2_2 _17159_ (.A(_10151_),
    .B(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__nor2_1 _17160_ (.A(_08587_),
    .B(_09861_),
    .Y(_10162_));
 sky130_fd_sc_hd__a21o_1 _17161_ (.A1(_09863_),
    .A2(_09864_),
    .B1(_08584_),
    .X(_10163_));
 sky130_fd_sc_hd__a21oi_1 _17162_ (.A1(_09732_),
    .A2(_09733_),
    .B1(_09086_),
    .Y(_10164_));
 sky130_fd_sc_hd__xnor2_1 _17163_ (.A(_10163_),
    .B(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__xor2_1 _17164_ (.A(_10162_),
    .B(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__and2_1 _17165_ (.A(net3502),
    .B(_09304_),
    .X(_10167_));
 sky130_fd_sc_hd__a21oi_4 _17166_ (.A1(_06211_),
    .A2(_09870_),
    .B1(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand2_1 _17167_ (.A(_08632_),
    .B(_08664_),
    .Y(_10169_));
 sky130_fd_sc_hd__o211a_1 _17168_ (.A1(net4954),
    .A2(_08664_),
    .B1(_09870_),
    .C1(_10169_),
    .X(_10170_));
 sky130_fd_sc_hd__or3b_1 _17169_ (.A(_09096_),
    .B(_10168_),
    .C_N(_10170_),
    .X(_10171_));
 sky130_fd_sc_hd__a21o_1 _17170_ (.A1(_09873_),
    .A2(_09738_),
    .B1(_09305_),
    .X(_10172_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(net3565),
    .B(_09305_),
    .Y(_10173_));
 sky130_fd_sc_hd__and2_2 _17172_ (.A(_10172_),
    .B(_10173_),
    .X(_10174_));
 sky130_fd_sc_hd__o21bai_1 _17173_ (.A1(_09096_),
    .A2(_10174_),
    .B1_N(_10170_),
    .Y(_10175_));
 sky130_fd_sc_hd__a21bo_1 _17174_ (.A1(_09871_),
    .A2(_09874_),
    .B1_N(_09872_),
    .X(_10176_));
 sky130_fd_sc_hd__nand3_2 _17175_ (.A(_10171_),
    .B(_10175_),
    .C(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__a21o_1 _17176_ (.A1(_10171_),
    .A2(_10175_),
    .B1(_10176_),
    .X(_10178_));
 sky130_fd_sc_hd__nand3_1 _17177_ (.A(_10166_),
    .B(_10177_),
    .C(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__a21o_1 _17178_ (.A1(_10177_),
    .A2(_10178_),
    .B1(_10166_),
    .X(_10180_));
 sky130_fd_sc_hd__a21bo_1 _17179_ (.A1(_09868_),
    .A2(_09880_),
    .B1_N(_09879_),
    .X(_10181_));
 sky130_fd_sc_hd__nand3_1 _17180_ (.A(_10179_),
    .B(_10180_),
    .C(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__a21o_1 _17181_ (.A1(_10179_),
    .A2(_10180_),
    .B1(_10181_),
    .X(_10183_));
 sky130_fd_sc_hd__and3_1 _17182_ (.A(_10161_),
    .B(_10182_),
    .C(_10183_),
    .X(_10184_));
 sky130_fd_sc_hd__a21oi_1 _17183_ (.A1(_10182_),
    .A2(_10183_),
    .B1(_10161_),
    .Y(_10185_));
 sky130_fd_sc_hd__or2_2 _17184_ (.A(_10184_),
    .B(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__and2_2 _17185_ (.A(_09885_),
    .B(_09887_),
    .X(_10187_));
 sky130_fd_sc_hd__xor2_2 _17186_ (.A(_10186_),
    .B(_10187_),
    .X(_10188_));
 sky130_fd_sc_hd__xnor2_2 _17187_ (.A(_10149_),
    .B(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__a21boi_2 _17188_ (.A1(_09850_),
    .A2(_09892_),
    .B1_N(_09891_),
    .Y(_10190_));
 sky130_fd_sc_hd__xor2_2 _17189_ (.A(_10189_),
    .B(_10190_),
    .X(_10191_));
 sky130_fd_sc_hd__xnor2_1 _17190_ (.A(_10125_),
    .B(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__nor2_1 _17191_ (.A(_09895_),
    .B(_09896_),
    .Y(_10193_));
 sky130_fd_sc_hd__a21oi_2 _17192_ (.A1(_09829_),
    .A2(_09897_),
    .B1(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__nor2_2 _17193_ (.A(_10192_),
    .B(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__and2_1 _17194_ (.A(_10192_),
    .B(_10194_),
    .X(_10196_));
 sky130_fd_sc_hd__nor2_4 _17195_ (.A(_10195_),
    .B(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__xnor2_4 _17196_ (.A(_10092_),
    .B(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__o2bb2a_4 _17197_ (.A1_N(_09792_),
    .A2_N(_09900_),
    .B1(_09899_),
    .B2(_09898_),
    .X(_10199_));
 sky130_fd_sc_hd__xor2_4 _17198_ (.A(_10198_),
    .B(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__xor2_4 _17199_ (.A(_10087_),
    .B(_10200_),
    .X(_10201_));
 sky130_fd_sc_hd__xnor2_4 _17200_ (.A(_09904_),
    .B(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__a21o_1 _17201_ (.A1(_09782_),
    .A2(_09780_),
    .B1(_09906_),
    .X(_10203_));
 sky130_fd_sc_hd__o31a_4 _17202_ (.A1(_09652_),
    .A2(_09779_),
    .A3(_09907_),
    .B1(_10203_),
    .X(_10204_));
 sky130_fd_sc_hd__xor2_4 _17203_ (.A(_10202_),
    .B(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__and2_1 _17204_ (.A(_06204_),
    .B(_10205_),
    .X(_10206_));
 sky130_fd_sc_hd__a31o_1 _17205_ (.A1(_09987_),
    .A2(_10085_),
    .A3(net7824),
    .B1(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__mux2_1 _17206_ (.A0(_10207_),
    .A1(net3578),
    .S(net4903),
    .X(_10208_));
 sky130_fd_sc_hd__clkbuf_1 _17207_ (.A(_10208_),
    .X(_00539_));
 sky130_fd_sc_hd__and2_1 _17208_ (.A(net4540),
    .B(net4411),
    .X(_10209_));
 sky130_fd_sc_hd__nor2_1 _17209_ (.A(net4540),
    .B(net4411),
    .Y(_10210_));
 sky130_fd_sc_hd__a211o_1 _17210_ (.A1(_10084_),
    .A2(_10086_),
    .B1(_10209_),
    .C1(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__o211ai_1 _17211_ (.A1(_10209_),
    .A2(_10210_),
    .B1(_10084_),
    .C1(net7824),
    .Y(_10212_));
 sky130_fd_sc_hd__or2_1 _17212_ (.A(_10198_),
    .B(_10199_),
    .X(_10213_));
 sky130_fd_sc_hd__nand2_1 _17213_ (.A(_10087_),
    .B(_10200_),
    .Y(_10214_));
 sky130_fd_sc_hd__or2b_1 _17214_ (.A(_10124_),
    .B_N(_10093_),
    .X(_10215_));
 sky130_fd_sc_hd__a21oi_2 _17215_ (.A1(_10104_),
    .A2(_10105_),
    .B1(_10102_),
    .Y(_10216_));
 sky130_fd_sc_hd__a21oi_4 _17216_ (.A1(_10122_),
    .A2(_10215_),
    .B1(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__and3_1 _17217_ (.A(_10122_),
    .B(_10215_),
    .C(_10216_),
    .X(_10218_));
 sky130_fd_sc_hd__nor2_2 _17218_ (.A(_10217_),
    .B(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__a21o_1 _17219_ (.A1(_10106_),
    .A2(_10120_),
    .B1(_10118_),
    .X(_10220_));
 sky130_fd_sc_hd__or2b_1 _17220_ (.A(_10147_),
    .B_N(_10129_),
    .X(_10221_));
 sky130_fd_sc_hd__or2b_1 _17221_ (.A(_10148_),
    .B_N(_10127_),
    .X(_10222_));
 sky130_fd_sc_hd__nor2_1 _17222_ (.A(_09328_),
    .B(_09538_),
    .Y(_10223_));
 sky130_fd_sc_hd__inv_2 _17223_ (.A(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__a2bb2o_1 _17224_ (.A1_N(_09328_),
    .A2_N(_09419_),
    .B1(_09794_),
    .B2(_09051_),
    .X(_10225_));
 sky130_fd_sc_hd__o21a_1 _17225_ (.A1(_09797_),
    .A2(_10224_),
    .B1(_10225_),
    .X(_10226_));
 sky130_fd_sc_hd__nor2_1 _17226_ (.A(_08724_),
    .B(_09666_),
    .Y(_10227_));
 sky130_fd_sc_hd__xnor2_1 _17227_ (.A(_10226_),
    .B(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__a21oi_1 _17228_ (.A1(_10098_),
    .A2(_10099_),
    .B1(_10096_),
    .Y(_10229_));
 sky130_fd_sc_hd__nor2_1 _17229_ (.A(_10228_),
    .B(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__and2_1 _17230_ (.A(_10228_),
    .B(_10229_),
    .X(_10231_));
 sky130_fd_sc_hd__nor2_1 _17231_ (.A(_10230_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__nor2_1 _17232_ (.A(_09133_),
    .B(_09784_),
    .Y(_10233_));
 sky130_fd_sc_hd__xor2_1 _17233_ (.A(_10232_),
    .B(_10233_),
    .X(_10234_));
 sky130_fd_sc_hd__o21ai_1 _17234_ (.A1(_09813_),
    .A2(_10109_),
    .B1(_10112_),
    .Y(_10235_));
 sky130_fd_sc_hd__or2_1 _17235_ (.A(_10130_),
    .B(_09251_),
    .X(_10236_));
 sky130_fd_sc_hd__a2bb2o_1 _17236_ (.A1_N(_09251_),
    .A2_N(_09562_),
    .B1(_08849_),
    .B2(_09306_),
    .X(_10237_));
 sky130_fd_sc_hd__o21a_1 _17237_ (.A1(_09813_),
    .A2(_10236_),
    .B1(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__and2b_1 _17238_ (.A_N(_09311_),
    .B(_09447_),
    .X(_10239_));
 sky130_fd_sc_hd__xnor2_1 _17239_ (.A(_10238_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__a21oi_1 _17240_ (.A1(_10132_),
    .A2(_10134_),
    .B1(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__and3_1 _17241_ (.A(_10132_),
    .B(_10134_),
    .C(_10240_),
    .X(_10242_));
 sky130_fd_sc_hd__nor2_1 _17242_ (.A(_10241_),
    .B(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__xnor2_1 _17243_ (.A(_10235_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__a32oi_4 _17244_ (.A1(_10108_),
    .A2(_10112_),
    .A3(_10113_),
    .B1(_10115_),
    .B2(_10107_),
    .Y(_10245_));
 sky130_fd_sc_hd__nor2_1 _17245_ (.A(_10244_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__and2_1 _17246_ (.A(_10244_),
    .B(_10245_),
    .X(_10247_));
 sky130_fd_sc_hd__nor2_1 _17247_ (.A(_10246_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__xnor2_1 _17248_ (.A(_10234_),
    .B(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__a21o_1 _17249_ (.A1(_10221_),
    .A2(_10222_),
    .B1(_10249_),
    .X(_10250_));
 sky130_fd_sc_hd__nand3_1 _17250_ (.A(_10221_),
    .B(_10222_),
    .C(_10249_),
    .Y(_10251_));
 sky130_fd_sc_hd__nand2_1 _17251_ (.A(_10250_),
    .B(_10251_),
    .Y(_10252_));
 sky130_fd_sc_hd__xnor2_2 _17252_ (.A(_10220_),
    .B(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__a21o_1 _17253_ (.A1(_10136_),
    .A2(_10146_),
    .B1(_10144_),
    .X(_10254_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(_10154_),
    .B(_10159_),
    .Y(_10255_));
 sky130_fd_sc_hd__nand2_1 _17255_ (.A(_10151_),
    .B(_10160_),
    .Y(_10256_));
 sky130_fd_sc_hd__buf_2 _17256_ (.A(_08556_),
    .X(_10257_));
 sky130_fd_sc_hd__or4_2 _17257_ (.A(_08315_),
    .B(_08331_),
    .C(_08641_),
    .D(_08548_),
    .X(_10258_));
 sky130_fd_sc_hd__buf_2 _17258_ (.A(_08315_),
    .X(_10259_));
 sky130_fd_sc_hd__a2bb2o_1 _17259_ (.A1_N(_10259_),
    .A2_N(_08641_),
    .B1(_08754_),
    .B2(_08701_),
    .X(_10260_));
 sky130_fd_sc_hd__nand2_1 _17260_ (.A(_10258_),
    .B(_10260_),
    .Y(_10261_));
 sky130_fd_sc_hd__or3_1 _17261_ (.A(_10257_),
    .B(_08708_),
    .C(_10261_),
    .X(_10262_));
 sky130_fd_sc_hd__o21ai_1 _17262_ (.A1(_10257_),
    .A2(_08708_),
    .B1(_10261_),
    .Y(_10263_));
 sky130_fd_sc_hd__and2_1 _17263_ (.A(_10262_),
    .B(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__nor2_1 _17264_ (.A(_08873_),
    .B(_09216_),
    .Y(_10265_));
 sky130_fd_sc_hd__nor2_1 _17265_ (.A(_08872_),
    .B(_09477_),
    .Y(_10266_));
 sky130_fd_sc_hd__xor2_1 _17266_ (.A(_10265_),
    .B(_10266_),
    .X(_10267_));
 sky130_fd_sc_hd__nor2_1 _17267_ (.A(_08717_),
    .B(_08582_),
    .Y(_10268_));
 sky130_fd_sc_hd__xnor2_1 _17268_ (.A(_10267_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__nand2_1 _17269_ (.A(_10139_),
    .B(_10140_),
    .Y(_10270_));
 sky130_fd_sc_hd__a21boi_2 _17270_ (.A1(_10141_),
    .A2(_10142_),
    .B1_N(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__nor2_1 _17271_ (.A(_10269_),
    .B(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__nand2_1 _17272_ (.A(_10269_),
    .B(_10271_),
    .Y(_10273_));
 sky130_fd_sc_hd__and2b_1 _17273_ (.A_N(_10272_),
    .B(_10273_),
    .X(_10274_));
 sky130_fd_sc_hd__xnor2_1 _17274_ (.A(_10264_),
    .B(_10274_),
    .Y(_10275_));
 sky130_fd_sc_hd__a21o_1 _17275_ (.A1(_10255_),
    .A2(_10256_),
    .B1(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__nand3_1 _17276_ (.A(_10255_),
    .B(_10256_),
    .C(_10275_),
    .Y(_10277_));
 sky130_fd_sc_hd__nand2_1 _17277_ (.A(_10276_),
    .B(_10277_),
    .Y(_10278_));
 sky130_fd_sc_hd__xnor2_2 _17278_ (.A(_10254_),
    .B(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__or3_1 _17279_ (.A(_09582_),
    .B(_09477_),
    .C(_10157_),
    .X(_10280_));
 sky130_fd_sc_hd__a21bo_1 _17280_ (.A1(_10155_),
    .A2(_10156_),
    .B1_N(_10280_),
    .X(_10281_));
 sky130_fd_sc_hd__or3_1 _17281_ (.A(_09139_),
    .B(_10152_),
    .C(_10163_),
    .X(_10282_));
 sky130_fd_sc_hd__a21bo_1 _17282_ (.A1(_10162_),
    .A2(_10165_),
    .B1_N(_10282_),
    .X(_10283_));
 sky130_fd_sc_hd__or4_1 _17283_ (.A(_09103_),
    .B(_09064_),
    .C(_09483_),
    .D(_09603_),
    .X(_10284_));
 sky130_fd_sc_hd__o22ai_1 _17284_ (.A1(_09064_),
    .A2(_09484_),
    .B1(_09603_),
    .B2(_09103_),
    .Y(_10285_));
 sky130_fd_sc_hd__nand2_1 _17285_ (.A(_10284_),
    .B(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__nor2_1 _17286_ (.A(_08684_),
    .B(_09595_),
    .Y(_10287_));
 sky130_fd_sc_hd__xnor2_1 _17287_ (.A(_10286_),
    .B(_10287_),
    .Y(_10288_));
 sky130_fd_sc_hd__xor2_1 _17288_ (.A(_10283_),
    .B(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(_10281_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__or2_1 _17290_ (.A(_10281_),
    .B(_10289_),
    .X(_10291_));
 sky130_fd_sc_hd__and2_1 _17291_ (.A(_10290_),
    .B(_10291_),
    .X(_10292_));
 sky130_fd_sc_hd__nor2_1 _17292_ (.A(_09593_),
    .B(_10152_),
    .Y(_10293_));
 sky130_fd_sc_hd__a21o_1 _17293_ (.A1(_09863_),
    .A2(_09864_),
    .B1(_09086_),
    .X(_10294_));
 sky130_fd_sc_hd__a21oi_1 _17294_ (.A1(_10172_),
    .A2(_10173_),
    .B1(_08584_),
    .Y(_10295_));
 sky130_fd_sc_hd__xnor2_1 _17295_ (.A(_10294_),
    .B(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__xor2_1 _17296_ (.A(_10293_),
    .B(_10296_),
    .X(_10297_));
 sky130_fd_sc_hd__and2_1 _17297_ (.A(_09870_),
    .B(_10169_),
    .X(_10298_));
 sky130_fd_sc_hd__nor2_1 _17298_ (.A(_09096_),
    .B(_10168_),
    .Y(_10299_));
 sky130_fd_sc_hd__nand2_1 _17299_ (.A(_08755_),
    .B(_09870_),
    .Y(_10300_));
 sky130_fd_sc_hd__or4_4 _17300_ (.A(_09096_),
    .B(net4954),
    .C(_10300_),
    .D(_10168_),
    .X(_10301_));
 sky130_fd_sc_hd__o21a_2 _17301_ (.A1(_10298_),
    .A2(_10299_),
    .B1(_10301_),
    .X(_10302_));
 sky130_fd_sc_hd__xnor2_1 _17302_ (.A(_10297_),
    .B(_10302_),
    .Y(_10303_));
 sky130_fd_sc_hd__a21oi_1 _17303_ (.A1(_10177_),
    .A2(_10179_),
    .B1(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__and3_1 _17304_ (.A(_10177_),
    .B(_10179_),
    .C(_10303_),
    .X(_10305_));
 sky130_fd_sc_hd__nor2_1 _17305_ (.A(_10304_),
    .B(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__xnor2_2 _17306_ (.A(_10292_),
    .B(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__a21boi_2 _17307_ (.A1(_10161_),
    .A2(_10183_),
    .B1_N(_10182_),
    .Y(_10308_));
 sky130_fd_sc_hd__xor2_2 _17308_ (.A(_10307_),
    .B(_10308_),
    .X(_10309_));
 sky130_fd_sc_hd__xnor2_1 _17309_ (.A(_10279_),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__nor2_1 _17310_ (.A(_10186_),
    .B(_10187_),
    .Y(_10311_));
 sky130_fd_sc_hd__a21oi_2 _17311_ (.A1(_10149_),
    .A2(_10188_),
    .B1(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__nor2_1 _17312_ (.A(_10310_),
    .B(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand2_1 _17313_ (.A(_10310_),
    .B(_10312_),
    .Y(_10314_));
 sky130_fd_sc_hd__and2b_1 _17314_ (.A_N(_10314_),
    .B(_10313_),
    .X(_10315_));
 sky130_fd_sc_hd__xnor2_2 _17315_ (.A(_10253_),
    .B(_10315_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_1 _17316_ (.A(_10189_),
    .B(_10190_),
    .Y(_10317_));
 sky130_fd_sc_hd__a21oi_2 _17317_ (.A1(_10125_),
    .A2(_10191_),
    .B1(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__xor2_2 _17318_ (.A(_10316_),
    .B(_10318_),
    .X(_10319_));
 sky130_fd_sc_hd__xnor2_2 _17319_ (.A(_10219_),
    .B(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__a21oi_2 _17320_ (.A1(_10092_),
    .A2(_10197_),
    .B1(_10195_),
    .Y(_10321_));
 sky130_fd_sc_hd__xor2_2 _17321_ (.A(_10320_),
    .B(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__xnor2_2 _17322_ (.A(_10090_),
    .B(_10322_),
    .Y(_10323_));
 sky130_fd_sc_hd__a21oi_1 _17323_ (.A1(_10213_),
    .A2(_10214_),
    .B1(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__and3_1 _17324_ (.A(_10213_),
    .B(_10214_),
    .C(_10323_),
    .X(_10325_));
 sky130_fd_sc_hd__nor2_2 _17325_ (.A(_10324_),
    .B(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__nand2_1 _17326_ (.A(_09904_),
    .B(_10201_),
    .Y(_10327_));
 sky130_fd_sc_hd__o21ai_2 _17327_ (.A1(_10202_),
    .A2(_10204_),
    .B1(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__xor2_4 _17328_ (.A(_10326_),
    .B(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__and2_1 _17329_ (.A(_06204_),
    .B(_10329_),
    .X(_10330_));
 sky130_fd_sc_hd__a31o_1 _17330_ (.A1(_09987_),
    .A2(_10211_),
    .A3(_10212_),
    .B1(_10330_),
    .X(_10331_));
 sky130_fd_sc_hd__mux2_1 _17331_ (.A0(_10331_),
    .A1(net4540),
    .S(net4903),
    .X(_10332_));
 sky130_fd_sc_hd__clkbuf_1 _17332_ (.A(_10332_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _17333_ (.A(net3474),
    .B(net4349),
    .Y(_10333_));
 sky130_fd_sc_hd__or2_1 _17334_ (.A(net3474),
    .B(net4349),
    .X(_10334_));
 sky130_fd_sc_hd__inv_2 _17335_ (.A(_10211_),
    .Y(_10335_));
 sky130_fd_sc_hd__a211o_1 _17336_ (.A1(_10333_),
    .A2(_10334_),
    .B1(_10209_),
    .C1(_10335_),
    .X(_10336_));
 sky130_fd_sc_hd__o211ai_2 _17337_ (.A1(_10209_),
    .A2(_10335_),
    .B1(_10333_),
    .C1(_10334_),
    .Y(_10337_));
 sky130_fd_sc_hd__or2b_1 _17338_ (.A(_10252_),
    .B_N(_10220_),
    .X(_10338_));
 sky130_fd_sc_hd__a21oi_1 _17339_ (.A1(_10232_),
    .A2(_10233_),
    .B1(_10230_),
    .Y(_10339_));
 sky130_fd_sc_hd__a21oi_2 _17340_ (.A1(_10250_),
    .A2(_10338_),
    .B1(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__and3_1 _17341_ (.A(_10250_),
    .B(_10338_),
    .C(_10339_),
    .X(_10341_));
 sky130_fd_sc_hd__nor2_2 _17342_ (.A(_10340_),
    .B(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__a21o_1 _17343_ (.A1(_10234_),
    .A2(_10248_),
    .B1(_10246_),
    .X(_10343_));
 sky130_fd_sc_hd__or2b_1 _17344_ (.A(_10278_),
    .B_N(_10254_),
    .X(_10344_));
 sky130_fd_sc_hd__a21oi_1 _17345_ (.A1(_09447_),
    .A2(_09662_),
    .B1(_10223_),
    .Y(_10345_));
 sky130_fd_sc_hd__or4bb_1 _17346_ (.A(_09538_),
    .B(_09328_),
    .C_N(_09447_),
    .D_N(_09662_),
    .X(_10346_));
 sky130_fd_sc_hd__and2b_1 _17347_ (.A_N(_10345_),
    .B(_10346_),
    .X(_10347_));
 sky130_fd_sc_hd__nor2_1 _17348_ (.A(_09091_),
    .B(_09666_),
    .Y(_10348_));
 sky130_fd_sc_hd__xnor2_1 _17349_ (.A(_10347_),
    .B(_10348_),
    .Y(_10349_));
 sky130_fd_sc_hd__o2bb2a_1 _17350_ (.A1_N(_10225_),
    .A2_N(_10227_),
    .B1(_10224_),
    .B2(_09797_),
    .X(_10350_));
 sky130_fd_sc_hd__nor2_1 _17351_ (.A(_10349_),
    .B(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__and2_1 _17352_ (.A(_10349_),
    .B(_10350_),
    .X(_10352_));
 sky130_fd_sc_hd__nor2_1 _17353_ (.A(_10351_),
    .B(_10352_),
    .Y(_10353_));
 sky130_fd_sc_hd__and2_1 _17354_ (.A(_08724_),
    .B(net7378),
    .X(_10354_));
 sky130_fd_sc_hd__xor2_1 _17355_ (.A(_10353_),
    .B(_10354_),
    .X(_10355_));
 sky130_fd_sc_hd__a2bb2o_1 _17356_ (.A1_N(_09813_),
    .A2_N(_10236_),
    .B1(_10239_),
    .B2(_10237_),
    .X(_10356_));
 sky130_fd_sc_hd__or2_1 _17357_ (.A(_08556_),
    .B(_08795_),
    .X(_10357_));
 sky130_fd_sc_hd__nor2_1 _17358_ (.A(_08556_),
    .B(_09251_),
    .Y(_10358_));
 sky130_fd_sc_hd__and3_1 _17359_ (.A(_08849_),
    .B(_09306_),
    .C(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__a21oi_1 _17360_ (.A1(_10236_),
    .A2(_10357_),
    .B1(_10359_),
    .Y(_10360_));
 sky130_fd_sc_hd__nor2_1 _17361_ (.A(_09562_),
    .B(_09312_),
    .Y(_10361_));
 sky130_fd_sc_hd__xnor2_1 _17362_ (.A(_10360_),
    .B(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__a21oi_1 _17363_ (.A1(_10258_),
    .A2(_10262_),
    .B1(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__and3_1 _17364_ (.A(_10258_),
    .B(_10262_),
    .C(_10362_),
    .X(_10364_));
 sky130_fd_sc_hd__nor2_1 _17365_ (.A(_10363_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__xnor2_1 _17366_ (.A(_10356_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__a21oi_1 _17367_ (.A1(_10235_),
    .A2(_10243_),
    .B1(_10241_),
    .Y(_10367_));
 sky130_fd_sc_hd__nor2_1 _17368_ (.A(_10366_),
    .B(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__and2_1 _17369_ (.A(_10366_),
    .B(_10367_),
    .X(_10369_));
 sky130_fd_sc_hd__nor2_1 _17370_ (.A(_10368_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__xnor2_1 _17371_ (.A(_10355_),
    .B(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a21o_1 _17372_ (.A1(_10276_),
    .A2(_10344_),
    .B1(_10371_),
    .X(_10372_));
 sky130_fd_sc_hd__nand3_1 _17373_ (.A(_10276_),
    .B(_10344_),
    .C(_10371_),
    .Y(_10373_));
 sky130_fd_sc_hd__nand2_1 _17374_ (.A(_10372_),
    .B(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__xnor2_2 _17375_ (.A(_10343_),
    .B(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__a21o_1 _17376_ (.A1(_10264_),
    .A2(_10273_),
    .B1(_10272_),
    .X(_10376_));
 sky130_fd_sc_hd__nand2_1 _17377_ (.A(_10283_),
    .B(_10288_),
    .Y(_10377_));
 sky130_fd_sc_hd__o2bb2a_1 _17378_ (.A1_N(_08701_),
    .A2_N(_08540_),
    .B1(_08643_),
    .B2(_08317_),
    .X(_10378_));
 sky130_fd_sc_hd__buf_2 _17379_ (.A(_08641_),
    .X(_10379_));
 sky130_fd_sc_hd__nand2_2 _17380_ (.A(_08579_),
    .B(_08580_),
    .Y(_10380_));
 sky130_fd_sc_hd__or4_1 _17381_ (.A(_10259_),
    .B(_08329_),
    .C(_10379_),
    .D(_10380_),
    .X(_10381_));
 sky130_fd_sc_hd__or2b_1 _17382_ (.A(_10378_),
    .B_N(_10381_),
    .X(_10382_));
 sky130_fd_sc_hd__clkbuf_4 _17383_ (.A(_08548_),
    .X(_10383_));
 sky130_fd_sc_hd__nor2_1 _17384_ (.A(_10383_),
    .B(_08708_),
    .Y(_10384_));
 sky130_fd_sc_hd__xnor2_2 _17385_ (.A(_10382_),
    .B(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__nor2_1 _17386_ (.A(_08873_),
    .B(_09477_),
    .Y(_10386_));
 sky130_fd_sc_hd__or2_1 _17387_ (.A(_08872_),
    .B(_09595_),
    .X(_10387_));
 sky130_fd_sc_hd__xnor2_1 _17388_ (.A(_10386_),
    .B(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__nor2_1 _17389_ (.A(_08717_),
    .B(_09216_),
    .Y(_10389_));
 sky130_fd_sc_hd__nand2_1 _17390_ (.A(_10388_),
    .B(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__or2_1 _17391_ (.A(_10388_),
    .B(_10389_),
    .X(_10391_));
 sky130_fd_sc_hd__nand2_1 _17392_ (.A(_10390_),
    .B(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__and2_1 _17393_ (.A(_10267_),
    .B(_10268_),
    .X(_10393_));
 sky130_fd_sc_hd__a21oi_1 _17394_ (.A1(_10265_),
    .A2(_10266_),
    .B1(_10393_),
    .Y(_10394_));
 sky130_fd_sc_hd__nor2_1 _17395_ (.A(_10392_),
    .B(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__and2_1 _17396_ (.A(_10392_),
    .B(_10394_),
    .X(_10396_));
 sky130_fd_sc_hd__nor2_1 _17397_ (.A(_10395_),
    .B(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__xnor2_1 _17398_ (.A(_10385_),
    .B(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__a21o_1 _17399_ (.A1(_10377_),
    .A2(_10290_),
    .B1(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__nand3_1 _17400_ (.A(_10377_),
    .B(_10290_),
    .C(_10398_),
    .Y(_10400_));
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(_10399_),
    .B(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__xnor2_2 _17402_ (.A(_10376_),
    .B(_10401_),
    .Y(_10402_));
 sky130_fd_sc_hd__a21bo_1 _17403_ (.A1(_10285_),
    .A2(_10287_),
    .B1_N(_10284_),
    .X(_10403_));
 sky130_fd_sc_hd__or3_1 _17404_ (.A(_09138_),
    .B(_10174_),
    .C(_10294_),
    .X(_10404_));
 sky130_fd_sc_hd__a21bo_1 _17405_ (.A1(_10293_),
    .A2(_10296_),
    .B1_N(_10404_),
    .X(_10405_));
 sky130_fd_sc_hd__buf_2 _17406_ (.A(_09064_),
    .X(_10406_));
 sky130_fd_sc_hd__clkbuf_4 _17407_ (.A(_10152_),
    .X(_10407_));
 sky130_fd_sc_hd__or4_1 _17408_ (.A(_09103_),
    .B(_10406_),
    .C(_09861_),
    .D(_10407_),
    .X(_10408_));
 sky130_fd_sc_hd__o22ai_1 _17409_ (.A1(_10406_),
    .A2(_09861_),
    .B1(_10407_),
    .B2(_09108_),
    .Y(_10409_));
 sky130_fd_sc_hd__nand2_1 _17410_ (.A(_10408_),
    .B(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__nor2_1 _17411_ (.A(_09582_),
    .B(_09484_),
    .Y(_10411_));
 sky130_fd_sc_hd__xnor2_1 _17412_ (.A(_10410_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__xnor2_1 _17413_ (.A(_10405_),
    .B(_10412_),
    .Y(_10413_));
 sky130_fd_sc_hd__xnor2_1 _17414_ (.A(_10403_),
    .B(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__and2_1 _17415_ (.A(_09863_),
    .B(_09864_),
    .X(_10415_));
 sky130_fd_sc_hd__clkbuf_4 _17416_ (.A(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__nor2_1 _17417_ (.A(_09593_),
    .B(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__o22ai_1 _17418_ (.A1(_09138_),
    .A2(_10168_),
    .B1(_10174_),
    .B2(_09139_),
    .Y(_10418_));
 sky130_fd_sc_hd__or4_1 _17419_ (.A(_09138_),
    .B(_09139_),
    .C(_10168_),
    .D(_10174_),
    .X(_10419_));
 sky130_fd_sc_hd__nand3_1 _17420_ (.A(_10417_),
    .B(_10418_),
    .C(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__a21o_1 _17421_ (.A1(_10418_),
    .A2(_10419_),
    .B1(_10417_),
    .X(_10421_));
 sky130_fd_sc_hd__nand3_1 _17422_ (.A(_10302_),
    .B(_10420_),
    .C(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__a21o_1 _17423_ (.A1(_10420_),
    .A2(_10421_),
    .B1(_10302_),
    .X(_10423_));
 sky130_fd_sc_hd__a21bo_1 _17424_ (.A1(_10297_),
    .A2(_10302_),
    .B1_N(_10301_),
    .X(_10424_));
 sky130_fd_sc_hd__nand3_1 _17425_ (.A(_10422_),
    .B(_10423_),
    .C(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__a21o_1 _17426_ (.A1(_10422_),
    .A2(_10423_),
    .B1(_10424_),
    .X(_10426_));
 sky130_fd_sc_hd__nand2_1 _17427_ (.A(_10425_),
    .B(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__xor2_1 _17428_ (.A(_10414_),
    .B(_10427_),
    .X(_10428_));
 sky130_fd_sc_hd__a21oi_1 _17429_ (.A1(_10292_),
    .A2(_10306_),
    .B1(_10304_),
    .Y(_10429_));
 sky130_fd_sc_hd__nor2_1 _17430_ (.A(_10428_),
    .B(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__and2_1 _17431_ (.A(_10428_),
    .B(_10429_),
    .X(_10431_));
 sky130_fd_sc_hd__nor2_1 _17432_ (.A(_10430_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__xnor2_2 _17433_ (.A(_10402_),
    .B(_10432_),
    .Y(_10433_));
 sky130_fd_sc_hd__nor2_1 _17434_ (.A(_10307_),
    .B(_10308_),
    .Y(_10434_));
 sky130_fd_sc_hd__a21oi_2 _17435_ (.A1(_10279_),
    .A2(_10309_),
    .B1(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__xor2_2 _17436_ (.A(_10433_),
    .B(_10435_),
    .X(_10436_));
 sky130_fd_sc_hd__xnor2_1 _17437_ (.A(_10375_),
    .B(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__a21oi_1 _17438_ (.A1(_10253_),
    .A2(_10314_),
    .B1(_10313_),
    .Y(_10438_));
 sky130_fd_sc_hd__nor2_1 _17439_ (.A(_10437_),
    .B(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__nand2_1 _17440_ (.A(_10437_),
    .B(_10438_),
    .Y(_10440_));
 sky130_fd_sc_hd__and2b_1 _17441_ (.A_N(_10439_),
    .B(_10440_),
    .X(_10441_));
 sky130_fd_sc_hd__xnor2_4 _17442_ (.A(_10342_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__nor2_1 _17443_ (.A(_10316_),
    .B(_10318_),
    .Y(_10443_));
 sky130_fd_sc_hd__a21oi_2 _17444_ (.A1(_10219_),
    .A2(_10319_),
    .B1(_10443_),
    .Y(_10444_));
 sky130_fd_sc_hd__xor2_4 _17445_ (.A(_10442_),
    .B(_10444_),
    .X(_10445_));
 sky130_fd_sc_hd__xnor2_4 _17446_ (.A(_10217_),
    .B(_10445_),
    .Y(_10446_));
 sky130_fd_sc_hd__nor2_1 _17447_ (.A(_10320_),
    .B(_10321_),
    .Y(_10447_));
 sky130_fd_sc_hd__a21oi_2 _17448_ (.A1(_10090_),
    .A2(_10322_),
    .B1(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__xor2_4 _17449_ (.A(_10446_),
    .B(_10448_),
    .X(_10449_));
 sky130_fd_sc_hd__a21o_1 _17450_ (.A1(_10213_),
    .A2(_10214_),
    .B1(_10323_),
    .X(_10450_));
 sky130_fd_sc_hd__or3b_1 _17451_ (.A(_10325_),
    .B(_10202_),
    .C_N(_10450_),
    .X(_10451_));
 sky130_fd_sc_hd__a21o_1 _17452_ (.A1(_10327_),
    .A2(_10450_),
    .B1(_10325_),
    .X(_10452_));
 sky130_fd_sc_hd__o21a_4 _17453_ (.A1(_10204_),
    .A2(_10451_),
    .B1(_10452_),
    .X(_10453_));
 sky130_fd_sc_hd__xnor2_4 _17454_ (.A(_10449_),
    .B(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__and2_1 _17455_ (.A(_06204_),
    .B(_10454_),
    .X(_10455_));
 sky130_fd_sc_hd__a31o_1 _17456_ (.A1(_09987_),
    .A2(_10336_),
    .A3(_10337_),
    .B1(_10455_),
    .X(_10456_));
 sky130_fd_sc_hd__mux2_1 _17457_ (.A0(_10456_),
    .A1(net3474),
    .S(net4903),
    .X(_10457_));
 sky130_fd_sc_hd__clkbuf_1 _17458_ (.A(_10457_),
    .X(_00541_));
 sky130_fd_sc_hd__and2_1 _17459_ (.A(net4501),
    .B(net4417),
    .X(_10458_));
 sky130_fd_sc_hd__nor2_1 _17460_ (.A(net4501),
    .B(net4417),
    .Y(_10459_));
 sky130_fd_sc_hd__a211oi_1 _17461_ (.A1(_10333_),
    .A2(_10337_),
    .B1(_10458_),
    .C1(_10459_),
    .Y(_10460_));
 sky130_fd_sc_hd__o211a_1 _17462_ (.A1(_10458_),
    .A2(_10459_),
    .B1(_10333_),
    .C1(_10337_),
    .X(_10461_));
 sky130_fd_sc_hd__or2_1 _17463_ (.A(_10446_),
    .B(_10448_),
    .X(_10462_));
 sky130_fd_sc_hd__inv_2 _17464_ (.A(_10449_),
    .Y(_10463_));
 sky130_fd_sc_hd__or2_1 _17465_ (.A(_10463_),
    .B(_10453_),
    .X(_10464_));
 sky130_fd_sc_hd__or2_1 _17466_ (.A(_10442_),
    .B(_10444_),
    .X(_10465_));
 sky130_fd_sc_hd__nand2_1 _17467_ (.A(_10217_),
    .B(_10445_),
    .Y(_10466_));
 sky130_fd_sc_hd__or2b_1 _17468_ (.A(_10374_),
    .B_N(_10343_),
    .X(_10467_));
 sky130_fd_sc_hd__a21oi_1 _17469_ (.A1(_10353_),
    .A2(_10354_),
    .B1(_10351_),
    .Y(_10468_));
 sky130_fd_sc_hd__a21oi_2 _17470_ (.A1(_10372_),
    .A2(_10467_),
    .B1(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__and3_1 _17471_ (.A(_10372_),
    .B(_10467_),
    .C(_10468_),
    .X(_10470_));
 sky130_fd_sc_hd__nor2_1 _17472_ (.A(_10469_),
    .B(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__a21o_1 _17473_ (.A1(_10355_),
    .A2(_10370_),
    .B1(_10368_),
    .X(_10472_));
 sky130_fd_sc_hd__or2b_1 _17474_ (.A(_10401_),
    .B_N(_10376_),
    .X(_10473_));
 sky130_fd_sc_hd__nor2_1 _17475_ (.A(_09562_),
    .B(_09420_),
    .Y(_10474_));
 sky130_fd_sc_hd__a21oi_1 _17476_ (.A1(_09447_),
    .A2(_09794_),
    .B1(_10474_),
    .Y(_10475_));
 sky130_fd_sc_hd__and3_1 _17477_ (.A(_09447_),
    .B(_09794_),
    .C(_10474_),
    .X(_10476_));
 sky130_fd_sc_hd__nor2_1 _17478_ (.A(_10475_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__nor2_1 _17479_ (.A(_09328_),
    .B(_09666_),
    .Y(_10478_));
 sky130_fd_sc_hd__xnor2_1 _17480_ (.A(_10477_),
    .B(_10478_),
    .Y(_10479_));
 sky130_fd_sc_hd__o31a_1 _17481_ (.A1(_09091_),
    .A2(_09666_),
    .A3(_10345_),
    .B1(_10346_),
    .X(_10480_));
 sky130_fd_sc_hd__or2_1 _17482_ (.A(_10479_),
    .B(_10480_),
    .X(_10481_));
 sky130_fd_sc_hd__nand2_1 _17483_ (.A(_10479_),
    .B(_10480_),
    .Y(_10482_));
 sky130_fd_sc_hd__nand2_1 _17484_ (.A(_10481_),
    .B(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__nor2_1 _17485_ (.A(_09051_),
    .B(_09784_),
    .Y(_10484_));
 sky130_fd_sc_hd__xnor2_1 _17486_ (.A(_10483_),
    .B(_10484_),
    .Y(_10485_));
 sky130_fd_sc_hd__a21o_1 _17487_ (.A1(_10360_),
    .A2(_10361_),
    .B1(_10359_),
    .X(_10486_));
 sky130_fd_sc_hd__nor2_1 _17488_ (.A(_10383_),
    .B(_08795_),
    .Y(_10487_));
 sky130_fd_sc_hd__xnor2_1 _17489_ (.A(_10358_),
    .B(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__or3_1 _17490_ (.A(_10130_),
    .B(_09312_),
    .C(_10488_),
    .X(_10489_));
 sky130_fd_sc_hd__o21ai_1 _17491_ (.A1(_10130_),
    .A2(_09312_),
    .B1(_10488_),
    .Y(_10490_));
 sky130_fd_sc_hd__nand2_1 _17492_ (.A(_10489_),
    .B(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__o31ai_1 _17493_ (.A1(_10383_),
    .A2(_08708_),
    .A3(_10378_),
    .B1(_10381_),
    .Y(_10492_));
 sky130_fd_sc_hd__and2b_1 _17494_ (.A_N(_10491_),
    .B(_10492_),
    .X(_10493_));
 sky130_fd_sc_hd__and2b_1 _17495_ (.A_N(_10492_),
    .B(_10491_),
    .X(_10494_));
 sky130_fd_sc_hd__nor2_1 _17496_ (.A(_10493_),
    .B(_10494_),
    .Y(_10495_));
 sky130_fd_sc_hd__xnor2_1 _17497_ (.A(_10486_),
    .B(_10495_),
    .Y(_10496_));
 sky130_fd_sc_hd__a21oi_1 _17498_ (.A1(_10356_),
    .A2(_10365_),
    .B1(_10363_),
    .Y(_10497_));
 sky130_fd_sc_hd__nor2_1 _17499_ (.A(_10496_),
    .B(_10497_),
    .Y(_10498_));
 sky130_fd_sc_hd__and2_1 _17500_ (.A(_10496_),
    .B(_10497_),
    .X(_10499_));
 sky130_fd_sc_hd__nor2_1 _17501_ (.A(_10498_),
    .B(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__xnor2_1 _17502_ (.A(_10485_),
    .B(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__a21o_1 _17503_ (.A1(_10399_),
    .A2(_10473_),
    .B1(_10501_),
    .X(_10502_));
 sky130_fd_sc_hd__nand3_1 _17504_ (.A(_10399_),
    .B(_10473_),
    .C(_10501_),
    .Y(_10503_));
 sky130_fd_sc_hd__nand2_1 _17505_ (.A(_10502_),
    .B(_10503_),
    .Y(_10504_));
 sky130_fd_sc_hd__xnor2_2 _17506_ (.A(_10472_),
    .B(_10504_),
    .Y(_10505_));
 sky130_fd_sc_hd__a21o_1 _17507_ (.A1(_10385_),
    .A2(_10397_),
    .B1(_10395_),
    .X(_10506_));
 sky130_fd_sc_hd__nand2_1 _17508_ (.A(_10405_),
    .B(_10412_),
    .Y(_10507_));
 sky130_fd_sc_hd__or2b_1 _17509_ (.A(_10413_),
    .B_N(_10403_),
    .X(_10508_));
 sky130_fd_sc_hd__nor2_1 _17510_ (.A(_08329_),
    .B(_10380_),
    .Y(_10509_));
 sky130_fd_sc_hd__nor2_1 _17511_ (.A(_08317_),
    .B(_08634_),
    .Y(_10510_));
 sky130_fd_sc_hd__xnor2_1 _17512_ (.A(_10509_),
    .B(_10510_),
    .Y(_10511_));
 sky130_fd_sc_hd__or3_1 _17513_ (.A(_10379_),
    .B(_08705_),
    .C(_10511_),
    .X(_10512_));
 sky130_fd_sc_hd__o21ai_1 _17514_ (.A1(_10379_),
    .A2(_08705_),
    .B1(_10511_),
    .Y(_10513_));
 sky130_fd_sc_hd__and2_1 _17515_ (.A(_10512_),
    .B(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__or2_1 _17516_ (.A(_08873_),
    .B(_09595_),
    .X(_10515_));
 sky130_fd_sc_hd__nor2_1 _17517_ (.A(_08872_),
    .B(_09484_),
    .Y(_10516_));
 sky130_fd_sc_hd__xor2_2 _17518_ (.A(_10515_),
    .B(_10516_),
    .X(_10517_));
 sky130_fd_sc_hd__or2_1 _17519_ (.A(_08717_),
    .B(_09477_),
    .X(_10518_));
 sky130_fd_sc_hd__xnor2_2 _17520_ (.A(_10517_),
    .B(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__clkbuf_4 _17521_ (.A(_08873_),
    .X(_10520_));
 sky130_fd_sc_hd__o31a_1 _17522_ (.A1(_10520_),
    .A2(_09477_),
    .A3(_10387_),
    .B1(_10390_),
    .X(_10521_));
 sky130_fd_sc_hd__xor2_1 _17523_ (.A(_10519_),
    .B(_10521_),
    .X(_10522_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_10514_),
    .B(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__or2_1 _17525_ (.A(_10514_),
    .B(_10522_),
    .X(_10524_));
 sky130_fd_sc_hd__nand2_1 _17526_ (.A(_10523_),
    .B(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__a21o_1 _17527_ (.A1(_10507_),
    .A2(_10508_),
    .B1(_10525_),
    .X(_10526_));
 sky130_fd_sc_hd__nand3_1 _17528_ (.A(_10507_),
    .B(_10508_),
    .C(_10525_),
    .Y(_10527_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_10526_),
    .B(_10527_),
    .Y(_10528_));
 sky130_fd_sc_hd__xnor2_1 _17530_ (.A(_10506_),
    .B(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__a21bo_1 _17531_ (.A1(_10409_),
    .A2(_10411_),
    .B1_N(_10408_),
    .X(_10530_));
 sky130_fd_sc_hd__nand2_1 _17532_ (.A(_10419_),
    .B(_10420_),
    .Y(_10531_));
 sky130_fd_sc_hd__or4_1 _17533_ (.A(_09103_),
    .B(_10406_),
    .C(_10407_),
    .D(_10415_),
    .X(_10532_));
 sky130_fd_sc_hd__o22ai_2 _17534_ (.A1(_10406_),
    .A2(_10407_),
    .B1(_10416_),
    .B2(_09108_),
    .Y(_10533_));
 sky130_fd_sc_hd__nand2_1 _17535_ (.A(_10532_),
    .B(_10533_),
    .Y(_10534_));
 sky130_fd_sc_hd__nor2_1 _17536_ (.A(_09582_),
    .B(_09861_),
    .Y(_10535_));
 sky130_fd_sc_hd__xor2_1 _17537_ (.A(_10534_),
    .B(_10535_),
    .X(_10536_));
 sky130_fd_sc_hd__xor2_1 _17538_ (.A(_10531_),
    .B(_10536_),
    .X(_10537_));
 sky130_fd_sc_hd__xnor2_1 _17539_ (.A(_10530_),
    .B(_10537_),
    .Y(_10538_));
 sky130_fd_sc_hd__buf_2 _17540_ (.A(_10174_),
    .X(_10539_));
 sky130_fd_sc_hd__nor2_1 _17541_ (.A(_09593_),
    .B(_10539_),
    .Y(_10540_));
 sky130_fd_sc_hd__or3_2 _17542_ (.A(_09138_),
    .B(_09139_),
    .C(_10168_),
    .X(_10541_));
 sky130_fd_sc_hd__a21oi_1 _17543_ (.A1(_09138_),
    .A2(_09139_),
    .B1(_10168_),
    .Y(_10542_));
 sky130_fd_sc_hd__nand2_2 _17544_ (.A(_10541_),
    .B(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__xnor2_1 _17545_ (.A(_10540_),
    .B(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__xnor2_1 _17546_ (.A(_10302_),
    .B(_10544_),
    .Y(_10545_));
 sky130_fd_sc_hd__and2_1 _17547_ (.A(_10301_),
    .B(_10422_),
    .X(_10546_));
 sky130_fd_sc_hd__xor2_1 _17548_ (.A(_10545_),
    .B(_10546_),
    .X(_10547_));
 sky130_fd_sc_hd__xnor2_1 _17549_ (.A(_10538_),
    .B(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__a21boi_1 _17550_ (.A1(_10414_),
    .A2(_10426_),
    .B1_N(_10425_),
    .Y(_10549_));
 sky130_fd_sc_hd__nor2_1 _17551_ (.A(_10548_),
    .B(_10549_),
    .Y(_10550_));
 sky130_fd_sc_hd__and2_1 _17552_ (.A(_10548_),
    .B(_10549_),
    .X(_10551_));
 sky130_fd_sc_hd__nor2_1 _17553_ (.A(_10550_),
    .B(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__xnor2_1 _17554_ (.A(_10529_),
    .B(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__a21oi_1 _17555_ (.A1(_10402_),
    .A2(_10432_),
    .B1(_10430_),
    .Y(_10554_));
 sky130_fd_sc_hd__nor2_1 _17556_ (.A(_10553_),
    .B(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__and2_1 _17557_ (.A(_10553_),
    .B(_10554_),
    .X(_10556_));
 sky130_fd_sc_hd__nor2_1 _17558_ (.A(_10555_),
    .B(_10556_),
    .Y(_10557_));
 sky130_fd_sc_hd__xnor2_2 _17559_ (.A(_10505_),
    .B(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__nor2_1 _17560_ (.A(_10433_),
    .B(_10435_),
    .Y(_10559_));
 sky130_fd_sc_hd__a21oi_2 _17561_ (.A1(_10375_),
    .A2(_10436_),
    .B1(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__xor2_2 _17562_ (.A(_10558_),
    .B(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__xnor2_2 _17563_ (.A(_10471_),
    .B(_10561_),
    .Y(_10562_));
 sky130_fd_sc_hd__a21oi_2 _17564_ (.A1(_10342_),
    .A2(_10440_),
    .B1(_10439_),
    .Y(_10563_));
 sky130_fd_sc_hd__xor2_2 _17565_ (.A(_10562_),
    .B(_10563_),
    .X(_10564_));
 sky130_fd_sc_hd__xnor2_2 _17566_ (.A(_10340_),
    .B(_10564_),
    .Y(_10565_));
 sky130_fd_sc_hd__a21oi_1 _17567_ (.A1(_10465_),
    .A2(_10466_),
    .B1(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__and3_1 _17568_ (.A(_10465_),
    .B(_10466_),
    .C(_10565_),
    .X(_10567_));
 sky130_fd_sc_hd__or2_1 _17569_ (.A(_10566_),
    .B(_10567_),
    .X(_10568_));
 sky130_fd_sc_hd__a21o_1 _17570_ (.A1(_10462_),
    .A2(_10464_),
    .B1(_10568_),
    .X(_10569_));
 sky130_fd_sc_hd__nand2_1 _17571_ (.A(_06204_),
    .B(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__a31o_2 _17572_ (.A1(_10462_),
    .A2(_10464_),
    .A3(_10568_),
    .B1(_10570_),
    .X(_10571_));
 sky130_fd_sc_hd__o31ai_1 _17573_ (.A1(_10010_),
    .A2(_10460_),
    .A3(_10461_),
    .B1(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__mux2_1 _17574_ (.A0(_10572_),
    .A1(net4501),
    .S(net4903),
    .X(_10573_));
 sky130_fd_sc_hd__clkbuf_1 _17575_ (.A(_10573_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_1 _17576_ (.A(net4403),
    .B(net7373),
    .Y(_10574_));
 sky130_fd_sc_hd__or2_1 _17577_ (.A(net4403),
    .B(net7373),
    .X(_10575_));
 sky130_fd_sc_hd__nand2_1 _17578_ (.A(net7374),
    .B(_10575_),
    .Y(_10576_));
 sky130_fd_sc_hd__nor2_1 _17579_ (.A(_10458_),
    .B(_10460_),
    .Y(_10577_));
 sky130_fd_sc_hd__xnor2_1 _17580_ (.A(net7375),
    .B(_10577_),
    .Y(_10578_));
 sky130_fd_sc_hd__or2b_1 _17581_ (.A(_10504_),
    .B_N(_10472_),
    .X(_10579_));
 sky130_fd_sc_hd__o31a_1 _17582_ (.A1(_09051_),
    .A2(_09784_),
    .A3(_10483_),
    .B1(_10481_),
    .X(_10580_));
 sky130_fd_sc_hd__a21oi_2 _17583_ (.A1(_10502_),
    .A2(_10579_),
    .B1(_10580_),
    .Y(_10581_));
 sky130_fd_sc_hd__and3_1 _17584_ (.A(_10502_),
    .B(_10579_),
    .C(_10580_),
    .X(_10582_));
 sky130_fd_sc_hd__nor2_1 _17585_ (.A(_10581_),
    .B(_10582_),
    .Y(_10583_));
 sky130_fd_sc_hd__a21o_1 _17586_ (.A1(_10485_),
    .A2(_10500_),
    .B1(_10498_),
    .X(_10584_));
 sky130_fd_sc_hd__or2b_1 _17587_ (.A(_10528_),
    .B_N(_10506_),
    .X(_10585_));
 sky130_fd_sc_hd__nor2_1 _17588_ (.A(_10130_),
    .B(_09538_),
    .Y(_10586_));
 sky130_fd_sc_hd__o22a_1 _17589_ (.A1(_10130_),
    .A2(_09420_),
    .B1(_09538_),
    .B2(_09562_),
    .X(_10587_));
 sky130_fd_sc_hd__a21oi_1 _17590_ (.A1(_10474_),
    .A2(_10586_),
    .B1(_10587_),
    .Y(_10588_));
 sky130_fd_sc_hd__and2b_1 _17591_ (.A_N(_09805_),
    .B(_09447_),
    .X(_10589_));
 sky130_fd_sc_hd__xnor2_1 _17592_ (.A(_10588_),
    .B(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__a21oi_1 _17593_ (.A1(_10477_),
    .A2(_10478_),
    .B1(_10476_),
    .Y(_10591_));
 sky130_fd_sc_hd__nor2_1 _17594_ (.A(_10590_),
    .B(_10591_),
    .Y(_10592_));
 sky130_fd_sc_hd__and2_1 _17595_ (.A(_10590_),
    .B(_10591_),
    .X(_10593_));
 sky130_fd_sc_hd__nor2_1 _17596_ (.A(_10592_),
    .B(_10593_),
    .Y(_10594_));
 sky130_fd_sc_hd__and2_1 _17597_ (.A(_09328_),
    .B(net7378),
    .X(_10595_));
 sky130_fd_sc_hd__xor2_1 _17598_ (.A(_10594_),
    .B(_10595_),
    .X(_10596_));
 sky130_fd_sc_hd__a21bo_1 _17599_ (.A1(_10358_),
    .A2(_10487_),
    .B1_N(_10489_),
    .X(_10597_));
 sky130_fd_sc_hd__nor2_1 _17600_ (.A(_08546_),
    .B(_09251_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_1 _17601_ (.A(_08641_),
    .B(_08793_),
    .Y(_01653_));
 sky130_fd_sc_hd__xnor2_1 _17602_ (.A(_01652_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__or3_1 _17603_ (.A(_10257_),
    .B(_09312_),
    .C(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__o21ai_1 _17604_ (.A1(_10257_),
    .A2(_09312_),
    .B1(_01654_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _17605_ (.A(_01655_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__a21bo_1 _17606_ (.A1(_10509_),
    .A2(_10510_),
    .B1_N(_10512_),
    .X(_01658_));
 sky130_fd_sc_hd__and2b_1 _17607_ (.A_N(_01657_),
    .B(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__and2b_1 _17608_ (.A_N(_01658_),
    .B(_01657_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_1 _17609_ (.A(_01659_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__xnor2_1 _17610_ (.A(_10597_),
    .B(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__a21oi_1 _17611_ (.A1(_10486_),
    .A2(_10495_),
    .B1(_10493_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_1 _17612_ (.A(_01662_),
    .B(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__and2_1 _17613_ (.A(_01662_),
    .B(_01663_),
    .X(_01665_));
 sky130_fd_sc_hd__nor2_1 _17614_ (.A(_01664_),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__xnor2_1 _17615_ (.A(_10596_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__a21o_1 _17616_ (.A1(_10526_),
    .A2(_10585_),
    .B1(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__nand3_1 _17617_ (.A(_10526_),
    .B(_10585_),
    .C(_01667_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_1 _17618_ (.A(_01668_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__xnor2_1 _17619_ (.A(_10584_),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__o21ai_2 _17620_ (.A1(_10519_),
    .A2(_10521_),
    .B1(_10523_),
    .Y(_01672_));
 sky130_fd_sc_hd__or2b_1 _17621_ (.A(_10536_),
    .B_N(_10531_),
    .X(_01673_));
 sky130_fd_sc_hd__or2b_1 _17622_ (.A(_10537_),
    .B_N(_10530_),
    .X(_01674_));
 sky130_fd_sc_hd__nand2_2 _17623_ (.A(_08596_),
    .B(_08597_),
    .Y(_01675_));
 sky130_fd_sc_hd__or2_1 _17624_ (.A(_08329_),
    .B(_01675_),
    .X(_01676_));
 sky130_fd_sc_hd__nor2_1 _17625_ (.A(_10259_),
    .B(_08630_),
    .Y(_01677_));
 sky130_fd_sc_hd__xnor2_1 _17626_ (.A(_01676_),
    .B(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor2_1 _17627_ (.A(_08643_),
    .B(_08708_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _17628_ (.A(_01678_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__or2_1 _17629_ (.A(_01678_),
    .B(_01679_),
    .X(_01681_));
 sky130_fd_sc_hd__and2_1 _17630_ (.A(_01680_),
    .B(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__or4_1 _17631_ (.A(_08872_),
    .B(_08873_),
    .C(_09484_),
    .D(_09861_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_2 _17632_ (.A(_08872_),
    .X(_01684_));
 sky130_fd_sc_hd__o22ai_1 _17633_ (.A1(_10520_),
    .A2(_09484_),
    .B1(_09861_),
    .B2(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__and2_1 _17634_ (.A(_01683_),
    .B(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_1 _17635_ (.A(_08717_),
    .B(_09595_),
    .Y(_01687_));
 sky130_fd_sc_hd__xnor2_2 _17636_ (.A(_01686_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__or2_1 _17637_ (.A(_10517_),
    .B(_10518_),
    .X(_01689_));
 sky130_fd_sc_hd__o31a_1 _17638_ (.A1(_01684_),
    .A2(_09484_),
    .A3(_10515_),
    .B1(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__xor2_1 _17639_ (.A(_01688_),
    .B(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(_01682_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__or2_1 _17641_ (.A(_01682_),
    .B(_01691_),
    .X(_01693_));
 sky130_fd_sc_hd__nand2_1 _17642_ (.A(_01692_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21o_1 _17643_ (.A1(_01673_),
    .A2(_01674_),
    .B1(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nand3_1 _17644_ (.A(_01673_),
    .B(_01674_),
    .C(_01694_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _17645_ (.A(_01695_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__xnor2_1 _17646_ (.A(_01672_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__a21bo_1 _17647_ (.A1(_10533_),
    .A2(_10535_),
    .B1_N(_10532_),
    .X(_01699_));
 sky130_fd_sc_hd__or3_1 _17648_ (.A(_09593_),
    .B(_10539_),
    .C(_10543_),
    .X(_01700_));
 sky130_fd_sc_hd__or4_1 _17649_ (.A(_09108_),
    .B(_10406_),
    .C(_10416_),
    .D(_10174_),
    .X(_01701_));
 sky130_fd_sc_hd__o22ai_1 _17650_ (.A1(_10406_),
    .A2(_10416_),
    .B1(_10539_),
    .B2(_09108_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_1 _17651_ (.A(_01701_),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__nor2_1 _17652_ (.A(_09582_),
    .B(_10407_),
    .Y(_01704_));
 sky130_fd_sc_hd__xor2_1 _17653_ (.A(_01703_),
    .B(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__a21o_1 _17654_ (.A1(_10541_),
    .A2(_01700_),
    .B1(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__nand3_1 _17655_ (.A(_10541_),
    .B(_01700_),
    .C(_01705_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _17656_ (.A(_01706_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__xnor2_1 _17657_ (.A(_01699_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _17658_ (.A(_10302_),
    .B(_10544_),
    .Y(_01710_));
 sky130_fd_sc_hd__buf_2 _17659_ (.A(_10168_),
    .X(_01711_));
 sky130_fd_sc_hd__nor2_1 _17660_ (.A(_09593_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__mux2_1 _17661_ (.A0(_09593_),
    .A1(_01712_),
    .S(_10543_),
    .X(_01713_));
 sky130_fd_sc_hd__xnor2_1 _17662_ (.A(_10302_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__a21oi_1 _17663_ (.A1(_10301_),
    .A2(_01710_),
    .B1(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__and3_1 _17664_ (.A(_10301_),
    .B(_01710_),
    .C(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__nor2_1 _17665_ (.A(_01715_),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__xnor2_1 _17666_ (.A(_01709_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__nor2_1 _17667_ (.A(_10545_),
    .B(_10546_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21oi_1 _17668_ (.A1(_10538_),
    .A2(_10547_),
    .B1(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _17669_ (.A(_01718_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__and2_1 _17670_ (.A(_01718_),
    .B(_01720_),
    .X(_01722_));
 sky130_fd_sc_hd__nor2_1 _17671_ (.A(_01721_),
    .B(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__xnor2_1 _17672_ (.A(_01698_),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__a21oi_1 _17673_ (.A1(_10529_),
    .A2(_10552_),
    .B1(_10550_),
    .Y(_01725_));
 sky130_fd_sc_hd__xor2_1 _17674_ (.A(_01724_),
    .B(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__xnor2_1 _17675_ (.A(_01671_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__a21oi_1 _17676_ (.A1(_10505_),
    .A2(_10557_),
    .B1(_10555_),
    .Y(_01728_));
 sky130_fd_sc_hd__nor2_1 _17677_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__and2_1 _17678_ (.A(_01727_),
    .B(_01728_),
    .X(_01730_));
 sky130_fd_sc_hd__nor2_1 _17679_ (.A(_01729_),
    .B(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__xnor2_1 _17680_ (.A(_10583_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_1 _17681_ (.A(_10558_),
    .B(_10560_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_1 _17682_ (.A1(_10471_),
    .A2(_10561_),
    .B1(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__xor2_1 _17683_ (.A(_01732_),
    .B(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__xnor2_1 _17684_ (.A(_10469_),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__nor2_1 _17685_ (.A(_10562_),
    .B(_10563_),
    .Y(_01737_));
 sky130_fd_sc_hd__a21oi_1 _17686_ (.A1(_10340_),
    .A2(_10564_),
    .B1(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _17687_ (.A(_01736_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__and2_1 _17688_ (.A(_01736_),
    .B(_01738_),
    .X(_01740_));
 sky130_fd_sc_hd__or2_1 _17689_ (.A(_01739_),
    .B(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__a21o_1 _17690_ (.A1(_10465_),
    .A2(_10466_),
    .B1(_10565_),
    .X(_01742_));
 sky130_fd_sc_hd__a21o_1 _17691_ (.A1(_10462_),
    .A2(_01742_),
    .B1(_10567_),
    .X(_01743_));
 sky130_fd_sc_hd__o31a_1 _17692_ (.A1(_10463_),
    .A2(_10453_),
    .A3(_10568_),
    .B1(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__and2_1 _17693_ (.A(_01741_),
    .B(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__nor2_1 _17694_ (.A(_01741_),
    .B(_01744_),
    .Y(_01746_));
 sky130_fd_sc_hd__or3_2 _17695_ (.A(_09999_),
    .B(_01745_),
    .C(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__o21ai_1 _17696_ (.A1(_06206_),
    .A2(net7376),
    .B1(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__clkbuf_8 _17697_ (.A(net4902),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _17698_ (.A0(_01748_),
    .A1(net4403),
    .S(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__clkbuf_1 _17699_ (.A(_01750_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_1 _17700_ (.A(net4433),
    .B(net4593),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _17701_ (.A(net4433),
    .B(net4593),
    .Y(_01752_));
 sky130_fd_sc_hd__or2b_1 _17702_ (.A(_01751_),
    .B_N(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__o21a_1 _17703_ (.A1(net7375),
    .A2(_10577_),
    .B1(net7374),
    .X(_01754_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_01753_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__or2_1 _17705_ (.A(_01732_),
    .B(_01734_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_1 _17706_ (.A(_10469_),
    .B(_01735_),
    .Y(_01757_));
 sky130_fd_sc_hd__or2b_1 _17707_ (.A(_01670_),
    .B_N(_10584_),
    .X(_01758_));
 sky130_fd_sc_hd__a21oi_2 _17708_ (.A1(_10594_),
    .A2(_10595_),
    .B1(_10592_),
    .Y(_01759_));
 sky130_fd_sc_hd__a21oi_2 _17709_ (.A1(_01668_),
    .A2(_01758_),
    .B1(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__and3_1 _17710_ (.A(_01668_),
    .B(_01758_),
    .C(_01759_),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_1 _17711_ (.A(_01760_),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__a21o_1 _17712_ (.A1(_10596_),
    .A2(_01666_),
    .B1(_01664_),
    .X(_01763_));
 sky130_fd_sc_hd__or2b_1 _17713_ (.A(_01697_),
    .B_N(_01672_),
    .X(_01764_));
 sky130_fd_sc_hd__nor2_1 _17714_ (.A(_10257_),
    .B(_09420_),
    .Y(_01765_));
 sky130_fd_sc_hd__or2_1 _17715_ (.A(_10257_),
    .B(_09538_),
    .X(_01766_));
 sky130_fd_sc_hd__or3_1 _17716_ (.A(_10130_),
    .B(_09420_),
    .C(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__o21a_1 _17717_ (.A1(_10586_),
    .A2(_01765_),
    .B1(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__nor2_1 _17718_ (.A(_09562_),
    .B(_09805_),
    .Y(_01769_));
 sky130_fd_sc_hd__xnor2_1 _17719_ (.A(_01768_),
    .B(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__a22oi_1 _17720_ (.A1(_10474_),
    .A2(_10586_),
    .B1(_10588_),
    .B2(_10589_),
    .Y(_01771_));
 sky130_fd_sc_hd__or2_1 _17721_ (.A(_01770_),
    .B(_01771_),
    .X(_01772_));
 sky130_fd_sc_hd__nand2_1 _17722_ (.A(_01770_),
    .B(_01771_),
    .Y(_01773_));
 sky130_fd_sc_hd__nand2_1 _17723_ (.A(_01772_),
    .B(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2_1 _17724_ (.A(_09447_),
    .B(_09784_),
    .Y(_01775_));
 sky130_fd_sc_hd__xnor2_2 _17725_ (.A(_01774_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__a21bo_1 _17726_ (.A1(_01652_),
    .A2(_01653_),
    .B1_N(_01655_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_2 _17727_ (.A(_08630_),
    .X(_01778_));
 sky130_fd_sc_hd__or3_1 _17728_ (.A(_10259_),
    .B(_01778_),
    .C(_01676_),
    .X(_01779_));
 sky130_fd_sc_hd__or2_1 _17729_ (.A(_08643_),
    .B(_08795_),
    .X(_01780_));
 sky130_fd_sc_hd__or3_1 _17730_ (.A(_10379_),
    .B(_09249_),
    .C(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__o21ai_1 _17731_ (.A1(_10379_),
    .A2(_09249_),
    .B1(_01780_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_1 _17732_ (.A(_01781_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_1 _17733_ (.A(_10383_),
    .B(_09312_),
    .Y(_01784_));
 sky130_fd_sc_hd__xor2_1 _17734_ (.A(_01783_),
    .B(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__a21oi_1 _17735_ (.A1(_01779_),
    .A2(_01680_),
    .B1(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__and3_1 _17736_ (.A(_01779_),
    .B(_01680_),
    .C(_01785_),
    .X(_01787_));
 sky130_fd_sc_hd__nor2_1 _17737_ (.A(_01786_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__xnor2_1 _17738_ (.A(_01777_),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21oi_1 _17739_ (.A1(_10597_),
    .A2(_01661_),
    .B1(_01659_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _17740_ (.A(_01789_),
    .B(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__and2_1 _17741_ (.A(_01789_),
    .B(_01790_),
    .X(_01792_));
 sky130_fd_sc_hd__nor2_1 _17742_ (.A(_01791_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__xnor2_2 _17743_ (.A(_01776_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21o_1 _17744_ (.A1(_01695_),
    .A2(_01764_),
    .B1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__nand3_1 _17745_ (.A(_01695_),
    .B(_01764_),
    .C(_01794_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand2_1 _17746_ (.A(_01795_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__xnor2_1 _17747_ (.A(_01763_),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__o21ai_2 _17748_ (.A1(_01688_),
    .A2(_01690_),
    .B1(_01692_),
    .Y(_01799_));
 sky130_fd_sc_hd__or2b_1 _17749_ (.A(_01708_),
    .B_N(_01699_),
    .X(_01800_));
 sky130_fd_sc_hd__or2_1 _17750_ (.A(_10259_),
    .B(_09231_),
    .X(_01801_));
 sky130_fd_sc_hd__buf_2 _17751_ (.A(_08329_),
    .X(_01802_));
 sky130_fd_sc_hd__nor2_1 _17752_ (.A(_01802_),
    .B(_01778_),
    .Y(_01803_));
 sky130_fd_sc_hd__xnor2_1 _17753_ (.A(_01801_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _17754_ (.A(_08634_),
    .B(_08708_),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2_1 _17755_ (.A(_01804_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__or2_1 _17756_ (.A(_01804_),
    .B(_01805_),
    .X(_01807_));
 sky130_fd_sc_hd__and2_1 _17757_ (.A(_01806_),
    .B(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__nor2_1 _17758_ (.A(_10520_),
    .B(_09861_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _17759_ (.A(_01684_),
    .B(_10407_),
    .Y(_01810_));
 sky130_fd_sc_hd__xnor2_1 _17760_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__buf_2 _17761_ (.A(_08717_),
    .X(_01812_));
 sky130_fd_sc_hd__nor2_1 _17762_ (.A(_01812_),
    .B(_09484_),
    .Y(_01813_));
 sky130_fd_sc_hd__xor2_1 _17763_ (.A(_01811_),
    .B(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__a21boi_1 _17764_ (.A1(_01685_),
    .A2(_01687_),
    .B1_N(_01683_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _17765_ (.A(_01814_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__and2_1 _17766_ (.A(_01814_),
    .B(_01815_),
    .X(_01817_));
 sky130_fd_sc_hd__nor2_1 _17767_ (.A(_01816_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__xnor2_1 _17768_ (.A(_01808_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__a21o_1 _17769_ (.A1(_01706_),
    .A2(_01800_),
    .B1(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__nand3_1 _17770_ (.A(_01706_),
    .B(_01800_),
    .C(_01819_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _17771_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__xnor2_1 _17772_ (.A(_01799_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__a21bo_1 _17773_ (.A1(_01702_),
    .A2(_01704_),
    .B1_N(_01701_),
    .X(_01824_));
 sky130_fd_sc_hd__o21ai_4 _17774_ (.A1(_09593_),
    .A2(_10543_),
    .B1(_10541_),
    .Y(_01825_));
 sky130_fd_sc_hd__o22ai_1 _17775_ (.A1(_09108_),
    .A2(_01711_),
    .B1(_10539_),
    .B2(_10406_),
    .Y(_01826_));
 sky130_fd_sc_hd__or4_1 _17776_ (.A(_09108_),
    .B(_10406_),
    .C(_01711_),
    .D(_10539_),
    .X(_01827_));
 sky130_fd_sc_hd__nand2_1 _17777_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__nor2_1 _17778_ (.A(_09582_),
    .B(_10416_),
    .Y(_01829_));
 sky130_fd_sc_hd__xnor2_1 _17779_ (.A(_01828_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__xnor2_1 _17780_ (.A(_01825_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__xnor2_1 _17781_ (.A(_01824_),
    .B(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2b_2 _17782_ (.A_N(_10301_),
    .B(_01713_),
    .Y(_01833_));
 sky130_fd_sc_hd__or3_1 _17783_ (.A(_10298_),
    .B(_10299_),
    .C(_01713_),
    .X(_01834_));
 sky130_fd_sc_hd__and2_1 _17784_ (.A(_01833_),
    .B(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__buf_2 _17785_ (.A(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__nand2_1 _17786_ (.A(_01832_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__or2_1 _17787_ (.A(_01832_),
    .B(_01836_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(_01837_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21oi_1 _17789_ (.A1(_01709_),
    .A2(_01717_),
    .B1(_01715_),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_1 _17790_ (.A(_01839_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__and2_1 _17791_ (.A(_01839_),
    .B(_01840_),
    .X(_01842_));
 sky130_fd_sc_hd__nor2_1 _17792_ (.A(_01841_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__xnor2_1 _17793_ (.A(_01823_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__a21oi_1 _17794_ (.A1(_01698_),
    .A2(_01723_),
    .B1(_01721_),
    .Y(_01845_));
 sky130_fd_sc_hd__nor2_1 _17795_ (.A(_01844_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__and2_1 _17796_ (.A(_01844_),
    .B(_01845_),
    .X(_01847_));
 sky130_fd_sc_hd__nor2_1 _17797_ (.A(_01846_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__xnor2_1 _17798_ (.A(_01798_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _17799_ (.A(_01724_),
    .B(_01725_),
    .Y(_01850_));
 sky130_fd_sc_hd__a21o_1 _17800_ (.A1(_01671_),
    .A2(_01726_),
    .B1(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__xnor2_1 _17801_ (.A(_01849_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__xnor2_1 _17802_ (.A(_01762_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__a21oi_1 _17803_ (.A1(_10583_),
    .A2(_01731_),
    .B1(_01729_),
    .Y(_01854_));
 sky130_fd_sc_hd__xor2_1 _17804_ (.A(_01853_),
    .B(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__xnor2_1 _17805_ (.A(_10581_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand3_1 _17806_ (.A(_01756_),
    .B(_01757_),
    .C(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21o_1 _17807_ (.A1(_01756_),
    .A2(_01757_),
    .B1(_01856_),
    .X(_01858_));
 sky130_fd_sc_hd__nand2_1 _17808_ (.A(_01857_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _17809_ (.A(_01739_),
    .B(_01746_),
    .Y(_01860_));
 sky130_fd_sc_hd__o21ai_1 _17810_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_06205_),
    .Y(_01861_));
 sky130_fd_sc_hd__a21o_2 _17811_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__o21ai_1 _17812_ (.A1(_06206_),
    .A2(_01755_),
    .B1(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__mux2_1 _17813_ (.A0(_01863_),
    .A1(net4433),
    .S(_01749_),
    .X(_01864_));
 sky130_fd_sc_hd__clkbuf_1 _17814_ (.A(_01864_),
    .X(_00544_));
 sky130_fd_sc_hd__nor2_1 _17815_ (.A(net4558),
    .B(net4639),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _17816_ (.A(net4558),
    .B(net4639),
    .Y(_01866_));
 sky130_fd_sc_hd__or2b_1 _17817_ (.A(_01865_),
    .B_N(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__o21a_1 _17818_ (.A1(_01751_),
    .A2(_01754_),
    .B1(_01752_),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_1 _17819_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__buf_4 _17820_ (.A(_06204_),
    .X(_01870_));
 sky130_fd_sc_hd__a21o_1 _17821_ (.A1(_01867_),
    .A2(_01868_),
    .B1(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__or2b_1 _17822_ (.A(_01797_),
    .B_N(_01763_),
    .X(_01872_));
 sky130_fd_sc_hd__o31a_1 _17823_ (.A1(_09447_),
    .A2(_09784_),
    .A3(_01774_),
    .B1(_01772_),
    .X(_01873_));
 sky130_fd_sc_hd__a21oi_2 _17824_ (.A1(_01795_),
    .A2(_01872_),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__and3_1 _17825_ (.A(_01795_),
    .B(_01872_),
    .C(_01873_),
    .X(_01875_));
 sky130_fd_sc_hd__nor2_1 _17826_ (.A(_01874_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a21o_1 _17827_ (.A1(_01776_),
    .A2(_01793_),
    .B1(_01791_),
    .X(_01877_));
 sky130_fd_sc_hd__or2b_1 _17828_ (.A(_01822_),
    .B_N(_01799_),
    .X(_01878_));
 sky130_fd_sc_hd__o21ai_1 _17829_ (.A1(_10383_),
    .A2(_09420_),
    .B1(_01766_),
    .Y(_01879_));
 sky130_fd_sc_hd__or3_1 _17830_ (.A(_10383_),
    .B(_09420_),
    .C(_01766_),
    .X(_01880_));
 sky130_fd_sc_hd__nand2_1 _17831_ (.A(_01879_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_1 _17832_ (.A(_10130_),
    .B(_09805_),
    .Y(_01882_));
 sky130_fd_sc_hd__xor2_1 _17833_ (.A(_01881_),
    .B(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__a21boi_1 _17834_ (.A1(_01768_),
    .A2(_01769_),
    .B1_N(_01767_),
    .Y(_01884_));
 sky130_fd_sc_hd__nor2_1 _17835_ (.A(_01883_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__and2_1 _17836_ (.A(_01883_),
    .B(_01884_),
    .X(_01886_));
 sky130_fd_sc_hd__nor2_1 _17837_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__and2_1 _17838_ (.A(_09562_),
    .B(net7378),
    .X(_01888_));
 sky130_fd_sc_hd__xor2_2 _17839_ (.A(_01887_),
    .B(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__o31ai_2 _17840_ (.A1(_10383_),
    .A2(_09312_),
    .A3(_01783_),
    .B1(_01781_),
    .Y(_01890_));
 sky130_fd_sc_hd__or3_1 _17841_ (.A(_01802_),
    .B(_01778_),
    .C(_01801_),
    .X(_01891_));
 sky130_fd_sc_hd__or2_1 _17842_ (.A(_01675_),
    .B(_08793_),
    .X(_01892_));
 sky130_fd_sc_hd__nor2_1 _17843_ (.A(_10380_),
    .B(_09249_),
    .Y(_01893_));
 sky130_fd_sc_hd__xnor2_1 _17844_ (.A(_01892_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__nor2_1 _17845_ (.A(_10379_),
    .B(_09310_),
    .Y(_01895_));
 sky130_fd_sc_hd__xnor2_1 _17846_ (.A(_01894_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__a21oi_1 _17847_ (.A1(_01891_),
    .A2(_01806_),
    .B1(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__and3_1 _17848_ (.A(_01891_),
    .B(_01806_),
    .C(_01896_),
    .X(_01898_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(_01897_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__xnor2_1 _17850_ (.A(_01890_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__a21oi_1 _17851_ (.A1(_01777_),
    .A2(_01788_),
    .B1(_01786_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _17852_ (.A(_01900_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__and2_1 _17853_ (.A(_01900_),
    .B(_01901_),
    .X(_01903_));
 sky130_fd_sc_hd__nor2_1 _17854_ (.A(_01902_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__xnor2_1 _17855_ (.A(_01889_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a21o_1 _17856_ (.A1(_01820_),
    .A2(_01878_),
    .B1(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__nand3_1 _17857_ (.A(_01820_),
    .B(_01878_),
    .C(_01905_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _17858_ (.A(_01906_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__xnor2_2 _17859_ (.A(_01877_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__a21o_1 _17860_ (.A1(_01808_),
    .A2(_01818_),
    .B1(_01816_),
    .X(_01910_));
 sky130_fd_sc_hd__nand2_1 _17861_ (.A(_01825_),
    .B(_01830_),
    .Y(_01911_));
 sky130_fd_sc_hd__or2b_1 _17862_ (.A(_01831_),
    .B_N(_01824_),
    .X(_01912_));
 sky130_fd_sc_hd__or2_1 _17863_ (.A(_10259_),
    .B(_09375_),
    .X(_01913_));
 sky130_fd_sc_hd__or3_1 _17864_ (.A(_01802_),
    .B(_09231_),
    .C(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__o21ai_1 _17865_ (.A1(_01802_),
    .A2(_09231_),
    .B1(_01913_),
    .Y(_01915_));
 sky130_fd_sc_hd__and2_1 _17866_ (.A(_01914_),
    .B(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__nor2_1 _17867_ (.A(_01778_),
    .B(_08705_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _17868_ (.A(_01916_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__or2_1 _17869_ (.A(_01916_),
    .B(_01917_),
    .X(_01919_));
 sky130_fd_sc_hd__and2_1 _17870_ (.A(_01918_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__or4_1 _17871_ (.A(_01684_),
    .B(_10520_),
    .C(_10407_),
    .D(_10416_),
    .X(_01921_));
 sky130_fd_sc_hd__o22ai_1 _17872_ (.A1(_10520_),
    .A2(_10407_),
    .B1(_10416_),
    .B2(_01684_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _17873_ (.A(_01921_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__or2_1 _17874_ (.A(_01812_),
    .B(_09861_),
    .X(_01924_));
 sky130_fd_sc_hd__xnor2_1 _17875_ (.A(_01923_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_01809_),
    .B(_01810_),
    .Y(_01926_));
 sky130_fd_sc_hd__o31a_1 _17877_ (.A1(_01812_),
    .A2(_09484_),
    .A3(_01811_),
    .B1(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__nor2_1 _17878_ (.A(_01925_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__and2_1 _17879_ (.A(_01925_),
    .B(_01927_),
    .X(_01929_));
 sky130_fd_sc_hd__nor2_1 _17880_ (.A(_01928_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__xnor2_1 _17881_ (.A(_01920_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__a21o_1 _17882_ (.A1(_01911_),
    .A2(_01912_),
    .B1(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__nand3_1 _17883_ (.A(_01911_),
    .B(_01912_),
    .C(_01931_),
    .Y(_01933_));
 sky130_fd_sc_hd__nand2_1 _17884_ (.A(_01932_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__xnor2_1 _17885_ (.A(_01910_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__a21bo_1 _17886_ (.A1(_01826_),
    .A2(_01829_),
    .B1_N(_01827_),
    .X(_01936_));
 sky130_fd_sc_hd__or2_1 _17887_ (.A(_09582_),
    .B(_10539_),
    .X(_01937_));
 sky130_fd_sc_hd__or3_1 _17888_ (.A(_09108_),
    .B(_10406_),
    .C(_01711_),
    .X(_01938_));
 sky130_fd_sc_hd__a21oi_1 _17889_ (.A1(_09108_),
    .A2(_10406_),
    .B1(_01711_),
    .Y(_01939_));
 sky130_fd_sc_hd__nand2_2 _17890_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__xor2_1 _17891_ (.A(_01937_),
    .B(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__xnor2_1 _17892_ (.A(_01825_),
    .B(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__xnor2_1 _17893_ (.A(_01936_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__xnor2_1 _17894_ (.A(_01836_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__a21oi_1 _17895_ (.A1(_01833_),
    .A2(_01837_),
    .B1(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__and3_1 _17896_ (.A(_01833_),
    .B(_01837_),
    .C(_01944_),
    .X(_01946_));
 sky130_fd_sc_hd__nor2_1 _17897_ (.A(_01945_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__xnor2_1 _17898_ (.A(_01935_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__a21oi_1 _17899_ (.A1(_01823_),
    .A2(_01843_),
    .B1(_01841_),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_1 _17900_ (.A(_01948_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__and2_1 _17901_ (.A(_01948_),
    .B(_01949_),
    .X(_01951_));
 sky130_fd_sc_hd__nor2_1 _17902_ (.A(_01950_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__xnor2_1 _17903_ (.A(_01909_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__a21oi_1 _17904_ (.A1(_01798_),
    .A2(_01848_),
    .B1(_01846_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor2_1 _17905_ (.A(_01953_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _17906_ (.A(_01953_),
    .B(_01954_),
    .Y(_01956_));
 sky130_fd_sc_hd__and2b_1 _17907_ (.A_N(_01955_),
    .B(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__xnor2_1 _17908_ (.A(_01876_),
    .B(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__and2b_1 _17909_ (.A_N(_01849_),
    .B(_01851_),
    .X(_01959_));
 sky130_fd_sc_hd__a21oi_1 _17910_ (.A1(_01762_),
    .A2(_01852_),
    .B1(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__xor2_1 _17911_ (.A(_01958_),
    .B(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__xnor2_1 _17912_ (.A(_01760_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _17913_ (.A(_01853_),
    .B(_01854_),
    .Y(_01963_));
 sky130_fd_sc_hd__a21oi_1 _17914_ (.A1(_10581_),
    .A2(_01855_),
    .B1(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__or2_1 _17915_ (.A(_01962_),
    .B(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _17916_ (.A(_01962_),
    .B(_01964_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_2 _17917_ (.A(_01965_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__a311o_1 _17918_ (.A1(_01756_),
    .A2(_01757_),
    .A3(_01856_),
    .B1(_01738_),
    .C1(_01736_),
    .X(_01968_));
 sky130_fd_sc_hd__o311a_4 _17919_ (.A1(_01741_),
    .A2(_01744_),
    .A3(_01859_),
    .B1(_01968_),
    .C1(_01858_),
    .X(_01969_));
 sky130_fd_sc_hd__o21ai_1 _17920_ (.A1(_01967_),
    .A2(_01969_),
    .B1(_06205_),
    .Y(_01970_));
 sky130_fd_sc_hd__a21o_1 _17921_ (.A1(_01967_),
    .A2(_01969_),
    .B1(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__o21ai_1 _17922_ (.A1(_01869_),
    .A2(_01871_),
    .B1(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__mux2_1 _17923_ (.A0(_01972_),
    .A1(net4558),
    .S(_01749_),
    .X(_01973_));
 sky130_fd_sc_hd__clkbuf_1 _17924_ (.A(_01973_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _17925_ (.A(net4599),
    .B(net4530),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _17926_ (.A(net4599),
    .B(net4530),
    .Y(_01975_));
 sky130_fd_sc_hd__or2b_1 _17927_ (.A(_01974_),
    .B_N(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__o21a_1 _17928_ (.A1(_01865_),
    .A2(_01868_),
    .B1(_01866_),
    .X(_01977_));
 sky130_fd_sc_hd__nor2_1 _17929_ (.A(_01976_),
    .B(net7798),
    .Y(_01978_));
 sky130_fd_sc_hd__a21o_1 _17930_ (.A1(_01976_),
    .A2(_01977_),
    .B1(_01870_),
    .X(_01979_));
 sky130_fd_sc_hd__or2_1 _17931_ (.A(_01958_),
    .B(_01960_),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_1 _17932_ (.A(_01760_),
    .B(_01961_),
    .Y(_01981_));
 sky130_fd_sc_hd__or2b_1 _17933_ (.A(_01908_),
    .B_N(_01877_),
    .X(_01982_));
 sky130_fd_sc_hd__a21oi_2 _17934_ (.A1(_01887_),
    .A2(_01888_),
    .B1(_01885_),
    .Y(_01983_));
 sky130_fd_sc_hd__a21oi_4 _17935_ (.A1(_01906_),
    .A2(_01982_),
    .B1(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__and3_1 _17936_ (.A(_01906_),
    .B(_01982_),
    .C(_01983_),
    .X(_01985_));
 sky130_fd_sc_hd__nor2_1 _17937_ (.A(_01984_),
    .B(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__a21o_1 _17938_ (.A1(_01889_),
    .A2(_01904_),
    .B1(_01902_),
    .X(_01987_));
 sky130_fd_sc_hd__or2b_1 _17939_ (.A(_01934_),
    .B_N(_01910_),
    .X(_01988_));
 sky130_fd_sc_hd__nor2_1 _17940_ (.A(_08546_),
    .B(_09538_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor2_1 _17941_ (.A(_10379_),
    .B(_09418_),
    .Y(_01990_));
 sky130_fd_sc_hd__xnor2_1 _17942_ (.A(_01989_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__or2_1 _17943_ (.A(_10257_),
    .B(_09805_),
    .X(_01992_));
 sky130_fd_sc_hd__xnor2_1 _17944_ (.A(_01991_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__o31a_1 _17945_ (.A1(_10130_),
    .A2(_09805_),
    .A3(_01881_),
    .B1(_01880_),
    .X(_01994_));
 sky130_fd_sc_hd__or2_1 _17946_ (.A(_01993_),
    .B(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__nand2_1 _17947_ (.A(_01993_),
    .B(_01994_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand2_1 _17948_ (.A(_01995_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _17949_ (.A(_08849_),
    .B(_09784_),
    .Y(_01998_));
 sky130_fd_sc_hd__xnor2_1 _17950_ (.A(_01997_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__or2_1 _17951_ (.A(_08634_),
    .B(_09251_),
    .X(_02000_));
 sky130_fd_sc_hd__o2bb2ai_1 _17952_ (.A1_N(_01894_),
    .A2_N(_01895_),
    .B1(_02000_),
    .B2(_01780_),
    .Y(_02001_));
 sky130_fd_sc_hd__or3_1 _17953_ (.A(_01778_),
    .B(_08793_),
    .C(_02000_),
    .X(_02002_));
 sky130_fd_sc_hd__o21ai_1 _17954_ (.A1(_01778_),
    .A2(_08793_),
    .B1(_02000_),
    .Y(_02003_));
 sky130_fd_sc_hd__and2_1 _17955_ (.A(_02002_),
    .B(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__nor2_1 _17956_ (.A(_10380_),
    .B(_09310_),
    .Y(_02005_));
 sky130_fd_sc_hd__xnor2_1 _17957_ (.A(_02004_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__a21oi_1 _17958_ (.A1(_01914_),
    .A2(_01918_),
    .B1(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__and3_1 _17959_ (.A(_01914_),
    .B(_01918_),
    .C(_02006_),
    .X(_02008_));
 sky130_fd_sc_hd__nor2_1 _17960_ (.A(_02007_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__xnor2_1 _17961_ (.A(_02001_),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__a21oi_1 _17962_ (.A1(_01890_),
    .A2(_01899_),
    .B1(_01897_),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _17963_ (.A(_02010_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__and2_1 _17964_ (.A(_02010_),
    .B(_02011_),
    .X(_02013_));
 sky130_fd_sc_hd__nor2_1 _17965_ (.A(_02012_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__xnor2_1 _17966_ (.A(_01999_),
    .B(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__a21o_1 _17967_ (.A1(_01932_),
    .A2(_01988_),
    .B1(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__nand3_1 _17968_ (.A(_01932_),
    .B(_01988_),
    .C(_02015_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand2_1 _17969_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__xnor2_2 _17970_ (.A(_01987_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__o21ai_1 _17971_ (.A1(_01937_),
    .A2(_01940_),
    .B1(_01938_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _17972_ (.A(_09582_),
    .B(_01711_),
    .Y(_02021_));
 sky130_fd_sc_hd__mux2_2 _17973_ (.A0(_09582_),
    .A1(_02021_),
    .S(_01940_),
    .X(_02022_));
 sky130_fd_sc_hd__xnor2_4 _17974_ (.A(_01825_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__xnor2_1 _17975_ (.A(_02020_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _17976_ (.A(_01836_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__or2_1 _17977_ (.A(_01836_),
    .B(_02024_),
    .X(_02026_));
 sky130_fd_sc_hd__nand2_1 _17978_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__a21boi_1 _17979_ (.A1(_01836_),
    .A2(_01943_),
    .B1_N(_01833_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _17980_ (.A(_02027_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__and2_1 _17981_ (.A(_02027_),
    .B(_02028_),
    .X(_02030_));
 sky130_fd_sc_hd__nor2_1 _17982_ (.A(_02029_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__a21o_1 _17983_ (.A1(_01920_),
    .A2(_01930_),
    .B1(_01928_),
    .X(_02032_));
 sky130_fd_sc_hd__nand2_1 _17984_ (.A(_01825_),
    .B(_01941_),
    .Y(_02033_));
 sky130_fd_sc_hd__or2b_1 _17985_ (.A(_01942_),
    .B_N(_01936_),
    .X(_02034_));
 sky130_fd_sc_hd__nor2_1 _17986_ (.A(_10259_),
    .B(_09602_),
    .Y(_02035_));
 sky130_fd_sc_hd__nor2_1 _17987_ (.A(_01802_),
    .B(_09375_),
    .Y(_02036_));
 sky130_fd_sc_hd__xnor2_1 _17988_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__or3_1 _17989_ (.A(_09231_),
    .B(_08705_),
    .C(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__o21ai_1 _17990_ (.A1(_09231_),
    .A2(_08705_),
    .B1(_02037_),
    .Y(_02039_));
 sky130_fd_sc_hd__and2_1 _17991_ (.A(_02038_),
    .B(_02039_),
    .X(_02040_));
 sky130_fd_sc_hd__nor2_1 _17992_ (.A(_10520_),
    .B(_10416_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_1 _17993_ (.A(_01684_),
    .B(_10539_),
    .Y(_02042_));
 sky130_fd_sc_hd__xnor2_1 _17994_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_1 _17995_ (.A(_01812_),
    .B(_10407_),
    .Y(_02044_));
 sky130_fd_sc_hd__xor2_1 _17996_ (.A(_02043_),
    .B(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__o31a_1 _17997_ (.A1(_01812_),
    .A2(_09861_),
    .A3(_01923_),
    .B1(_01921_),
    .X(_02046_));
 sky130_fd_sc_hd__xor2_1 _17998_ (.A(_02045_),
    .B(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__xnor2_1 _17999_ (.A(_02040_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__a21o_1 _18000_ (.A1(_02033_),
    .A2(_02034_),
    .B1(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__nand3_1 _18001_ (.A(_02033_),
    .B(_02034_),
    .C(_02048_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _18002_ (.A(_02049_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__xnor2_1 _18003_ (.A(_02032_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_02031_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__a21oi_1 _18005_ (.A1(_01935_),
    .A2(_01947_),
    .B1(_01945_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _18006_ (.A(_02053_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__and2_1 _18007_ (.A(_02053_),
    .B(_02054_),
    .X(_02056_));
 sky130_fd_sc_hd__nor2_1 _18008_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__xnor2_2 _18009_ (.A(_02019_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21oi_2 _18010_ (.A1(_01909_),
    .A2(_01952_),
    .B1(_01950_),
    .Y(_02059_));
 sky130_fd_sc_hd__xor2_2 _18011_ (.A(_02058_),
    .B(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__xnor2_2 _18012_ (.A(_01986_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__a21oi_2 _18013_ (.A1(_01876_),
    .A2(_01956_),
    .B1(_01955_),
    .Y(_02062_));
 sky130_fd_sc_hd__xor2_2 _18014_ (.A(_02061_),
    .B(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__xnor2_1 _18015_ (.A(_01874_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__a21oi_1 _18016_ (.A1(_01980_),
    .A2(_01981_),
    .B1(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__and3_1 _18017_ (.A(_01980_),
    .B(_01981_),
    .C(_02064_),
    .X(_02066_));
 sky130_fd_sc_hd__or2_2 _18018_ (.A(_02065_),
    .B(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__o21a_1 _18019_ (.A1(_01967_),
    .A2(_01969_),
    .B1(_01965_),
    .X(_02068_));
 sky130_fd_sc_hd__o21ai_1 _18020_ (.A1(_02067_),
    .A2(_02068_),
    .B1(_06205_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21o_1 _18021_ (.A1(_02067_),
    .A2(_02068_),
    .B1(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__o21ai_1 _18022_ (.A1(net7799),
    .A2(_01979_),
    .B1(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__mux2_1 _18023_ (.A0(_02071_),
    .A1(net4599),
    .S(_01749_),
    .X(_02072_));
 sky130_fd_sc_hd__clkbuf_1 _18024_ (.A(_02072_),
    .X(_00546_));
 sky130_fd_sc_hd__or2_1 _18025_ (.A(net4497),
    .B(net4619),
    .X(_02073_));
 sky130_fd_sc_hd__nand2_1 _18026_ (.A(net4497),
    .B(net4619),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _18027_ (.A(_02073_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__o21ai_1 _18028_ (.A1(_01974_),
    .A2(_01977_),
    .B1(_01975_),
    .Y(_02076_));
 sky130_fd_sc_hd__xnor2_1 _18029_ (.A(_02075_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__or2b_1 _18030_ (.A(_02018_),
    .B_N(_01987_),
    .X(_02078_));
 sky130_fd_sc_hd__o31a_1 _18031_ (.A1(_08849_),
    .A2(_09784_),
    .A3(_01997_),
    .B1(_01995_),
    .X(_02079_));
 sky130_fd_sc_hd__a21oi_2 _18032_ (.A1(_02016_),
    .A2(_02078_),
    .B1(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__and3_1 _18033_ (.A(_02016_),
    .B(_02078_),
    .C(_02079_),
    .X(_02081_));
 sky130_fd_sc_hd__nor2_1 _18034_ (.A(_02080_),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__o21a_1 _18035_ (.A1(_09582_),
    .A2(_01940_),
    .B1(_01938_),
    .X(_02083_));
 sky130_fd_sc_hd__xor2_2 _18036_ (.A(_02023_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__xnor2_1 _18037_ (.A(_01836_),
    .B(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__a21o_1 _18038_ (.A1(_01833_),
    .A2(_02025_),
    .B1(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__nand3_1 _18039_ (.A(_01833_),
    .B(_02025_),
    .C(_02085_),
    .Y(_02087_));
 sky130_fd_sc_hd__and2_1 _18040_ (.A(_02086_),
    .B(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__nor2_1 _18041_ (.A(_02045_),
    .B(_02046_),
    .Y(_02089_));
 sky130_fd_sc_hd__a21o_1 _18042_ (.A1(_02040_),
    .A2(_02047_),
    .B1(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__nand2_1 _18043_ (.A(_01825_),
    .B(_02022_),
    .Y(_02091_));
 sky130_fd_sc_hd__or2b_1 _18044_ (.A(_02023_),
    .B_N(_02020_),
    .X(_02092_));
 sky130_fd_sc_hd__nand2_1 _18045_ (.A(_02091_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__or2_1 _18046_ (.A(_10259_),
    .B(_09732_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_1 _18047_ (.A(_01802_),
    .B(_09602_),
    .Y(_02095_));
 sky130_fd_sc_hd__xnor2_1 _18048_ (.A(_02094_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _18049_ (.A(_08705_),
    .B(_09375_),
    .Y(_02097_));
 sky130_fd_sc_hd__xnor2_1 _18050_ (.A(_02096_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__or4_1 _18051_ (.A(_01684_),
    .B(_10520_),
    .C(_10168_),
    .D(_10539_),
    .X(_02099_));
 sky130_fd_sc_hd__o22ai_1 _18052_ (.A1(_01684_),
    .A2(_01711_),
    .B1(_10539_),
    .B2(_10520_),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _18053_ (.A(_02099_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_1 _18054_ (.A(_01812_),
    .B(_10416_),
    .Y(_02102_));
 sky130_fd_sc_hd__xor2_1 _18055_ (.A(_02101_),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__nand2_1 _18056_ (.A(_02041_),
    .B(_02042_),
    .Y(_02104_));
 sky130_fd_sc_hd__o31a_1 _18057_ (.A1(_01812_),
    .A2(_10407_),
    .A3(_02043_),
    .B1(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__xor2_1 _18058_ (.A(_02103_),
    .B(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__xnor2_1 _18059_ (.A(_02098_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__xnor2_1 _18060_ (.A(_02093_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__xnor2_1 _18061_ (.A(_02090_),
    .B(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _18062_ (.A(_02088_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__or2_1 _18063_ (.A(_02088_),
    .B(_02109_),
    .X(_02111_));
 sky130_fd_sc_hd__nand2_1 _18064_ (.A(_02110_),
    .B(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__a21oi_1 _18065_ (.A1(_02031_),
    .A2(_02052_),
    .B1(_02029_),
    .Y(_02113_));
 sky130_fd_sc_hd__xor2_1 _18066_ (.A(_02112_),
    .B(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__a21o_1 _18067_ (.A1(_01999_),
    .A2(_02014_),
    .B1(_02012_),
    .X(_02115_));
 sky130_fd_sc_hd__or2b_1 _18068_ (.A(_02051_),
    .B_N(_02032_),
    .X(_02116_));
 sky130_fd_sc_hd__or2_1 _18069_ (.A(_08643_),
    .B(_09420_),
    .X(_02117_));
 sky130_fd_sc_hd__or3_1 _18070_ (.A(_10379_),
    .B(_09536_),
    .C(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__o21ai_1 _18071_ (.A1(_10379_),
    .A2(_09536_),
    .B1(_02117_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _18072_ (.A(_02118_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__nor2_1 _18073_ (.A(_10383_),
    .B(_09805_),
    .Y(_02121_));
 sky130_fd_sc_hd__xor2_1 _18074_ (.A(_02120_),
    .B(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__nand2_1 _18075_ (.A(_01989_),
    .B(_01990_),
    .Y(_02123_));
 sky130_fd_sc_hd__o31a_1 _18076_ (.A1(_10257_),
    .A2(_09805_),
    .A3(_01991_),
    .B1(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__xor2_1 _18077_ (.A(_02122_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__and3_1 _18078_ (.A(_10257_),
    .B(net7378),
    .C(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__a21oi_1 _18079_ (.A1(_10257_),
    .A2(net7378),
    .B1(_02125_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _18080_ (.A(_02126_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__a21bo_1 _18081_ (.A1(_02004_),
    .A2(_02005_),
    .B1_N(_02002_),
    .X(_02129_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_02035_),
    .B(_02036_),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _18083_ (.A(_01778_),
    .B(_09249_),
    .Y(_02131_));
 sky130_fd_sc_hd__nor2_1 _18084_ (.A(_09231_),
    .B(_08793_),
    .Y(_02132_));
 sky130_fd_sc_hd__xnor2_1 _18085_ (.A(_02131_),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__or3_1 _18086_ (.A(_01675_),
    .B(_09310_),
    .C(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__o21ai_1 _18087_ (.A1(_01675_),
    .A2(_09310_),
    .B1(_02133_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _18088_ (.A(_02134_),
    .B(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__a21oi_1 _18089_ (.A1(_02130_),
    .A2(_02038_),
    .B1(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__and3_1 _18090_ (.A(_02130_),
    .B(_02038_),
    .C(_02136_),
    .X(_02138_));
 sky130_fd_sc_hd__nor2_1 _18091_ (.A(_02137_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__xnor2_1 _18092_ (.A(_02129_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__a21oi_1 _18093_ (.A1(_02001_),
    .A2(_02009_),
    .B1(_02007_),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_1 _18094_ (.A(_02140_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__and2_1 _18095_ (.A(_02140_),
    .B(_02141_),
    .X(_02143_));
 sky130_fd_sc_hd__nor2_1 _18096_ (.A(_02142_),
    .B(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__xnor2_1 _18097_ (.A(_02128_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__a21oi_1 _18098_ (.A1(_02049_),
    .A2(_02116_),
    .B1(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__and3_1 _18099_ (.A(_02049_),
    .B(_02116_),
    .C(_02145_),
    .X(_02147_));
 sky130_fd_sc_hd__or2_1 _18100_ (.A(_02146_),
    .B(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__xnor2_1 _18101_ (.A(_02115_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(_02114_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__or2_1 _18103_ (.A(_02114_),
    .B(_02149_),
    .X(_02151_));
 sky130_fd_sc_hd__nand2_1 _18104_ (.A(_02150_),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21oi_1 _18105_ (.A1(_02019_),
    .A2(_02057_),
    .B1(_02055_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor2_1 _18106_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__and2_1 _18107_ (.A(_02152_),
    .B(_02153_),
    .X(_02155_));
 sky130_fd_sc_hd__nor2_1 _18108_ (.A(_02154_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__xnor2_1 _18109_ (.A(_02082_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__nor2_1 _18110_ (.A(_02058_),
    .B(_02059_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21oi_2 _18111_ (.A1(_01986_),
    .A2(_02060_),
    .B1(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__xor2_1 _18112_ (.A(_02157_),
    .B(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__xnor2_1 _18113_ (.A(_01984_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _18114_ (.A(_02061_),
    .B(_02062_),
    .Y(_02162_));
 sky130_fd_sc_hd__a21oi_2 _18115_ (.A1(_01874_),
    .A2(_02063_),
    .B1(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__or2_1 _18116_ (.A(_02161_),
    .B(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__nand2_1 _18117_ (.A(_02161_),
    .B(_02163_),
    .Y(_02165_));
 sky130_fd_sc_hd__and2_1 _18118_ (.A(_02164_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__a21o_1 _18119_ (.A1(_01980_),
    .A2(_01981_),
    .B1(_02064_),
    .X(_02167_));
 sky130_fd_sc_hd__a21o_1 _18120_ (.A1(_01965_),
    .A2(_02167_),
    .B1(_02066_),
    .X(_02168_));
 sky130_fd_sc_hd__o31ai_4 _18121_ (.A1(_01967_),
    .A2(_01969_),
    .A3(_02067_),
    .B1(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__a21oi_1 _18122_ (.A1(_02166_),
    .A2(_02169_),
    .B1(net3508),
    .Y(_02170_));
 sky130_fd_sc_hd__o21a_1 _18123_ (.A1(_02166_),
    .A2(_02169_),
    .B1(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__a21o_1 _18124_ (.A1(_09987_),
    .A2(net7815),
    .B1(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_1 _18125_ (.A0(_02172_),
    .A1(net4497),
    .S(_01749_),
    .X(_02173_));
 sky130_fd_sc_hd__clkbuf_1 _18126_ (.A(_02173_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _18127_ (.A(_02157_),
    .B(_02159_),
    .X(_02174_));
 sky130_fd_sc_hd__nand2_1 _18128_ (.A(_01984_),
    .B(_02160_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _18129_ (.A(_01834_),
    .B(_02084_),
    .Y(_02176_));
 sky130_fd_sc_hd__and2b_1 _18130_ (.A_N(_01833_),
    .B(_02084_),
    .X(_02177_));
 sky130_fd_sc_hd__nor2_1 _18131_ (.A(_02176_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__or2b_1 _18132_ (.A(_02098_),
    .B_N(_02106_),
    .X(_02179_));
 sky130_fd_sc_hd__o21a_1 _18133_ (.A1(_02103_),
    .A2(_02105_),
    .B1(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__o21ai_2 _18134_ (.A1(_02023_),
    .A2(_02083_),
    .B1(_02091_),
    .Y(_02181_));
 sky130_fd_sc_hd__or2_1 _18135_ (.A(_10259_),
    .B(_09863_),
    .X(_02182_));
 sky130_fd_sc_hd__nor2_1 _18136_ (.A(_01802_),
    .B(_09732_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_1 _18137_ (.A(_02182_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _18138_ (.A(_08705_),
    .B(_09602_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_1 _18139_ (.A(_02184_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__or2_1 _18140_ (.A(_02184_),
    .B(_02185_),
    .X(_02187_));
 sky130_fd_sc_hd__nand2_1 _18141_ (.A(_02186_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__o31a_1 _18142_ (.A1(_01812_),
    .A2(_10416_),
    .A3(_02101_),
    .B1(_02099_),
    .X(_02189_));
 sky130_fd_sc_hd__a21o_1 _18143_ (.A1(_01684_),
    .A2(_10520_),
    .B1(_01711_),
    .X(_02190_));
 sky130_fd_sc_hd__nor3_1 _18144_ (.A(_01684_),
    .B(_10520_),
    .C(_01711_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _18145_ (.A(_02190_),
    .B(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__nor2_1 _18146_ (.A(_01812_),
    .B(_10539_),
    .Y(_02193_));
 sky130_fd_sc_hd__xnor2_2 _18147_ (.A(_02192_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__xor2_1 _18148_ (.A(_02189_),
    .B(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__xnor2_1 _18149_ (.A(_02188_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _18150_ (.A(_02181_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__or2_1 _18151_ (.A(_02181_),
    .B(_02196_),
    .X(_02198_));
 sky130_fd_sc_hd__nand2_1 _18152_ (.A(_02197_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__xor2_2 _18153_ (.A(_02180_),
    .B(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__xnor2_1 _18154_ (.A(_02178_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__a21o_1 _18155_ (.A1(_02086_),
    .A2(_02110_),
    .B1(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__nand3_1 _18156_ (.A(_02086_),
    .B(_02110_),
    .C(_02201_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _18157_ (.A(_02202_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21o_1 _18158_ (.A1(_02128_),
    .A2(_02144_),
    .B1(_02142_),
    .X(_02205_));
 sky130_fd_sc_hd__or2b_1 _18159_ (.A(_02108_),
    .B_N(_02090_),
    .X(_02206_));
 sky130_fd_sc_hd__a21bo_1 _18160_ (.A1(_02093_),
    .A2(_02107_),
    .B1_N(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__o22a_1 _18161_ (.A1(_08634_),
    .A2(_09420_),
    .B1(_09538_),
    .B2(_08643_),
    .X(_02208_));
 sky130_fd_sc_hd__or3_1 _18162_ (.A(_08634_),
    .B(_09538_),
    .C(_02117_),
    .X(_02209_));
 sky130_fd_sc_hd__or2b_1 _18163_ (.A(_02208_),
    .B_N(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__or3b_1 _18164_ (.A(_09486_),
    .B(_10379_),
    .C_N(net8017),
    .X(_02211_));
 sky130_fd_sc_hd__xnor2_1 _18165_ (.A(_02210_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__o31a_1 _18166_ (.A1(_10383_),
    .A2(_09805_),
    .A3(_02120_),
    .B1(_02118_),
    .X(_02213_));
 sky130_fd_sc_hd__xnor2_1 _18167_ (.A(_02212_),
    .B(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _18168_ (.A(_10383_),
    .B(net7378),
    .Y(_02215_));
 sky130_fd_sc_hd__xnor2_1 _18169_ (.A(_02214_),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21bo_1 _18170_ (.A1(_02131_),
    .A2(_02132_),
    .B1_N(_02134_),
    .X(_02217_));
 sky130_fd_sc_hd__or3_1 _18171_ (.A(_01802_),
    .B(_09602_),
    .C(_02094_),
    .X(_02218_));
 sky130_fd_sc_hd__a21bo_1 _18172_ (.A1(_02096_),
    .A2(_02097_),
    .B1_N(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__nor2_1 _18173_ (.A(_09231_),
    .B(_09249_),
    .Y(_02220_));
 sky130_fd_sc_hd__nor2_1 _18174_ (.A(_08793_),
    .B(_09375_),
    .Y(_02221_));
 sky130_fd_sc_hd__xnor2_1 _18175_ (.A(_02220_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _18176_ (.A(_01778_),
    .B(_09310_),
    .Y(_02223_));
 sky130_fd_sc_hd__xnor2_1 _18177_ (.A(_02222_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _18178_ (.A(_02219_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__or2_1 _18179_ (.A(_02219_),
    .B(_02224_),
    .X(_02226_));
 sky130_fd_sc_hd__and2_1 _18180_ (.A(_02225_),
    .B(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__xnor2_1 _18181_ (.A(_02217_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__a21oi_1 _18182_ (.A1(_02129_),
    .A2(_02139_),
    .B1(_02137_),
    .Y(_02229_));
 sky130_fd_sc_hd__xor2_1 _18183_ (.A(_02228_),
    .B(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__xnor2_1 _18184_ (.A(_02216_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__xor2_1 _18185_ (.A(_02207_),
    .B(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__and2_1 _18186_ (.A(_02205_),
    .B(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__nor2_1 _18187_ (.A(_02205_),
    .B(_02232_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _18188_ (.A(_02233_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__xor2_1 _18189_ (.A(_02204_),
    .B(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__o21a_1 _18190_ (.A1(_02112_),
    .A2(_02113_),
    .B1(_02150_),
    .X(_02237_));
 sky130_fd_sc_hd__xor2_1 _18191_ (.A(_02236_),
    .B(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__and2b_1 _18192_ (.A_N(_02148_),
    .B(_02115_),
    .X(_02239_));
 sky130_fd_sc_hd__o21ba_1 _18193_ (.A1(_02122_),
    .A2(_02124_),
    .B1_N(_02126_),
    .X(_02240_));
 sky130_fd_sc_hd__o21ba_1 _18194_ (.A1(_02146_),
    .A2(_02239_),
    .B1_N(_02240_),
    .X(_02241_));
 sky130_fd_sc_hd__or3b_1 _18195_ (.A(_02146_),
    .B(_02239_),
    .C_N(_02240_),
    .X(_02242_));
 sky130_fd_sc_hd__and2b_1 _18196_ (.A_N(_02241_),
    .B(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__nand2_1 _18197_ (.A(_02238_),
    .B(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__or2_1 _18198_ (.A(_02238_),
    .B(_02243_),
    .X(_02245_));
 sky130_fd_sc_hd__nand2_1 _18199_ (.A(_02244_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21oi_1 _18200_ (.A1(_02082_),
    .A2(_02156_),
    .B1(_02154_),
    .Y(_02247_));
 sky130_fd_sc_hd__xor2_1 _18201_ (.A(_02246_),
    .B(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__xnor2_1 _18202_ (.A(_02080_),
    .B(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__a21oi_1 _18203_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__and3_1 _18204_ (.A(_02174_),
    .B(_02175_),
    .C(_02249_),
    .X(_02251_));
 sky130_fd_sc_hd__nor2_1 _18205_ (.A(_02250_),
    .B(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__a21bo_1 _18206_ (.A1(_02166_),
    .A2(_02169_),
    .B1_N(_02164_),
    .X(_02253_));
 sky130_fd_sc_hd__or2_1 _18207_ (.A(_02252_),
    .B(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__a21oi_2 _18208_ (.A1(_02252_),
    .A2(_02253_),
    .B1(_09999_),
    .Y(_02255_));
 sky130_fd_sc_hd__nand2_1 _18209_ (.A(net3780),
    .B(net4605),
    .Y(_02256_));
 sky130_fd_sc_hd__or2_1 _18210_ (.A(net3780),
    .B(net4605),
    .X(_02257_));
 sky130_fd_sc_hd__nand2_1 _18211_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__a21bo_1 _18212_ (.A1(_02073_),
    .A2(_02076_),
    .B1_N(_02074_),
    .X(_02259_));
 sky130_fd_sc_hd__xnor2_1 _18213_ (.A(_02258_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__clkbuf_8 _18214_ (.A(net3508),
    .X(_02261_));
 sky130_fd_sc_hd__a22o_1 _18215_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02260_),
    .B2(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_2 _18216_ (.A0(_02262_),
    .A1(net3780),
    .S(_01749_),
    .X(_02263_));
 sky130_fd_sc_hd__clkbuf_1 _18217_ (.A(_02263_),
    .X(_00548_));
 sky130_fd_sc_hd__a21bo_1 _18218_ (.A1(_02257_),
    .A2(_02259_),
    .B1_N(_02256_),
    .X(_02264_));
 sky130_fd_sc_hd__xor2_1 _18219_ (.A(net4577),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__nor2_1 _18220_ (.A(net4575),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__a21o_1 _18221_ (.A1(net4575),
    .A2(_02265_),
    .B1(_01870_),
    .X(_02267_));
 sky130_fd_sc_hd__a21o_1 _18222_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_02249_),
    .X(_02268_));
 sky130_fd_sc_hd__a21oi_1 _18223_ (.A1(_02164_),
    .A2(_02268_),
    .B1(_02251_),
    .Y(_02269_));
 sky130_fd_sc_hd__a31o_1 _18224_ (.A1(_02166_),
    .A2(_02169_),
    .A3(_02252_),
    .B1(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__nor2_1 _18225_ (.A(_02246_),
    .B(_02247_),
    .Y(_02271_));
 sky130_fd_sc_hd__a21oi_1 _18226_ (.A1(_02080_),
    .A2(_02248_),
    .B1(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__o22a_1 _18227_ (.A1(_02212_),
    .A2(_02213_),
    .B1(_02214_),
    .B2(_02215_),
    .X(_02273_));
 sky130_fd_sc_hd__xnor2_1 _18228_ (.A(_02272_),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__o21a_1 _18229_ (.A1(_02236_),
    .A2(_02237_),
    .B1(_02244_),
    .X(_02275_));
 sky130_fd_sc_hd__o21bai_1 _18230_ (.A1(_02190_),
    .A2(_02193_),
    .B1_N(_02191_),
    .Y(_02276_));
 sky130_fd_sc_hd__a21oi_1 _18231_ (.A1(_02207_),
    .A2(_02231_),
    .B1(_02233_),
    .Y(_02277_));
 sky130_fd_sc_hd__o31a_1 _18232_ (.A1(_02204_),
    .A2(_02233_),
    .A3(_02234_),
    .B1(_02202_),
    .X(_02278_));
 sky130_fd_sc_hd__xnor2_1 _18233_ (.A(_02277_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__xnor2_1 _18234_ (.A(_02276_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__o21ba_1 _18235_ (.A1(_02176_),
    .A2(_02200_),
    .B1_N(_02177_),
    .X(_02281_));
 sky130_fd_sc_hd__xnor2_1 _18236_ (.A(_02181_),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__and2_1 _18237_ (.A(_02189_),
    .B(_02194_),
    .X(_02283_));
 sky130_fd_sc_hd__or2_1 _18238_ (.A(_02189_),
    .B(_02194_),
    .X(_02284_));
 sky130_fd_sc_hd__o21a_1 _18239_ (.A1(_02188_),
    .A2(_02283_),
    .B1(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__nor2_1 _18240_ (.A(_08705_),
    .B(_09732_),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _18241_ (.A(_02285_),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__or2b_1 _18242_ (.A(_02216_),
    .B_N(_02230_),
    .X(_02288_));
 sky130_fd_sc_hd__o21a_1 _18243_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__nor2_1 _18244_ (.A(_08540_),
    .B(_09784_),
    .Y(_02290_));
 sky130_fd_sc_hd__xnor2_1 _18245_ (.A(_02289_),
    .B(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__nor2_1 _18246_ (.A(_09375_),
    .B(_09249_),
    .Y(_02292_));
 sky130_fd_sc_hd__a21bo_1 _18247_ (.A1(_02217_),
    .A2(_02227_),
    .B1_N(_02225_),
    .X(_02293_));
 sky130_fd_sc_hd__xor2_1 _18248_ (.A(_02292_),
    .B(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__xnor2_1 _18249_ (.A(_02291_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__o31a_1 _18250_ (.A1(_01802_),
    .A2(_09732_),
    .A3(_02182_),
    .B1(_02186_),
    .X(_02296_));
 sky130_fd_sc_hd__nand2_1 _18251_ (.A(_02220_),
    .B(_02221_),
    .Y(_02297_));
 sky130_fd_sc_hd__o31a_1 _18252_ (.A1(_01778_),
    .A2(_09310_),
    .A3(_02222_),
    .B1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__or2_1 _18253_ (.A(_09231_),
    .B(_09310_),
    .X(_02299_));
 sky130_fd_sc_hd__xnor2_1 _18254_ (.A(_02298_),
    .B(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _18255_ (.A(_02181_),
    .B(_02196_),
    .Y(_02301_));
 sky130_fd_sc_hd__o21ai_2 _18256_ (.A1(_02180_),
    .A2(_02301_),
    .B1(_02197_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _18257_ (.A(_08634_),
    .B(_09538_),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _18258_ (.A(_01778_),
    .B(_09418_),
    .Y(_02304_));
 sky130_fd_sc_hd__xnor2_1 _18259_ (.A(_02303_),
    .B(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__xnor2_1 _18260_ (.A(_02302_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__o21a_1 _18261_ (.A1(_02208_),
    .A2(_02211_),
    .B1(_02209_),
    .X(_02307_));
 sky130_fd_sc_hd__nor2_1 _18262_ (.A(_08643_),
    .B(_09805_),
    .Y(_02308_));
 sky130_fd_sc_hd__xnor2_1 _18263_ (.A(_02307_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__xnor2_1 _18264_ (.A(_02306_),
    .B(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__xnor2_1 _18265_ (.A(_02300_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__xnor2_1 _18266_ (.A(_02296_),
    .B(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _18267_ (.A(_08793_),
    .B(_09602_),
    .Y(_02313_));
 sky130_fd_sc_hd__xnor2_1 _18268_ (.A(_02312_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__xnor2_1 _18269_ (.A(_02295_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _18270_ (.A(_01812_),
    .B(_01711_),
    .Y(_02316_));
 sky130_fd_sc_hd__nor2_1 _18271_ (.A(_01802_),
    .B(_09863_),
    .Y(_02317_));
 sky130_fd_sc_hd__nor2_1 _18272_ (.A(_10259_),
    .B(_10172_),
    .Y(_02318_));
 sky130_fd_sc_hd__xnor2_1 _18273_ (.A(_02317_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__xnor2_1 _18274_ (.A(_02316_),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__xnor2_1 _18275_ (.A(_02315_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_1 _18276_ (.A(_02287_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__xnor2_1 _18277_ (.A(_02282_),
    .B(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__xnor2_1 _18278_ (.A(_02241_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _18279_ (.A(_02280_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__xnor2_1 _18280_ (.A(_02275_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand2_1 _18281_ (.A(_02274_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__or2_1 _18282_ (.A(_02274_),
    .B(_02326_),
    .X(_02328_));
 sky130_fd_sc_hd__and2_1 _18283_ (.A(_02327_),
    .B(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__a311oi_1 _18284_ (.A1(_02166_),
    .A2(_02169_),
    .A3(_02252_),
    .B1(_02269_),
    .C1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__a311o_1 _18285_ (.A1(_02270_),
    .A2(_02327_),
    .A3(_02328_),
    .B1(_02330_),
    .C1(_09999_),
    .X(_02331_));
 sky130_fd_sc_hd__o21ai_1 _18286_ (.A1(_02266_),
    .A2(_02267_),
    .B1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__mux2_4 _18287_ (.A0(_02332_),
    .A1(net4577),
    .S(_01749_),
    .X(_02333_));
 sky130_fd_sc_hd__clkbuf_1 _18288_ (.A(_02333_),
    .X(_00549_));
 sky130_fd_sc_hd__nand2_1 _18289_ (.A(net4475),
    .B(net4315),
    .Y(_02334_));
 sky130_fd_sc_hd__or2_1 _18290_ (.A(net4475),
    .B(net4315),
    .X(_02335_));
 sky130_fd_sc_hd__a31o_1 _18291_ (.A1(_09987_),
    .A2(_02334_),
    .A3(_02335_),
    .B1(_09992_),
    .X(_02336_));
 sky130_fd_sc_hd__a211o_1 _18292_ (.A1(_06204_),
    .A2(_08314_),
    .B1(_06388_),
    .C1(net4919),
    .X(_02337_));
 sky130_fd_sc_hd__buf_4 _18293_ (.A(net4920),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _18294_ (.A0(_02336_),
    .A1(net4475),
    .S(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__clkbuf_1 _18295_ (.A(_02339_),
    .X(_00550_));
 sky130_fd_sc_hd__nand2_1 _18296_ (.A(net4467),
    .B(net4310),
    .Y(_02340_));
 sky130_fd_sc_hd__or2_1 _18297_ (.A(net4467),
    .B(net4310),
    .X(_02341_));
 sky130_fd_sc_hd__nand2_1 _18298_ (.A(_02340_),
    .B(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__xnor2_1 _18299_ (.A(_02334_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__o21ai_1 _18300_ (.A1(_06206_),
    .A2(net7793),
    .B1(_10002_),
    .Y(_02344_));
 sky130_fd_sc_hd__mux2_1 _18301_ (.A0(_02344_),
    .A1(net4467),
    .S(_02338_),
    .X(_02345_));
 sky130_fd_sc_hd__clkbuf_1 _18302_ (.A(_02345_),
    .X(_00551_));
 sky130_fd_sc_hd__o21a_1 _18303_ (.A1(_02334_),
    .A2(_02342_),
    .B1(_02340_),
    .X(_02346_));
 sky130_fd_sc_hd__nor2_1 _18304_ (.A(net4687),
    .B(net4455),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _18305_ (.A(net4687),
    .B(net4455),
    .Y(_02348_));
 sky130_fd_sc_hd__or2b_1 _18306_ (.A(_02347_),
    .B_N(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__xnor2_1 _18307_ (.A(_02346_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__o21ai_1 _18308_ (.A1(_06206_),
    .A2(net7805),
    .B1(_10011_),
    .Y(_02351_));
 sky130_fd_sc_hd__mux2_1 _18309_ (.A0(_02351_),
    .A1(net4687),
    .S(_02338_),
    .X(_02352_));
 sky130_fd_sc_hd__clkbuf_1 _18310_ (.A(_02352_),
    .X(_00552_));
 sky130_fd_sc_hd__o21a_1 _18311_ (.A1(_02346_),
    .A2(_02347_),
    .B1(_02348_),
    .X(_02353_));
 sky130_fd_sc_hd__nor2_1 _18312_ (.A(net4499),
    .B(net4435),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _18313_ (.A(net4499),
    .B(net4435),
    .Y(_02355_));
 sky130_fd_sc_hd__or2b_1 _18314_ (.A(_02354_),
    .B_N(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__nor2_1 _18315_ (.A(_02353_),
    .B(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__a21o_1 _18316_ (.A1(_02353_),
    .A2(_02356_),
    .B1(_01870_),
    .X(_02358_));
 sky130_fd_sc_hd__o21ai_1 _18317_ (.A1(_02357_),
    .A2(_02358_),
    .B1(_10021_),
    .Y(_02359_));
 sky130_fd_sc_hd__mux2_1 _18318_ (.A0(_02359_),
    .A1(net4499),
    .S(_02338_),
    .X(_02360_));
 sky130_fd_sc_hd__clkbuf_1 _18319_ (.A(_02360_),
    .X(_00553_));
 sky130_fd_sc_hd__or2_1 _18320_ (.A(net4591),
    .B(net4382),
    .X(_02361_));
 sky130_fd_sc_hd__nand2_1 _18321_ (.A(net4591),
    .B(net4382),
    .Y(_02362_));
 sky130_fd_sc_hd__o21ai_2 _18322_ (.A1(_02353_),
    .A2(_02354_),
    .B1(_02355_),
    .Y(_02363_));
 sky130_fd_sc_hd__a21oi_1 _18323_ (.A1(_02361_),
    .A2(_02362_),
    .B1(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__a31o_1 _18324_ (.A1(_02363_),
    .A2(_02361_),
    .A3(_02362_),
    .B1(_06205_),
    .X(_02365_));
 sky130_fd_sc_hd__o21ai_1 _18325_ (.A1(net7782),
    .A2(_02365_),
    .B1(_10029_),
    .Y(_02366_));
 sky130_fd_sc_hd__mux2_1 _18326_ (.A0(_02366_),
    .A1(net4591),
    .S(_02338_),
    .X(_02367_));
 sky130_fd_sc_hd__clkbuf_1 _18327_ (.A(_02367_),
    .X(_00554_));
 sky130_fd_sc_hd__a21boi_2 _18328_ (.A1(_02363_),
    .A2(_02361_),
    .B1_N(_02362_),
    .Y(_02368_));
 sky130_fd_sc_hd__nor2_1 _18329_ (.A(net4511),
    .B(net4374),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_1 _18330_ (.A(net4511),
    .B(net4374),
    .Y(_02370_));
 sky130_fd_sc_hd__or2b_1 _18331_ (.A(_02369_),
    .B_N(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__xnor2_1 _18332_ (.A(_02368_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__o21ai_1 _18333_ (.A1(_10010_),
    .A2(_02372_),
    .B1(_10037_),
    .Y(_02373_));
 sky130_fd_sc_hd__mux2_1 _18334_ (.A0(_02373_),
    .A1(net4511),
    .S(_02338_),
    .X(_02374_));
 sky130_fd_sc_hd__clkbuf_1 _18335_ (.A(_02374_),
    .X(_00555_));
 sky130_fd_sc_hd__o21a_1 _18336_ (.A1(_02368_),
    .A2(_02369_),
    .B1(_02370_),
    .X(_02375_));
 sky130_fd_sc_hd__nor2_1 _18337_ (.A(net4491),
    .B(net4473),
    .Y(_02376_));
 sky130_fd_sc_hd__nand2_1 _18338_ (.A(net4491),
    .B(net4473),
    .Y(_02377_));
 sky130_fd_sc_hd__or2b_1 _18339_ (.A(_02376_),
    .B_N(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__nor2_1 _18340_ (.A(_02375_),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21o_1 _18341_ (.A1(_02375_),
    .A2(_02378_),
    .B1(_01870_),
    .X(_02380_));
 sky130_fd_sc_hd__o21ai_1 _18342_ (.A1(net7818),
    .A2(_02380_),
    .B1(_10047_),
    .Y(_02381_));
 sky130_fd_sc_hd__mux2_1 _18343_ (.A0(_02381_),
    .A1(net4491),
    .S(_02338_),
    .X(_02382_));
 sky130_fd_sc_hd__clkbuf_1 _18344_ (.A(_02382_),
    .X(_00556_));
 sky130_fd_sc_hd__o21a_1 _18345_ (.A1(_02375_),
    .A2(_02376_),
    .B1(_02377_),
    .X(_02383_));
 sky130_fd_sc_hd__nor2_1 _18346_ (.A(net4485),
    .B(net4353),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(net4485),
    .B(net4353),
    .Y(_02385_));
 sky130_fd_sc_hd__or2b_1 _18348_ (.A(_02384_),
    .B_N(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__xnor2_1 _18349_ (.A(_02383_),
    .B(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__o21ai_1 _18350_ (.A1(_10010_),
    .A2(_02387_),
    .B1(_10055_),
    .Y(_02388_));
 sky130_fd_sc_hd__mux2_1 _18351_ (.A0(_02388_),
    .A1(net4485),
    .S(_02338_),
    .X(_02389_));
 sky130_fd_sc_hd__clkbuf_1 _18352_ (.A(_02389_),
    .X(_00557_));
 sky130_fd_sc_hd__o21a_1 _18353_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02385_),
    .X(_02390_));
 sky130_fd_sc_hd__nor2_1 _18354_ (.A(net4453),
    .B(net3505),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_1 _18355_ (.A(net4453),
    .B(net3505),
    .Y(_02392_));
 sky130_fd_sc_hd__or2b_1 _18356_ (.A(_02391_),
    .B_N(net3393),
    .X(_02393_));
 sky130_fd_sc_hd__nor2_1 _18357_ (.A(net7801),
    .B(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__a21o_1 _18358_ (.A1(_02390_),
    .A2(_02393_),
    .B1(_01870_),
    .X(_02395_));
 sky130_fd_sc_hd__o21ai_1 _18359_ (.A1(_02394_),
    .A2(_02395_),
    .B1(_10064_),
    .Y(_02396_));
 sky130_fd_sc_hd__mux2_1 _18360_ (.A0(_02396_),
    .A1(net4453),
    .S(_02338_),
    .X(_02397_));
 sky130_fd_sc_hd__clkbuf_1 _18361_ (.A(_02397_),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _18362_ (.A(net4489),
    .B(net4393),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_1 _18363_ (.A(net4489),
    .B(net4393),
    .Y(_02399_));
 sky130_fd_sc_hd__o21ai_1 _18364_ (.A1(_02390_),
    .A2(_02391_),
    .B1(net3393),
    .Y(_02400_));
 sky130_fd_sc_hd__a21oi_1 _18365_ (.A1(_02398_),
    .A2(_02399_),
    .B1(net3394),
    .Y(_02401_));
 sky130_fd_sc_hd__a31o_1 _18366_ (.A1(net3394),
    .A2(_02398_),
    .A3(_02399_),
    .B1(_06205_),
    .X(_02402_));
 sky130_fd_sc_hd__o21ai_1 _18367_ (.A1(_02401_),
    .A2(_02402_),
    .B1(_10072_),
    .Y(_02403_));
 sky130_fd_sc_hd__mux2_1 _18368_ (.A0(_02403_),
    .A1(net4489),
    .S(_02338_),
    .X(_02404_));
 sky130_fd_sc_hd__clkbuf_1 _18369_ (.A(_02404_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_1 _18370_ (.A(net3394),
    .B(_02398_),
    .Y(_02405_));
 sky130_fd_sc_hd__and2_1 _18371_ (.A(net4538),
    .B(net4405),
    .X(_02406_));
 sky130_fd_sc_hd__nor2_1 _18372_ (.A(net4538),
    .B(net4405),
    .Y(_02407_));
 sky130_fd_sc_hd__a211oi_1 _18373_ (.A1(_02399_),
    .A2(net3395),
    .B1(net3234),
    .C1(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__o211a_1 _18374_ (.A1(_02407_),
    .A2(net3234),
    .B1(net3395),
    .C1(_02399_),
    .X(_02409_));
 sky130_fd_sc_hd__o31ai_1 _18375_ (.A1(_10010_),
    .A2(net3396),
    .A3(_02409_),
    .B1(_10080_),
    .Y(_02410_));
 sky130_fd_sc_hd__buf_4 _18376_ (.A(net4920),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _18377_ (.A0(_02410_),
    .A1(net4538),
    .S(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__clkbuf_1 _18378_ (.A(_02412_),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _18379_ (.A(net4429),
    .B(net4451),
    .X(_02413_));
 sky130_fd_sc_hd__nand2_1 _18380_ (.A(net4429),
    .B(net4451),
    .Y(_02414_));
 sky130_fd_sc_hd__a211o_1 _18381_ (.A1(_02413_),
    .A2(_02414_),
    .B1(net3234),
    .C1(net3396),
    .X(_02415_));
 sky130_fd_sc_hd__o211ai_1 _18382_ (.A1(net3234),
    .A2(net3396),
    .B1(_02413_),
    .C1(_02414_),
    .Y(_02416_));
 sky130_fd_sc_hd__a31o_1 _18383_ (.A1(_09987_),
    .A2(_02415_),
    .A3(net3235),
    .B1(_10206_),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _18384_ (.A0(_02417_),
    .A1(net4429),
    .S(_02411_),
    .X(_02418_));
 sky130_fd_sc_hd__clkbuf_1 _18385_ (.A(_02418_),
    .X(_00561_));
 sky130_fd_sc_hd__and2_1 _18386_ (.A(net4536),
    .B(net4372),
    .X(_02419_));
 sky130_fd_sc_hd__nor2_1 _18387_ (.A(net4536),
    .B(net4372),
    .Y(_02420_));
 sky130_fd_sc_hd__a211o_1 _18388_ (.A1(_02414_),
    .A2(net3235),
    .B1(_02419_),
    .C1(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__o211ai_1 _18389_ (.A1(_02419_),
    .A2(_02420_),
    .B1(_02414_),
    .C1(net3235),
    .Y(_02422_));
 sky130_fd_sc_hd__a31o_1 _18390_ (.A1(_09987_),
    .A2(_02421_),
    .A3(net3236),
    .B1(_10330_),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _18391_ (.A0(_02423_),
    .A1(net4536),
    .S(_02411_),
    .X(_02424_));
 sky130_fd_sc_hd__clkbuf_1 _18392_ (.A(_02424_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _18393_ (.A(net4487),
    .B(net4423),
    .Y(_02425_));
 sky130_fd_sc_hd__or2_1 _18394_ (.A(net4487),
    .B(net4423),
    .X(_02426_));
 sky130_fd_sc_hd__inv_2 _18395_ (.A(_02421_),
    .Y(_02427_));
 sky130_fd_sc_hd__a211o_1 _18396_ (.A1(_02425_),
    .A2(_02426_),
    .B1(_02419_),
    .C1(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__o211ai_2 _18397_ (.A1(_02419_),
    .A2(_02427_),
    .B1(_02425_),
    .C1(_02426_),
    .Y(_02429_));
 sky130_fd_sc_hd__a31o_1 _18398_ (.A1(_02261_),
    .A2(_02428_),
    .A3(_02429_),
    .B1(_10455_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _18399_ (.A0(_02430_),
    .A1(net4487),
    .S(_02411_),
    .X(_02431_));
 sky130_fd_sc_hd__clkbuf_1 _18400_ (.A(_02431_),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _18401_ (.A(net4613),
    .B(net4378),
    .X(_02432_));
 sky130_fd_sc_hd__nor2_1 _18402_ (.A(net4613),
    .B(net4378),
    .Y(_02433_));
 sky130_fd_sc_hd__a211oi_1 _18403_ (.A1(_02425_),
    .A2(_02429_),
    .B1(_02432_),
    .C1(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__o211a_1 _18404_ (.A1(_02432_),
    .A2(_02433_),
    .B1(_02425_),
    .C1(_02429_),
    .X(_02435_));
 sky130_fd_sc_hd__o31ai_1 _18405_ (.A1(_10010_),
    .A2(_02434_),
    .A3(_02435_),
    .B1(_10571_),
    .Y(_02436_));
 sky130_fd_sc_hd__mux2_1 _18406_ (.A0(_02436_),
    .A1(net4613),
    .S(_02411_),
    .X(_02437_));
 sky130_fd_sc_hd__clkbuf_1 _18407_ (.A(_02437_),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _18408_ (.A(net4458),
    .B(net5684),
    .Y(_02438_));
 sky130_fd_sc_hd__or2_1 _18409_ (.A(net4458),
    .B(net5684),
    .X(_02439_));
 sky130_fd_sc_hd__nand2_1 _18410_ (.A(_02438_),
    .B(_02439_),
    .Y(_02440_));
 sky130_fd_sc_hd__nor2_1 _18411_ (.A(_02432_),
    .B(_02434_),
    .Y(_02441_));
 sky130_fd_sc_hd__xnor2_1 _18412_ (.A(_02440_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__o21ai_1 _18413_ (.A1(_10010_),
    .A2(_02442_),
    .B1(_01747_),
    .Y(_02443_));
 sky130_fd_sc_hd__mux2_1 _18414_ (.A0(_02443_),
    .A1(net4458),
    .S(_02411_),
    .X(_02444_));
 sky130_fd_sc_hd__clkbuf_1 _18415_ (.A(_02444_),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _18416_ (.A(net4483),
    .B(net4368),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _18417_ (.A(net4483),
    .B(net4368),
    .Y(_02446_));
 sky130_fd_sc_hd__or2b_1 _18418_ (.A(_02445_),
    .B_N(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__o21a_1 _18419_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02438_),
    .X(_02448_));
 sky130_fd_sc_hd__xnor2_1 _18420_ (.A(_02447_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__o21ai_1 _18421_ (.A1(_10010_),
    .A2(_02449_),
    .B1(_01862_),
    .Y(_02450_));
 sky130_fd_sc_hd__mux2_1 _18422_ (.A0(_02450_),
    .A1(net4483),
    .S(_02411_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _18423_ (.A(_02451_),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _18424_ (.A(net4573),
    .B(net4386),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_1 _18425_ (.A(net4573),
    .B(net4386),
    .Y(_02453_));
 sky130_fd_sc_hd__or2b_1 _18426_ (.A(_02452_),
    .B_N(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__o21a_1 _18427_ (.A1(_02445_),
    .A2(_02448_),
    .B1(_02446_),
    .X(_02455_));
 sky130_fd_sc_hd__nor2_1 _18428_ (.A(_02454_),
    .B(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__a21o_1 _18429_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_01870_),
    .X(_02457_));
 sky130_fd_sc_hd__o21ai_1 _18430_ (.A1(_02456_),
    .A2(_02457_),
    .B1(_01971_),
    .Y(_02458_));
 sky130_fd_sc_hd__mux2_1 _18431_ (.A0(_02458_),
    .A1(net4573),
    .S(_02411_),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_1 _18432_ (.A(_02459_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _18433_ (.A(net4513),
    .B(net4431),
    .Y(_02460_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(net4513),
    .B(net4431),
    .Y(_02461_));
 sky130_fd_sc_hd__or2b_1 _18435_ (.A(_02460_),
    .B_N(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__o21a_1 _18436_ (.A1(_02452_),
    .A2(_02455_),
    .B1(_02453_),
    .X(_02463_));
 sky130_fd_sc_hd__nor2_1 _18437_ (.A(_02462_),
    .B(net7789),
    .Y(_02464_));
 sky130_fd_sc_hd__a21o_1 _18438_ (.A1(_02462_),
    .A2(_02463_),
    .B1(_01870_),
    .X(_02465_));
 sky130_fd_sc_hd__o21ai_1 _18439_ (.A1(net7790),
    .A2(_02465_),
    .B1(_02070_),
    .Y(_02466_));
 sky130_fd_sc_hd__mux2_1 _18440_ (.A0(_02466_),
    .A1(net4513),
    .S(_02411_),
    .X(_02467_));
 sky130_fd_sc_hd__clkbuf_1 _18441_ (.A(_02467_),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _18442_ (.A(net4437),
    .B(net4380),
    .X(_02468_));
 sky130_fd_sc_hd__nand2_1 _18443_ (.A(net4437),
    .B(net4380),
    .Y(_02469_));
 sky130_fd_sc_hd__nand2_1 _18444_ (.A(_02468_),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__o21ai_1 _18445_ (.A1(_02460_),
    .A2(_02463_),
    .B1(_02461_),
    .Y(_02471_));
 sky130_fd_sc_hd__xnor2_1 _18446_ (.A(_02470_),
    .B(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__a21o_1 _18447_ (.A1(_09987_),
    .A2(_02472_),
    .B1(_02171_),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _18448_ (.A0(_02473_),
    .A1(net4437),
    .S(_02411_),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_1 _18449_ (.A(_02474_),
    .X(_00569_));
 sky130_fd_sc_hd__nand2_1 _18450_ (.A(net3742),
    .B(net4586),
    .Y(_02475_));
 sky130_fd_sc_hd__or2_1 _18451_ (.A(net3742),
    .B(net4586),
    .X(_02476_));
 sky130_fd_sc_hd__nand2_1 _18452_ (.A(net3059),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__a21bo_1 _18453_ (.A1(_02468_),
    .A2(_02471_),
    .B1_N(_02469_),
    .X(_02478_));
 sky130_fd_sc_hd__xnor2_1 _18454_ (.A(_02477_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__a22o_1 _18455_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02479_),
    .B2(_02261_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_2 _18456_ (.A0(_02480_),
    .A1(net3742),
    .S(net4920),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_1 _18457_ (.A(_02481_),
    .X(_00570_));
 sky130_fd_sc_hd__a21bo_1 _18458_ (.A1(_02476_),
    .A2(_02478_),
    .B1_N(net3059),
    .X(_02482_));
 sky130_fd_sc_hd__xnor2_1 _18459_ (.A(_06269_),
    .B(net3060),
    .Y(_02483_));
 sky130_fd_sc_hd__nor2_1 _18460_ (.A(net4332),
    .B(net3061),
    .Y(_02484_));
 sky130_fd_sc_hd__a21o_1 _18461_ (.A1(net4332),
    .A2(net3061),
    .B1(_01870_),
    .X(_02485_));
 sky130_fd_sc_hd__o21ai_1 _18462_ (.A1(net3062),
    .A2(_02485_),
    .B1(_02331_),
    .Y(_02486_));
 sky130_fd_sc_hd__mux2_4 _18463_ (.A0(_02486_),
    .A1(net4342),
    .S(net4920),
    .X(_02487_));
 sky130_fd_sc_hd__clkbuf_1 _18464_ (.A(_02487_),
    .X(_00571_));
 sky130_fd_sc_hd__buf_4 _18465_ (.A(_08274_),
    .X(_02488_));
 sky130_fd_sc_hd__and2_1 _18466_ (.A(net43),
    .B(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__clkbuf_1 _18467_ (.A(_02489_),
    .X(_00572_));
 sky130_fd_sc_hd__and2_1 _18468_ (.A(net7205),
    .B(_02488_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _18469_ (.A(net1212),
    .X(_00573_));
 sky130_fd_sc_hd__buf_2 _18470_ (.A(net4326),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_4 _18471_ (.A(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _18472_ (.A(net3074),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _18473_ (.A(net3150),
    .X(_02494_));
 sky130_fd_sc_hd__and2_2 _18474_ (.A(net3075),
    .B(net3151),
    .X(_02495_));
 sky130_fd_sc_hd__and2b_1 _18475_ (.A_N(net3925),
    .B(net3960),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_4 _18476_ (.A(net7315),
    .X(_02497_));
 sky130_fd_sc_hd__nor2_4 _18477_ (.A(net3074),
    .B(net3150),
    .Y(_02498_));
 sky130_fd_sc_hd__nand2_1 _18478_ (.A(_02497_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__and2b_2 _18479_ (.A_N(net3151),
    .B(net3074),
    .X(_02500_));
 sky130_fd_sc_hd__nand2_1 _18480_ (.A(net3074),
    .B(net3150),
    .Y(_02501_));
 sky130_fd_sc_hd__mux2_1 _18481_ (.A0(net7360),
    .A1(\rbzero.spi_registers.spi_cmd[2] ),
    .S(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__nand2_1 _18482_ (.A(_02499_),
    .B(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__a21o_1 _18483_ (.A1(_02497_),
    .A2(_02500_),
    .B1(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__o311a_1 _18484_ (.A1(net3925),
    .A2(net3960),
    .A3(_02495_),
    .B1(_02499_),
    .C1(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__xor2_1 _18485_ (.A(net3889),
    .B(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__nor2_1 _18486_ (.A(net3925),
    .B(net3960),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_02495_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__a21oi_1 _18488_ (.A1(_02504_),
    .A2(_02508_),
    .B1(net3211),
    .Y(_02509_));
 sky130_fd_sc_hd__or2_1 _18489_ (.A(net3747),
    .B(_02504_),
    .X(_02510_));
 sky130_fd_sc_hd__nand2_1 _18490_ (.A(net3747),
    .B(_02504_),
    .Y(_02511_));
 sky130_fd_sc_hd__a32o_1 _18491_ (.A1(net3211),
    .A2(_02504_),
    .A3(_02508_),
    .B1(_02510_),
    .B2(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__xor2_1 _18492_ (.A(net3904),
    .B(_02503_),
    .X(_02513_));
 sky130_fd_sc_hd__and2b_1 _18493_ (.A_N(net3960),
    .B(net3925),
    .X(_02514_));
 sky130_fd_sc_hd__and2_1 _18494_ (.A(_02501_),
    .B(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__a21oi_1 _18495_ (.A1(net3075),
    .A2(_02497_),
    .B1(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__xnor2_1 _18496_ (.A(net3885),
    .B(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__or3_1 _18497_ (.A(net3885),
    .B(net3904),
    .C(net3913),
    .X(_02518_));
 sky130_fd_sc_hd__nor3_1 _18498_ (.A(net1296),
    .B(net3969),
    .C(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__or3_1 _18499_ (.A(net1296),
    .B(net3374),
    .C(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__or3_1 _18500_ (.A(_02513_),
    .B(_02517_),
    .C(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__or4_1 _18501_ (.A(_02506_),
    .B(net3212),
    .C(_02512_),
    .D(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__nor2_1 _18502_ (.A(net3945),
    .B(_04241_),
    .Y(_02523_));
 sky130_fd_sc_hd__and2b_1 _18503_ (.A_N(net2977),
    .B(net1577),
    .X(_02524_));
 sky130_fd_sc_hd__and4bb_1 _18504_ (.A_N(_02492_),
    .B_N(net3213),
    .C(_02523_),
    .D(net2978),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_1 _18505_ (.A(net3214),
    .X(_00574_));
 sky130_fd_sc_hd__and2_1 _18506_ (.A(net44),
    .B(_02488_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _18507_ (.A(_02526_),
    .X(_00575_));
 sky130_fd_sc_hd__and2_2 _18508_ (.A(net6328),
    .B(_02488_),
    .X(_02527_));
 sky130_fd_sc_hd__clkbuf_1 _18509_ (.A(net628),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_4 _18510_ (.A(_09932_),
    .X(_02528_));
 sky130_fd_sc_hd__clkbuf_4 _18511_ (.A(_09935_),
    .X(_02529_));
 sky130_fd_sc_hd__nor2_1 _18512_ (.A(net4493),
    .B(net4791),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _18513_ (.A(net4446),
    .B(net4806),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _18514_ (.A(_05403_),
    .B(net715),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _18515_ (.A(net4424),
    .B(net701),
    .Y(_02533_));
 sky130_fd_sc_hd__or2_1 _18516_ (.A(net4656),
    .B(net715),
    .X(_02534_));
 sky130_fd_sc_hd__nand3b_1 _18517_ (.A_N(net4425),
    .B(net4657),
    .C(_02532_),
    .Y(_02535_));
 sky130_fd_sc_hd__and2_1 _18518_ (.A(_02532_),
    .B(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__nand2_1 _18519_ (.A(net4446),
    .B(net4806),
    .Y(_02537_));
 sky130_fd_sc_hd__o21a_1 _18520_ (.A1(_02531_),
    .A2(_02536_),
    .B1(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__nand2_1 _18521_ (.A(net4476),
    .B(net908),
    .Y(_02539_));
 sky130_fd_sc_hd__o21a_1 _18522_ (.A1(_02530_),
    .A2(_02538_),
    .B1(net4477),
    .X(_02540_));
 sky130_fd_sc_hd__nor2_1 _18523_ (.A(net3837),
    .B(net1076),
    .Y(_02541_));
 sky130_fd_sc_hd__nand2_1 _18524_ (.A(net3838),
    .B(net1076),
    .Y(_02542_));
 sky130_fd_sc_hd__or2b_1 _18525_ (.A(_02541_),
    .B_N(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__xor2_1 _18526_ (.A(net4478),
    .B(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__inv_2 _18527_ (.A(net4424),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _18528_ (.A(_02545_),
    .B(_08195_),
    .Y(_02546_));
 sky130_fd_sc_hd__a221o_1 _18529_ (.A1(net1076),
    .A2(_02528_),
    .B1(_02529_),
    .B2(net4479),
    .C1(_02546_),
    .X(_00577_));
 sky130_fd_sc_hd__nand2_1 _18530_ (.A(_05403_),
    .B(net4424),
    .Y(_02547_));
 sky130_fd_sc_hd__or2_1 _18531_ (.A(_05403_),
    .B(net4424),
    .X(_02548_));
 sky130_fd_sc_hd__o21a_1 _18532_ (.A1(net4478),
    .A2(_02541_),
    .B1(_02542_),
    .X(_02549_));
 sky130_fd_sc_hd__nor2_1 _18533_ (.A(net6237),
    .B(net2919),
    .Y(_02550_));
 sky130_fd_sc_hd__nand2_1 _18534_ (.A(net6237),
    .B(net2919),
    .Y(_02551_));
 sky130_fd_sc_hd__or2b_1 _18535_ (.A(_02550_),
    .B_N(net6238),
    .X(_02552_));
 sky130_fd_sc_hd__or2_1 _18536_ (.A(_02549_),
    .B(net6239),
    .X(_02553_));
 sky130_fd_sc_hd__a21oi_1 _18537_ (.A1(_02549_),
    .A2(net6239),
    .B1(_08246_),
    .Y(_02554_));
 sky130_fd_sc_hd__a32o_1 _18538_ (.A1(_04632_),
    .A2(_02547_),
    .A3(_02548_),
    .B1(net6240),
    .B2(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _18539_ (.A(_04623_),
    .B(_09930_),
    .Y(_02556_));
 sky130_fd_sc_hd__buf_4 _18540_ (.A(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _18541_ (.A0(net2919),
    .A1(net6241),
    .S(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_1 _18542_ (.A(net6243),
    .X(_00578_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(net4446),
    .B(_02548_),
    .Y(_02559_));
 sky130_fd_sc_hd__or2_1 _18544_ (.A(net4446),
    .B(_02548_),
    .X(_02560_));
 sky130_fd_sc_hd__o21a_1 _18545_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02551_),
    .X(_02561_));
 sky130_fd_sc_hd__nor2_1 _18546_ (.A(net4463),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02562_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(net4463),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02563_));
 sky130_fd_sc_hd__or2b_1 _18548_ (.A(_02562_),
    .B_N(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__or2_1 _18549_ (.A(_02561_),
    .B(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__a21oi_1 _18550_ (.A1(_02561_),
    .A2(_02564_),
    .B1(_08246_),
    .Y(_02566_));
 sky130_fd_sc_hd__a32o_1 _18551_ (.A1(_04632_),
    .A2(_02559_),
    .A3(_02560_),
    .B1(_02565_),
    .B2(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _18552_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_02567_),
    .S(_02557_),
    .X(_02568_));
 sky130_fd_sc_hd__clkbuf_1 _18553_ (.A(net6080),
    .X(_00579_));
 sky130_fd_sc_hd__or4_1 _18554_ (.A(net4476),
    .B(net4446),
    .C(_05403_),
    .D(net4424),
    .X(_02569_));
 sky130_fd_sc_hd__a21oi_1 _18555_ (.A1(net4476),
    .A2(_02560_),
    .B1(_04623_),
    .Y(_02570_));
 sky130_fd_sc_hd__o21ai_1 _18556_ (.A1(_02561_),
    .A2(_02562_),
    .B1(_02563_),
    .Y(_02571_));
 sky130_fd_sc_hd__buf_1 _18557_ (.A(net3241),
    .X(_02572_));
 sky130_fd_sc_hd__nor2_1 _18558_ (.A(_02572_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02573_));
 sky130_fd_sc_hd__and2_1 _18559_ (.A(net3241),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02574_));
 sky130_fd_sc_hd__or2_1 _18560_ (.A(_02573_),
    .B(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__xnor2_1 _18561_ (.A(_02571_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__a22o_1 _18562_ (.A1(_02569_),
    .A2(_02570_),
    .B1(_02576_),
    .B2(_04624_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _18563_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_02577_),
    .S(_02557_),
    .X(_02578_));
 sky130_fd_sc_hd__clkbuf_1 _18564_ (.A(net6086),
    .X(_00580_));
 sky130_fd_sc_hd__clkbuf_4 _18565_ (.A(_09935_),
    .X(_02579_));
 sky130_fd_sc_hd__o21a_1 _18566_ (.A1(net3241),
    .A2(\rbzero.wall_tracer.rayAddendX[-2] ),
    .B1(_02571_),
    .X(_02580_));
 sky130_fd_sc_hd__nand2_1 _18567_ (.A(_05401_),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02581_));
 sky130_fd_sc_hd__or2_1 _18568_ (.A(net4690),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02582_));
 sky130_fd_sc_hd__o211a_1 _18569_ (.A1(_02574_),
    .A2(_02580_),
    .B1(net7585),
    .C1(net4691),
    .X(_02583_));
 sky130_fd_sc_hd__inv_2 _18570_ (.A(net7586),
    .Y(_02584_));
 sky130_fd_sc_hd__a211o_1 _18571_ (.A1(net4691),
    .A2(_02581_),
    .B1(_02580_),
    .C1(_02574_),
    .X(_02585_));
 sky130_fd_sc_hd__o31a_1 _18572_ (.A1(net4476),
    .A2(net4446),
    .A3(_05403_),
    .B1(_02545_),
    .X(_02586_));
 sky130_fd_sc_hd__or2_1 _18573_ (.A(net3838),
    .B(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__nand2_1 _18574_ (.A(net3838),
    .B(_02586_),
    .Y(_02588_));
 sky130_fd_sc_hd__a32o_1 _18575_ (.A1(_04633_),
    .A2(_02587_),
    .A3(_02588_),
    .B1(_09933_),
    .B2(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02589_));
 sky130_fd_sc_hd__a31o_1 _18576_ (.A1(_02579_),
    .A2(_02584_),
    .A3(net4692),
    .B1(net3406),
    .X(_00581_));
 sky130_fd_sc_hd__xor2_1 _18577_ (.A(net6237),
    .B(_05403_),
    .X(_02590_));
 sky130_fd_sc_hd__nand2_1 _18578_ (.A(net3838),
    .B(net4424),
    .Y(_02591_));
 sky130_fd_sc_hd__o21ai_1 _18579_ (.A1(net3838),
    .A2(_02569_),
    .B1(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__xnor2_1 _18580_ (.A(_02590_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__nand2_1 _18581_ (.A(net7585),
    .B(_02584_),
    .Y(_02594_));
 sky130_fd_sc_hd__or2_1 _18582_ (.A(net4587),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02595_));
 sky130_fd_sc_hd__nand2_1 _18583_ (.A(net4587),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02596_));
 sky130_fd_sc_hd__nand2_1 _18584_ (.A(_02595_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__xnor2_1 _18585_ (.A(_02594_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__mux2_1 _18586_ (.A0(_02593_),
    .A1(_02598_),
    .S(_04623_),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _18587_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_02599_),
    .S(_02557_),
    .X(_02600_));
 sky130_fd_sc_hd__clkbuf_1 _18588_ (.A(net6117),
    .X(_00582_));
 sky130_fd_sc_hd__nand2_1 _18589_ (.A(net4666),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02601_));
 sky130_fd_sc_hd__or2_1 _18590_ (.A(net4666),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02602_));
 sky130_fd_sc_hd__a21bo_1 _18591_ (.A1(_02594_),
    .A2(_02595_),
    .B1_N(_02596_),
    .X(_02603_));
 sky130_fd_sc_hd__a21o_1 _18592_ (.A1(net4667),
    .A2(_02602_),
    .B1(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__and3_1 _18593_ (.A(net4667),
    .B(net7601),
    .C(_02603_),
    .X(_02605_));
 sky130_fd_sc_hd__inv_2 _18594_ (.A(net7602),
    .Y(_02606_));
 sky130_fd_sc_hd__nor2_1 _18595_ (.A(net4463),
    .B(net4446),
    .Y(_02607_));
 sky130_fd_sc_hd__and2_1 _18596_ (.A(net4463),
    .B(net4446),
    .X(_02608_));
 sky130_fd_sc_hd__nor4_1 _18597_ (.A(net6237),
    .B(_05403_),
    .C(_02607_),
    .D(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__o22a_1 _18598_ (.A1(net6237),
    .A2(_05403_),
    .B1(_02607_),
    .B2(_02608_),
    .X(_02610_));
 sky130_fd_sc_hd__or2_1 _18599_ (.A(_02609_),
    .B(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__o2bb2a_1 _18600_ (.A1_N(_02590_),
    .A2_N(_02591_),
    .B1(net3838),
    .B2(_02569_),
    .X(_02612_));
 sky130_fd_sc_hd__nor2_1 _18601_ (.A(_02611_),
    .B(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21o_1 _18602_ (.A1(_02611_),
    .A2(_02612_),
    .B1(_04624_),
    .X(_02614_));
 sky130_fd_sc_hd__a2bb2o_1 _18603_ (.A1_N(_02613_),
    .A2_N(_02614_),
    .B1(\rbzero.wall_tracer.rayAddendX[1] ),
    .B2(_09932_),
    .X(_02615_));
 sky130_fd_sc_hd__a31o_1 _18604_ (.A1(_02579_),
    .A2(net4668),
    .A3(_02606_),
    .B1(net3603),
    .X(_00583_));
 sky130_fd_sc_hd__xor2_1 _18605_ (.A(net4666),
    .B(net3796),
    .X(_02616_));
 sky130_fd_sc_hd__and2_1 _18606_ (.A(net4667),
    .B(_02606_),
    .X(_02617_));
 sky130_fd_sc_hd__xnor2_1 _18607_ (.A(_02616_),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__xor2_1 _18608_ (.A(net3242),
    .B(net4493),
    .X(_02619_));
 sky130_fd_sc_hd__or3_1 _18609_ (.A(net87),
    .B(_02613_),
    .C(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__o21ai_1 _18610_ (.A1(net87),
    .A2(_02613_),
    .B1(_02619_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand2_1 _18611_ (.A(_02620_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xnor2_1 _18612_ (.A(_02607_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__mux2_1 _18613_ (.A0(_02618_),
    .A1(_02623_),
    .S(_04632_),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _18614_ (.A0(net3796),
    .A1(_02624_),
    .S(_02557_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _18615_ (.A(net3797),
    .X(_00584_));
 sky130_fd_sc_hd__inv_2 _18616_ (.A(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02626_));
 sky130_fd_sc_hd__or2_1 _18617_ (.A(_05401_),
    .B(net3838),
    .X(_02627_));
 sky130_fd_sc_hd__nand2_1 _18618_ (.A(_05401_),
    .B(net3838),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__or3_1 _18620_ (.A(net3242),
    .B(net4476),
    .C(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__o21ai_1 _18621_ (.A1(net3242),
    .A2(net4493),
    .B1(_02629_),
    .Y(_02631_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(_02630_),
    .B(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__o21ai_1 _18623_ (.A1(_02613_),
    .A2(_02619_),
    .B1(_02607_),
    .Y(_02633_));
 sky130_fd_sc_hd__a21o_1 _18624_ (.A1(_02621_),
    .A2(_02633_),
    .B1(_02632_),
    .X(_02634_));
 sky130_fd_sc_hd__nand2_1 _18625_ (.A(_04633_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__a31o_1 _18626_ (.A1(_02621_),
    .A2(_02632_),
    .A3(_02633_),
    .B1(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_4 _18627_ (.A(net4666),
    .X(_02637_));
 sky130_fd_sc_hd__nand2_1 _18628_ (.A(_02637_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02638_));
 sky130_fd_sc_hd__or2_1 _18629_ (.A(_02637_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02639_));
 sky130_fd_sc_hd__o21a_1 _18630_ (.A1(net3796),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(net4666),
    .X(_02640_));
 sky130_fd_sc_hd__a21o_1 _18631_ (.A1(_02605_),
    .A2(_02616_),
    .B1(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__a21oi_1 _18632_ (.A1(net4752),
    .A2(_02639_),
    .B1(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__and3_1 _18633_ (.A(net4752),
    .B(_02639_),
    .C(_02641_),
    .X(_02643_));
 sky130_fd_sc_hd__or3_1 _18634_ (.A(_09943_),
    .B(net4753),
    .C(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__o211ai_1 _18635_ (.A1(net1999),
    .A2(_02557_),
    .B1(_02636_),
    .C1(net4754),
    .Y(_00585_));
 sky130_fd_sc_hd__xor2_1 _18636_ (.A(_02637_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02645_));
 sky130_fd_sc_hd__buf_2 _18637_ (.A(_02637_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_4 _18638_ (.A(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__a21oi_1 _18639_ (.A1(_02647_),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02643_),
    .Y(_02648_));
 sky130_fd_sc_hd__xnor2_1 _18640_ (.A(_02645_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__nor2_1 _18641_ (.A(net4587),
    .B(net6237),
    .Y(_02650_));
 sky130_fd_sc_hd__and2_1 _18642_ (.A(net4587),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_02651_));
 sky130_fd_sc_hd__or2_1 _18643_ (.A(_02650_),
    .B(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__nand3_1 _18644_ (.A(_02630_),
    .B(_02634_),
    .C(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__a21o_1 _18645_ (.A1(_02630_),
    .A2(_02634_),
    .B1(_02652_),
    .X(_02654_));
 sky130_fd_sc_hd__a21oi_1 _18646_ (.A1(_02653_),
    .A2(_02654_),
    .B1(_02627_),
    .Y(_02655_));
 sky130_fd_sc_hd__and3_1 _18647_ (.A(_02627_),
    .B(_02653_),
    .C(_02654_),
    .X(_02656_));
 sky130_fd_sc_hd__or2_1 _18648_ (.A(_02655_),
    .B(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _18649_ (.A0(_02649_),
    .A1(_02657_),
    .S(_04632_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _18650_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02658_),
    .S(_02557_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_1 _18651_ (.A(net6095),
    .X(_00586_));
 sky130_fd_sc_hd__nand2_1 _18652_ (.A(_02637_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02660_));
 sky130_fd_sc_hd__or2_1 _18653_ (.A(_02637_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02661_));
 sky130_fd_sc_hd__and2_1 _18654_ (.A(net4696),
    .B(net7608),
    .X(_02662_));
 sky130_fd_sc_hd__and2_1 _18655_ (.A(_02643_),
    .B(_02645_),
    .X(_02663_));
 sky130_fd_sc_hd__o21a_1 _18656_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02637_),
    .X(_02664_));
 sky130_fd_sc_hd__or3_1 _18657_ (.A(_02662_),
    .B(_02663_),
    .C(net4767),
    .X(_02665_));
 sky130_fd_sc_hd__o21ai_1 _18658_ (.A1(_02663_),
    .A2(net4767),
    .B1(_02662_),
    .Y(_02666_));
 sky130_fd_sc_hd__a21o_1 _18659_ (.A1(_02634_),
    .A2(_02652_),
    .B1(_02627_),
    .X(_02667_));
 sky130_fd_sc_hd__xor2_1 _18660_ (.A(_02637_),
    .B(net4463),
    .X(_02668_));
 sky130_fd_sc_hd__xnor2_1 _18661_ (.A(_02650_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a21oi_1 _18662_ (.A1(_02654_),
    .A2(_02667_),
    .B1(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__a31o_1 _18663_ (.A1(_02654_),
    .A2(_02669_),
    .A3(_02667_),
    .B1(_04623_),
    .X(_02671_));
 sky130_fd_sc_hd__a2bb2o_1 _18664_ (.A1_N(_02670_),
    .A2_N(_02671_),
    .B1(\rbzero.wall_tracer.rayAddendX[5] ),
    .B2(_09932_),
    .X(_02672_));
 sky130_fd_sc_hd__a31o_1 _18665_ (.A1(_02579_),
    .A2(net4768),
    .A3(net7609),
    .B1(net3552),
    .X(_00587_));
 sky130_fd_sc_hd__xnor2_2 _18666_ (.A(_02637_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02673_));
 sky130_fd_sc_hd__a21o_1 _18667_ (.A1(net4696),
    .A2(_02666_),
    .B1(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__nand3_1 _18668_ (.A(net4696),
    .B(_02666_),
    .C(net7571),
    .Y(_02675_));
 sky130_fd_sc_hd__inv_2 _18669_ (.A(_02646_),
    .Y(_02676_));
 sky130_fd_sc_hd__inv_2 _18670_ (.A(net4463),
    .Y(_02677_));
 sky130_fd_sc_hd__or2_1 _18671_ (.A(_02646_),
    .B(net3242),
    .X(_02678_));
 sky130_fd_sc_hd__nand2_1 _18672_ (.A(_02646_),
    .B(net3242),
    .Y(_02679_));
 sky130_fd_sc_hd__a22o_1 _18673_ (.A1(_02676_),
    .A2(_02677_),
    .B1(_02678_),
    .B2(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__or3b_1 _18674_ (.A(_02646_),
    .B(net4463),
    .C_N(net3242),
    .X(_02681_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(_02680_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__a21o_1 _18676_ (.A1(_02650_),
    .A2(_02668_),
    .B1(_02670_),
    .X(_02683_));
 sky130_fd_sc_hd__xnor2_1 _18677_ (.A(_02682_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__a22o_1 _18678_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_09933_),
    .B1(_02684_),
    .B2(_04633_),
    .X(_02685_));
 sky130_fd_sc_hd__a31o_1 _18679_ (.A1(_02579_),
    .A2(net4697),
    .A3(net7572),
    .B1(net3689),
    .X(_00588_));
 sky130_fd_sc_hd__nand2_2 _18680_ (.A(_02646_),
    .B(net3043),
    .Y(_02686_));
 sky130_fd_sc_hd__or2_1 _18681_ (.A(_02646_),
    .B(net3043),
    .X(_02687_));
 sky130_fd_sc_hd__inv_2 _18682_ (.A(_02673_),
    .Y(_02688_));
 sky130_fd_sc_hd__o21a_1 _18683_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .B1(_02637_),
    .X(_02689_));
 sky130_fd_sc_hd__a311o_1 _18684_ (.A1(_02662_),
    .A2(_02663_),
    .A3(_02688_),
    .B1(net4810),
    .C1(net4767),
    .X(_02690_));
 sky130_fd_sc_hd__a21o_1 _18685_ (.A1(_02686_),
    .A2(_02687_),
    .B1(net4811),
    .X(_02691_));
 sky130_fd_sc_hd__nand3_2 _18686_ (.A(_02686_),
    .B(_02687_),
    .C(net4811),
    .Y(_02692_));
 sky130_fd_sc_hd__or2_1 _18687_ (.A(_02646_),
    .B(_05401_),
    .X(_02693_));
 sky130_fd_sc_hd__nand2_1 _18688_ (.A(_02647_),
    .B(_05401_),
    .Y(_02694_));
 sky130_fd_sc_hd__a21bo_1 _18689_ (.A1(_02693_),
    .A2(_02694_),
    .B1_N(_02678_),
    .X(_02695_));
 sky130_fd_sc_hd__or3b_4 _18690_ (.A(_02647_),
    .B(net3242),
    .C_N(_05401_),
    .X(_02696_));
 sky130_fd_sc_hd__and3_1 _18691_ (.A(_02676_),
    .B(net3242),
    .C(_02677_),
    .X(_02697_));
 sky130_fd_sc_hd__and3_1 _18692_ (.A(_02680_),
    .B(_02681_),
    .C(_02683_),
    .X(_02698_));
 sky130_fd_sc_hd__a211o_1 _18693_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02697_),
    .C1(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__o211ai_4 _18694_ (.A1(_02697_),
    .A2(_02698_),
    .B1(_02695_),
    .C1(_02696_),
    .Y(_02700_));
 sky130_fd_sc_hd__a32o_1 _18695_ (.A1(_04633_),
    .A2(_02699_),
    .A3(_02700_),
    .B1(_09933_),
    .B2(net3043),
    .X(_02701_));
 sky130_fd_sc_hd__a31o_1 _18696_ (.A1(_02579_),
    .A2(net4812),
    .A3(_02692_),
    .B1(net3044),
    .X(_00589_));
 sky130_fd_sc_hd__nand2_1 _18697_ (.A(_02646_),
    .B(net7146),
    .Y(_02702_));
 sky130_fd_sc_hd__or2_1 _18698_ (.A(_02646_),
    .B(net7146),
    .X(_02703_));
 sky130_fd_sc_hd__nand2_1 _18699_ (.A(_02702_),
    .B(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__a21oi_1 _18700_ (.A1(_02686_),
    .A2(_02692_),
    .B1(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__a31o_1 _18701_ (.A1(_02686_),
    .A2(_02692_),
    .A3(_02704_),
    .B1(_08246_),
    .X(_02706_));
 sky130_fd_sc_hd__or2_1 _18702_ (.A(_02647_),
    .B(net4587),
    .X(_02707_));
 sky130_fd_sc_hd__nand2_1 _18703_ (.A(_02647_),
    .B(net4587),
    .Y(_02708_));
 sky130_fd_sc_hd__nand2_1 _18704_ (.A(_02707_),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__xnor2_1 _18705_ (.A(_02693_),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__a21oi_1 _18706_ (.A1(_02696_),
    .A2(_02700_),
    .B1(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a31o_1 _18707_ (.A1(_02696_),
    .A2(_02700_),
    .A3(_02710_),
    .B1(_04623_),
    .X(_02712_));
 sky130_fd_sc_hd__o22ai_1 _18708_ (.A1(_02705_),
    .A2(_02706_),
    .B1(_02711_),
    .B2(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__buf_4 _18709_ (.A(_02556_),
    .X(_02714_));
 sky130_fd_sc_hd__mux2_1 _18710_ (.A0(net7146),
    .A1(_02713_),
    .S(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_1 _18711_ (.A(net3195),
    .X(_00590_));
 sky130_fd_sc_hd__or2_1 _18712_ (.A(_02647_),
    .B(net4787),
    .X(_02716_));
 sky130_fd_sc_hd__nand2_1 _18713_ (.A(_02647_),
    .B(net4787),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2_1 _18714_ (.A(_02716_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__o211a_1 _18715_ (.A1(_02692_),
    .A2(_02704_),
    .B1(_02702_),
    .C1(_02686_),
    .X(_02719_));
 sky130_fd_sc_hd__xor2_1 _18716_ (.A(_02718_),
    .B(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__a211oi_1 _18717_ (.A1(net4587),
    .A2(_05401_),
    .B1(_02711_),
    .C1(_02647_),
    .Y(_02721_));
 sky130_fd_sc_hd__a211o_1 _18718_ (.A1(_02707_),
    .A2(_02711_),
    .B1(_02721_),
    .C1(_04624_),
    .X(_02722_));
 sky130_fd_sc_hd__o221a_1 _18719_ (.A1(net4787),
    .A2(_02557_),
    .B1(_09943_),
    .B2(_02720_),
    .C1(_02722_),
    .X(_00591_));
 sky130_fd_sc_hd__o21a_1 _18720_ (.A1(_02718_),
    .A2(_02719_),
    .B1(_02717_),
    .X(_02723_));
 sky130_fd_sc_hd__xor2_1 _18721_ (.A(_02647_),
    .B(net6304),
    .X(_02724_));
 sky130_fd_sc_hd__xnor2_1 _18722_ (.A(_02723_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__o311a_1 _18723_ (.A1(net4587),
    .A2(_05401_),
    .A3(_02700_),
    .B1(_08246_),
    .C1(_02676_),
    .X(_02726_));
 sky130_fd_sc_hd__a21o_1 _18724_ (.A1(_04624_),
    .A2(_02725_),
    .B1(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__mux2_1 _18725_ (.A0(net6304),
    .A1(_02727_),
    .S(_02714_),
    .X(_02728_));
 sky130_fd_sc_hd__clkbuf_1 _18726_ (.A(net3198),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _18727_ (.A0(net3917),
    .A1(_06227_),
    .S(_02261_),
    .X(_02729_));
 sky130_fd_sc_hd__mux2_1 _18728_ (.A0(net3918),
    .A1(_06185_),
    .S(_06394_),
    .X(_02730_));
 sky130_fd_sc_hd__clkbuf_1 _18729_ (.A(net3919),
    .X(_00593_));
 sky130_fd_sc_hd__nor2_1 _18730_ (.A(_06185_),
    .B(_06188_),
    .Y(_02731_));
 sky130_fd_sc_hd__or3_1 _18731_ (.A(_06205_),
    .B(_06189_),
    .C(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__o21ai_1 _18732_ (.A1(net3881),
    .A2(_09987_),
    .B1(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__mux2_1 _18733_ (.A0(net3882),
    .A1(_06186_),
    .S(_06394_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_1 _18734_ (.A(net3883),
    .X(_00594_));
 sky130_fd_sc_hd__or3_1 _18735_ (.A(net6186),
    .B(_06189_),
    .C(_06191_),
    .X(_02735_));
 sky130_fd_sc_hd__nor2_1 _18736_ (.A(_01870_),
    .B(_06192_),
    .Y(_02736_));
 sky130_fd_sc_hd__a22o_1 _18737_ (.A1(net4387),
    .A2(_10019_),
    .B1(net6187),
    .B2(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__mux2_1 _18738_ (.A0(net6188),
    .A1(net3804),
    .S(_06394_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_1 _18739_ (.A(net3805),
    .X(_00595_));
 sky130_fd_sc_hd__xnor2_1 _18740_ (.A(_06183_),
    .B(_06396_),
    .Y(_02739_));
 sky130_fd_sc_hd__xnor2_1 _18741_ (.A(_06193_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__mux2_1 _18742_ (.A0(net3893),
    .A1(_02740_),
    .S(_02261_),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _18743_ (.A0(net3894),
    .A1(_06183_),
    .S(_06394_),
    .X(_02742_));
 sky130_fd_sc_hd__clkbuf_1 _18744_ (.A(net3895),
    .X(_00596_));
 sky130_fd_sc_hd__xnor2_1 _18745_ (.A(_06197_),
    .B(_06195_),
    .Y(_02743_));
 sky130_fd_sc_hd__mux2_1 _18746_ (.A0(net3279),
    .A1(_02743_),
    .S(_02261_),
    .X(_02744_));
 sky130_fd_sc_hd__mux2_1 _18747_ (.A0(net3280),
    .A1(net4821),
    .S(_06394_),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_1 _18748_ (.A(net3281),
    .X(_00597_));
 sky130_fd_sc_hd__a21oi_1 _18749_ (.A1(net4821),
    .A2(_06396_),
    .B1(_06198_),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_1 _18750_ (.A(_06182_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__mux2_1 _18751_ (.A0(net3952),
    .A1(_02747_),
    .S(_09999_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _18752_ (.A0(_02748_),
    .A1(net6309),
    .S(_06392_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_1 _18753_ (.A(net3035),
    .X(_00598_));
 sky130_fd_sc_hd__nor2_1 _18754_ (.A(net4799),
    .B(net941),
    .Y(_02750_));
 sky130_fd_sc_hd__nor2_1 _18755_ (.A(net4640),
    .B(net4905),
    .Y(_02751_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_05393_),
    .B(net738),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_1 _18757_ (.A(net4438),
    .B(net723),
    .Y(_02753_));
 sky130_fd_sc_hd__or2_1 _18758_ (.A(net4620),
    .B(net738),
    .X(_02754_));
 sky130_fd_sc_hd__nand3b_1 _18759_ (.A_N(net4439),
    .B(net4621),
    .C(_02752_),
    .Y(_02755_));
 sky130_fd_sc_hd__and2_1 _18760_ (.A(_02752_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__nand2_1 _18761_ (.A(net4640),
    .B(net4905),
    .Y(_02757_));
 sky130_fd_sc_hd__o21a_1 _18762_ (.A1(_02751_),
    .A2(_02756_),
    .B1(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__nand2_1 _18763_ (.A(net4799),
    .B(net941),
    .Y(_02759_));
 sky130_fd_sc_hd__o21a_1 _18764_ (.A1(_02750_),
    .A2(_02758_),
    .B1(net4800),
    .X(_02760_));
 sky130_fd_sc_hd__nor2_1 _18765_ (.A(net4549),
    .B(net1091),
    .Y(_02761_));
 sky130_fd_sc_hd__nand2_1 _18766_ (.A(_05396_),
    .B(net1091),
    .Y(_02762_));
 sky130_fd_sc_hd__or2b_1 _18767_ (.A(net4550),
    .B_N(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__xor2_1 _18768_ (.A(_02760_),
    .B(net4551),
    .X(_02764_));
 sky130_fd_sc_hd__inv_2 _18769_ (.A(net4438),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_1 _18770_ (.A(_02765_),
    .B(_08195_),
    .Y(_02766_));
 sky130_fd_sc_hd__a221o_1 _18771_ (.A1(net1091),
    .A2(_02528_),
    .B1(_02529_),
    .B2(net4552),
    .C1(_02766_),
    .X(_00599_));
 sky130_fd_sc_hd__nand2_1 _18772_ (.A(_05393_),
    .B(net4438),
    .Y(_02767_));
 sky130_fd_sc_hd__or2_1 _18773_ (.A(_05393_),
    .B(net4438),
    .X(_02768_));
 sky130_fd_sc_hd__o21a_1 _18774_ (.A1(_02760_),
    .A2(net4550),
    .B1(_02762_),
    .X(_02769_));
 sky130_fd_sc_hd__nor2_1 _18775_ (.A(net3807),
    .B(net2884),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _18776_ (.A(net3807),
    .B(net2884),
    .Y(_02771_));
 sky130_fd_sc_hd__or2b_1 _18777_ (.A(_02770_),
    .B_N(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__or2_1 _18778_ (.A(_02769_),
    .B(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__a21oi_1 _18779_ (.A1(_02769_),
    .A2(_02772_),
    .B1(_08246_),
    .Y(_02774_));
 sky130_fd_sc_hd__a32o_1 _18780_ (.A1(_04632_),
    .A2(_02767_),
    .A3(_02768_),
    .B1(_02773_),
    .B2(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _18781_ (.A0(net6222),
    .A1(_02775_),
    .S(_02714_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _18782_ (.A(net2885),
    .X(_00600_));
 sky130_fd_sc_hd__nand2_1 _18783_ (.A(net4640),
    .B(_02768_),
    .Y(_02777_));
 sky130_fd_sc_hd__or2_1 _18784_ (.A(net4640),
    .B(_02768_),
    .X(_02778_));
 sky130_fd_sc_hd__o21a_1 _18785_ (.A1(_02769_),
    .A2(_02770_),
    .B1(_02771_),
    .X(_02779_));
 sky130_fd_sc_hd__nor2_1 _18786_ (.A(net4459),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_1 _18787_ (.A(net4459),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02781_));
 sky130_fd_sc_hd__or2b_1 _18788_ (.A(_02780_),
    .B_N(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__or2_1 _18789_ (.A(_02779_),
    .B(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__a21oi_1 _18790_ (.A1(_02779_),
    .A2(_02782_),
    .B1(_08246_),
    .Y(_02784_));
 sky130_fd_sc_hd__a32o_1 _18791_ (.A1(_04632_),
    .A2(_02777_),
    .A3(_02778_),
    .B1(_02783_),
    .B2(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _18792_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(_02785_),
    .S(_02714_),
    .X(_02786_));
 sky130_fd_sc_hd__clkbuf_1 _18793_ (.A(net6089),
    .X(_00601_));
 sky130_fd_sc_hd__or4_1 _18794_ (.A(net4799),
    .B(net4640),
    .C(_05393_),
    .D(net4438),
    .X(_02787_));
 sky130_fd_sc_hd__a21oi_1 _18795_ (.A1(net4799),
    .A2(_02778_),
    .B1(_04623_),
    .Y(_02788_));
 sky130_fd_sc_hd__o21ai_1 _18796_ (.A1(_02779_),
    .A2(_02780_),
    .B1(_02781_),
    .Y(_02789_));
 sky130_fd_sc_hd__clkbuf_1 _18797_ (.A(net3699),
    .X(_02790_));
 sky130_fd_sc_hd__nor2_1 _18798_ (.A(net3700),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_02791_));
 sky130_fd_sc_hd__and2_1 _18799_ (.A(net3699),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02792_));
 sky130_fd_sc_hd__or2_1 _18800_ (.A(_02791_),
    .B(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__xnor2_1 _18801_ (.A(_02789_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__a22o_1 _18802_ (.A1(_02787_),
    .A2(_02788_),
    .B1(_02794_),
    .B2(_04624_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _18803_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(_02795_),
    .S(_02714_),
    .X(_02796_));
 sky130_fd_sc_hd__clkbuf_1 _18804_ (.A(net6109),
    .X(_00602_));
 sky130_fd_sc_hd__o21a_1 _18805_ (.A1(net3699),
    .A2(\rbzero.wall_tracer.rayAddendY[-2] ),
    .B1(_02789_),
    .X(_02797_));
 sky130_fd_sc_hd__nand2_1 _18806_ (.A(_05391_),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_02798_));
 sky130_fd_sc_hd__or2_1 _18807_ (.A(net4625),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02799_));
 sky130_fd_sc_hd__o211a_1 _18808_ (.A1(_02792_),
    .A2(_02797_),
    .B1(net7575),
    .C1(net4626),
    .X(_02800_));
 sky130_fd_sc_hd__inv_2 _18809_ (.A(net7576),
    .Y(_02801_));
 sky130_fd_sc_hd__a211o_1 _18810_ (.A1(net4626),
    .A2(_02798_),
    .B1(_02797_),
    .C1(_02792_),
    .X(_02802_));
 sky130_fd_sc_hd__o31a_1 _18811_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .A3(_05393_),
    .B1(_02765_),
    .X(_02803_));
 sky130_fd_sc_hd__or2_1 _18812_ (.A(_05396_),
    .B(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__nand2_1 _18813_ (.A(_05396_),
    .B(_02803_),
    .Y(_02805_));
 sky130_fd_sc_hd__a32o_1 _18814_ (.A1(_04633_),
    .A2(_02804_),
    .A3(_02805_),
    .B1(_09933_),
    .B2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02806_));
 sky130_fd_sc_hd__a31o_1 _18815_ (.A1(_02579_),
    .A2(_02801_),
    .A3(net4627),
    .B1(net3133),
    .X(_00603_));
 sky130_fd_sc_hd__xor2_1 _18816_ (.A(net3807),
    .B(_05393_),
    .X(_02807_));
 sky130_fd_sc_hd__nand2_1 _18817_ (.A(_05396_),
    .B(net4438),
    .Y(_02808_));
 sky130_fd_sc_hd__o21ai_1 _18818_ (.A1(_05396_),
    .A2(_02787_),
    .B1(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__xnor2_1 _18819_ (.A(_02807_),
    .B(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__nand2_1 _18820_ (.A(net7575),
    .B(_02801_),
    .Y(_02811_));
 sky130_fd_sc_hd__or2_1 _18821_ (.A(net4634),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02812_));
 sky130_fd_sc_hd__nand2_1 _18822_ (.A(net4634),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_1 _18823_ (.A(_02812_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__xnor2_1 _18824_ (.A(_02811_),
    .B(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__mux2_1 _18825_ (.A0(_02810_),
    .A1(_02815_),
    .S(_04623_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _18826_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_02816_),
    .S(_02714_),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _18827_ (.A(net6120),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _18828_ (.A(net4708),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_02818_));
 sky130_fd_sc_hd__or2_1 _18829_ (.A(net4708),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02819_));
 sky130_fd_sc_hd__a21bo_1 _18830_ (.A1(_02811_),
    .A2(_02812_),
    .B1_N(_02813_),
    .X(_02820_));
 sky130_fd_sc_hd__a21o_1 _18831_ (.A1(net4709),
    .A2(_02819_),
    .B1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__and3_1 _18832_ (.A(net4709),
    .B(net7611),
    .C(_02820_),
    .X(_02822_));
 sky130_fd_sc_hd__inv_2 _18833_ (.A(net7612),
    .Y(_02823_));
 sky130_fd_sc_hd__nor2_1 _18834_ (.A(net4459),
    .B(net4640),
    .Y(_02824_));
 sky130_fd_sc_hd__and2_1 _18835_ (.A(net4459),
    .B(net4640),
    .X(_02825_));
 sky130_fd_sc_hd__nor4_1 _18836_ (.A(net3807),
    .B(_05393_),
    .C(_02824_),
    .D(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__o22a_1 _18837_ (.A1(net3807),
    .A2(_05393_),
    .B1(_02824_),
    .B2(_02825_),
    .X(_02827_));
 sky130_fd_sc_hd__or2_1 _18838_ (.A(net1580),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__o2bb2a_1 _18839_ (.A1_N(_02807_),
    .A2_N(_02808_),
    .B1(_05396_),
    .B2(_02787_),
    .X(_02829_));
 sky130_fd_sc_hd__nor2_1 _18840_ (.A(_02828_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__a21o_1 _18841_ (.A1(_02828_),
    .A2(_02829_),
    .B1(_04624_),
    .X(_02831_));
 sky130_fd_sc_hd__a2bb2o_1 _18842_ (.A1_N(_02830_),
    .A2_N(_02831_),
    .B1(\rbzero.wall_tracer.rayAddendY[1] ),
    .B2(_09932_),
    .X(_02832_));
 sky130_fd_sc_hd__a31o_1 _18843_ (.A1(_02529_),
    .A2(net4710),
    .A3(_02823_),
    .B1(net3862),
    .X(_00605_));
 sky130_fd_sc_hd__xor2_1 _18844_ (.A(net4708),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_02833_));
 sky130_fd_sc_hd__and2_1 _18845_ (.A(net4709),
    .B(_02823_),
    .X(_02834_));
 sky130_fd_sc_hd__xnor2_1 _18846_ (.A(_02833_),
    .B(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__xor2_1 _18847_ (.A(net3700),
    .B(net4799),
    .X(_02836_));
 sky130_fd_sc_hd__or3_1 _18848_ (.A(net1580),
    .B(_02830_),
    .C(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__o21ai_1 _18849_ (.A1(net1580),
    .A2(_02830_),
    .B1(_02836_),
    .Y(_02838_));
 sky130_fd_sc_hd__nand2_1 _18850_ (.A(_02837_),
    .B(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__xnor2_1 _18851_ (.A(_02824_),
    .B(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__mux2_1 _18852_ (.A0(_02835_),
    .A1(_02840_),
    .S(_04632_),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _18853_ (.A0(\rbzero.wall_tracer.rayAddendY[2] ),
    .A1(_02841_),
    .S(_02714_),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _18854_ (.A(net6069),
    .X(_00606_));
 sky130_fd_sc_hd__inv_2 _18855_ (.A(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02843_));
 sky130_fd_sc_hd__or2_1 _18856_ (.A(_05391_),
    .B(_05396_),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_1 _18857_ (.A(_05391_),
    .B(_05396_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _18858_ (.A(_02844_),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__or3_1 _18859_ (.A(net3700),
    .B(net4799),
    .C(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__o21ai_1 _18860_ (.A1(net3700),
    .A2(net4799),
    .B1(_02846_),
    .Y(_02848_));
 sky130_fd_sc_hd__nand2_1 _18861_ (.A(_02847_),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__o21ai_1 _18862_ (.A1(_02830_),
    .A2(_02836_),
    .B1(_02824_),
    .Y(_02850_));
 sky130_fd_sc_hd__a21o_1 _18863_ (.A1(_02838_),
    .A2(_02850_),
    .B1(_02849_),
    .X(_02851_));
 sky130_fd_sc_hd__nand2_1 _18864_ (.A(_04633_),
    .B(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__a31o_1 _18865_ (.A1(_02838_),
    .A2(_02849_),
    .A3(_02850_),
    .B1(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_4 _18866_ (.A(net4708),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _18867_ (.A(_02854_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02855_));
 sky130_fd_sc_hd__or2_1 _18868_ (.A(_02854_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02856_));
 sky130_fd_sc_hd__o21a_1 _18869_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(net4708),
    .X(_02857_));
 sky130_fd_sc_hd__a21o_1 _18870_ (.A1(_02822_),
    .A2(_02833_),
    .B1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__a21oi_1 _18871_ (.A1(net4721),
    .A2(_02856_),
    .B1(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__and3_1 _18872_ (.A(net4721),
    .B(_02856_),
    .C(_02858_),
    .X(_02860_));
 sky130_fd_sc_hd__or3_1 _18873_ (.A(_09943_),
    .B(net4722),
    .C(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__o211ai_1 _18874_ (.A1(net1581),
    .A2(_02557_),
    .B1(_02853_),
    .C1(net4723),
    .Y(_00607_));
 sky130_fd_sc_hd__xor2_1 _18875_ (.A(_02854_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_02862_));
 sky130_fd_sc_hd__buf_2 _18876_ (.A(_02854_),
    .X(_02863_));
 sky130_fd_sc_hd__buf_2 _18877_ (.A(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__a21oi_1 _18878_ (.A1(_02864_),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02860_),
    .Y(_02865_));
 sky130_fd_sc_hd__xnor2_1 _18879_ (.A(_02862_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__nor2_1 _18880_ (.A(net4634),
    .B(net3807),
    .Y(_02867_));
 sky130_fd_sc_hd__and2_1 _18881_ (.A(net4634),
    .B(net3807),
    .X(_02868_));
 sky130_fd_sc_hd__or2_1 _18882_ (.A(_02867_),
    .B(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__nand3_1 _18883_ (.A(_02847_),
    .B(_02851_),
    .C(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__a21o_1 _18884_ (.A1(_02847_),
    .A2(_02851_),
    .B1(_02869_),
    .X(_02871_));
 sky130_fd_sc_hd__a21oi_1 _18885_ (.A1(_02870_),
    .A2(_02871_),
    .B1(_02844_),
    .Y(_02872_));
 sky130_fd_sc_hd__and3_1 _18886_ (.A(_02844_),
    .B(_02870_),
    .C(_02871_),
    .X(_02873_));
 sky130_fd_sc_hd__or2_1 _18887_ (.A(_02872_),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _18888_ (.A0(_02866_),
    .A1(_02874_),
    .S(_04632_),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _18889_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_02875_),
    .S(_02714_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_1 _18890_ (.A(net6102),
    .X(_00608_));
 sky130_fd_sc_hd__nand2_1 _18891_ (.A(_02854_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_02877_));
 sky130_fd_sc_hd__or2_1 _18892_ (.A(_02854_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_02878_));
 sky130_fd_sc_hd__and2_1 _18893_ (.A(net4662),
    .B(net7598),
    .X(_02879_));
 sky130_fd_sc_hd__and2_1 _18894_ (.A(_02860_),
    .B(_02862_),
    .X(_02880_));
 sky130_fd_sc_hd__o21a_1 _18895_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02854_),
    .X(_02881_));
 sky130_fd_sc_hd__or3_1 _18896_ (.A(_02879_),
    .B(_02880_),
    .C(net4758),
    .X(_02882_));
 sky130_fd_sc_hd__o21ai_1 _18897_ (.A1(_02880_),
    .A2(net4758),
    .B1(_02879_),
    .Y(_02883_));
 sky130_fd_sc_hd__a21o_1 _18898_ (.A1(_02851_),
    .A2(_02869_),
    .B1(_02844_),
    .X(_02884_));
 sky130_fd_sc_hd__xor2_1 _18899_ (.A(_02854_),
    .B(net4459),
    .X(_02885_));
 sky130_fd_sc_hd__xnor2_1 _18900_ (.A(_02867_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__a21oi_1 _18901_ (.A1(_02871_),
    .A2(_02884_),
    .B1(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__a31o_1 _18902_ (.A1(_02871_),
    .A2(_02886_),
    .A3(_02884_),
    .B1(_04623_),
    .X(_02888_));
 sky130_fd_sc_hd__a2bb2o_1 _18903_ (.A1_N(_02887_),
    .A2_N(_02888_),
    .B1(\rbzero.wall_tracer.rayAddendY[5] ),
    .B2(_09932_),
    .X(_02889_));
 sky130_fd_sc_hd__a31o_1 _18904_ (.A1(_02529_),
    .A2(net4759),
    .A3(net7599),
    .B1(net3445),
    .X(_00609_));
 sky130_fd_sc_hd__xnor2_2 _18905_ (.A(_02854_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02890_));
 sky130_fd_sc_hd__a21o_1 _18906_ (.A1(net4662),
    .A2(_02883_),
    .B1(net7580),
    .X(_02891_));
 sky130_fd_sc_hd__nand3_1 _18907_ (.A(net4662),
    .B(_02883_),
    .C(_02890_),
    .Y(_02892_));
 sky130_fd_sc_hd__inv_2 _18908_ (.A(_02863_),
    .Y(_02893_));
 sky130_fd_sc_hd__inv_2 _18909_ (.A(net4459),
    .Y(_02894_));
 sky130_fd_sc_hd__or2_1 _18910_ (.A(_02863_),
    .B(net3700),
    .X(_02895_));
 sky130_fd_sc_hd__nand2_1 _18911_ (.A(_02863_),
    .B(net3700),
    .Y(_02896_));
 sky130_fd_sc_hd__a22o_1 _18912_ (.A1(_02893_),
    .A2(_02894_),
    .B1(_02895_),
    .B2(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__or3b_1 _18913_ (.A(_02863_),
    .B(net4459),
    .C_N(net3700),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _18914_ (.A(_02897_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__a21o_1 _18915_ (.A1(_02867_),
    .A2(_02885_),
    .B1(_02887_),
    .X(_02900_));
 sky130_fd_sc_hd__xnor2_1 _18916_ (.A(_02899_),
    .B(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__a22o_1 _18917_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(_09932_),
    .B1(_02901_),
    .B2(_04633_),
    .X(_02902_));
 sky130_fd_sc_hd__a31o_1 _18918_ (.A1(_02529_),
    .A2(net7581),
    .A3(net4663),
    .B1(net3481),
    .X(_00610_));
 sky130_fd_sc_hd__nand2_2 _18919_ (.A(_02863_),
    .B(net3090),
    .Y(_02903_));
 sky130_fd_sc_hd__or2_1 _18920_ (.A(_02863_),
    .B(net3090),
    .X(_02904_));
 sky130_fd_sc_hd__inv_2 _18921_ (.A(_02890_),
    .Y(_02905_));
 sky130_fd_sc_hd__o21a_1 _18922_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .B1(_02854_),
    .X(_02906_));
 sky130_fd_sc_hd__a311o_1 _18923_ (.A1(_02879_),
    .A2(_02880_),
    .A3(_02905_),
    .B1(net4816),
    .C1(net4758),
    .X(_02907_));
 sky130_fd_sc_hd__a21o_1 _18924_ (.A1(_02903_),
    .A2(_02904_),
    .B1(net4817),
    .X(_02908_));
 sky130_fd_sc_hd__nand3_2 _18925_ (.A(_02903_),
    .B(_02904_),
    .C(net4817),
    .Y(_02909_));
 sky130_fd_sc_hd__or2_1 _18926_ (.A(_02863_),
    .B(_05391_),
    .X(_02910_));
 sky130_fd_sc_hd__nand2_1 _18927_ (.A(_02864_),
    .B(_05391_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21bo_1 _18928_ (.A1(_02910_),
    .A2(_02911_),
    .B1_N(_02895_),
    .X(_02912_));
 sky130_fd_sc_hd__or3b_2 _18929_ (.A(_02864_),
    .B(net3700),
    .C_N(_05391_),
    .X(_02913_));
 sky130_fd_sc_hd__and3_1 _18930_ (.A(_02893_),
    .B(net3700),
    .C(_02894_),
    .X(_02914_));
 sky130_fd_sc_hd__and3_1 _18931_ (.A(_02897_),
    .B(_02898_),
    .C(_02900_),
    .X(_02915_));
 sky130_fd_sc_hd__a211o_1 _18932_ (.A1(_02912_),
    .A2(_02913_),
    .B1(_02914_),
    .C1(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__o211ai_2 _18933_ (.A1(_02914_),
    .A2(_02915_),
    .B1(_02912_),
    .C1(_02913_),
    .Y(_02917_));
 sky130_fd_sc_hd__a32o_1 _18934_ (.A1(_04633_),
    .A2(_02916_),
    .A3(_02917_),
    .B1(_09933_),
    .B2(net3090),
    .X(_02918_));
 sky130_fd_sc_hd__a31o_1 _18935_ (.A1(_02529_),
    .A2(net4818),
    .A3(_02909_),
    .B1(net3091),
    .X(_00611_));
 sky130_fd_sc_hd__nand2_1 _18936_ (.A(_02863_),
    .B(net3135),
    .Y(_02919_));
 sky130_fd_sc_hd__or2_1 _18937_ (.A(_02863_),
    .B(net3135),
    .X(_02920_));
 sky130_fd_sc_hd__nand2_1 _18938_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__a21oi_1 _18939_ (.A1(_02903_),
    .A2(_02909_),
    .B1(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__a31o_1 _18940_ (.A1(_02903_),
    .A2(_02909_),
    .A3(_02921_),
    .B1(_08246_),
    .X(_02923_));
 sky130_fd_sc_hd__or2_1 _18941_ (.A(_02864_),
    .B(net4634),
    .X(_02924_));
 sky130_fd_sc_hd__nand2_1 _18942_ (.A(_02864_),
    .B(net4634),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _18943_ (.A(_02924_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__xnor2_1 _18944_ (.A(_02910_),
    .B(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__a21oi_1 _18945_ (.A1(_02913_),
    .A2(_02917_),
    .B1(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__a31o_1 _18946_ (.A1(_02913_),
    .A2(_02917_),
    .A3(_02927_),
    .B1(_04623_),
    .X(_02929_));
 sky130_fd_sc_hd__o22ai_1 _18947_ (.A1(_02922_),
    .A2(_02923_),
    .B1(_02928_),
    .B2(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__mux2_1 _18948_ (.A0(net3135),
    .A1(_02930_),
    .S(_02714_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _18949_ (.A(net3136),
    .X(_00612_));
 sky130_fd_sc_hd__or2_1 _18950_ (.A(_02864_),
    .B(net3085),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_1 _18951_ (.A(_02864_),
    .B(net3085),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _18952_ (.A(_02932_),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__o211a_1 _18953_ (.A1(_02909_),
    .A2(_02921_),
    .B1(_02919_),
    .C1(_02903_),
    .X(_02935_));
 sky130_fd_sc_hd__xor2_1 _18954_ (.A(_02934_),
    .B(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__a211oi_1 _18955_ (.A1(net4634),
    .A2(_05391_),
    .B1(_02928_),
    .C1(_02864_),
    .Y(_02937_));
 sky130_fd_sc_hd__a211o_1 _18956_ (.A1(_02924_),
    .A2(_02928_),
    .B1(_02937_),
    .C1(_04624_),
    .X(_02938_));
 sky130_fd_sc_hd__o221a_1 _18957_ (.A1(net3085),
    .A2(_02557_),
    .B1(_09943_),
    .B2(_02936_),
    .C1(_02938_),
    .X(_00613_));
 sky130_fd_sc_hd__o21a_1 _18958_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02933_),
    .X(_02939_));
 sky130_fd_sc_hd__xor2_1 _18959_ (.A(_02864_),
    .B(net3018),
    .X(_02940_));
 sky130_fd_sc_hd__xnor2_1 _18960_ (.A(_02939_),
    .B(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__o311a_1 _18961_ (.A1(net4634),
    .A2(_05391_),
    .A3(_02917_),
    .B1(_08246_),
    .C1(_02893_),
    .X(_02942_));
 sky130_fd_sc_hd__a21o_1 _18962_ (.A1(_04624_),
    .A2(_02941_),
    .B1(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _18963_ (.A0(net3018),
    .A1(_02943_),
    .S(_02714_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _18964_ (.A(net3019),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _18965_ (.A0(net3821),
    .A1(_06219_),
    .S(_09999_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _18966_ (.A0(net3822),
    .A1(_06217_),
    .S(_01749_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _18967_ (.A(net3823),
    .X(_00615_));
 sky130_fd_sc_hd__or2_1 _18968_ (.A(_06217_),
    .B(_09950_),
    .X(_02947_));
 sky130_fd_sc_hd__nor2_1 _18969_ (.A(net3996),
    .B(_02261_),
    .Y(_02948_));
 sky130_fd_sc_hd__a31o_1 _18970_ (.A1(_02261_),
    .A2(_09951_),
    .A3(_02947_),
    .B1(net3997),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _18971_ (.A0(net3998),
    .A1(net6249),
    .S(_01749_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _18972_ (.A(net3999),
    .X(_00616_));
 sky130_fd_sc_hd__or2_1 _18973_ (.A(_09952_),
    .B(_09953_),
    .X(_02951_));
 sky130_fd_sc_hd__nor2_1 _18974_ (.A(_04823_),
    .B(_02261_),
    .Y(_02952_));
 sky130_fd_sc_hd__a31o_1 _18975_ (.A1(_02261_),
    .A2(_09954_),
    .A3(_02951_),
    .B1(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _18976_ (.A0(_02953_),
    .A1(net3984),
    .S(_01749_),
    .X(_02954_));
 sky130_fd_sc_hd__clkbuf_1 _18977_ (.A(net3985),
    .X(_00617_));
 sky130_fd_sc_hd__nand2_1 _18978_ (.A(_09956_),
    .B(_09949_),
    .Y(_02955_));
 sky130_fd_sc_hd__xnor2_1 _18979_ (.A(_09955_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__mux2_1 _18980_ (.A0(net3921),
    .A1(_02956_),
    .S(_09999_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _18981_ (.A0(net3922),
    .A1(net6217),
    .S(net4902),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_1 _18982_ (.A(net3923),
    .X(_00618_));
 sky130_fd_sc_hd__xor2_1 _18983_ (.A(_09948_),
    .B(_09957_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _18984_ (.A0(net3853),
    .A1(_02959_),
    .S(_09999_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _18985_ (.A0(net3854),
    .A1(net4874),
    .S(net4902),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _18986_ (.A(net3855),
    .X(_00619_));
 sky130_fd_sc_hd__a21oi_1 _18987_ (.A1(net4874),
    .A2(_09968_),
    .B1(_09974_),
    .Y(_02962_));
 sky130_fd_sc_hd__xnor2_1 _18988_ (.A(_09947_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__mux2_1 _18989_ (.A0(net6140),
    .A1(_02963_),
    .S(_09999_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _18990_ (.A0(net6141),
    .A1(net3265),
    .S(net4902),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _18991_ (.A(net3266),
    .X(_00620_));
 sky130_fd_sc_hd__and3_1 _18992_ (.A(net3747),
    .B(net3213),
    .C(net2978),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_2 _18993_ (.A(_02523_),
    .X(_02967_));
 sky130_fd_sc_hd__a21o_1 _18994_ (.A1(net3213),
    .A2(net2978),
    .B1(net3747),
    .X(_02968_));
 sky130_fd_sc_hd__and3b_1 _18995_ (.A_N(_02966_),
    .B(_02967_),
    .C(net3748),
    .X(_02969_));
 sky130_fd_sc_hd__clkbuf_1 _18996_ (.A(net3749),
    .X(_00621_));
 sky130_fd_sc_hd__and2_1 _18997_ (.A(net3889),
    .B(_02966_),
    .X(_02970_));
 sky130_fd_sc_hd__or2_1 _18998_ (.A(net3889),
    .B(_02966_),
    .X(_02971_));
 sky130_fd_sc_hd__and3b_1 _18999_ (.A_N(net7355),
    .B(_02967_),
    .C(net3890),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _19000_ (.A(net3891),
    .X(_00622_));
 sky130_fd_sc_hd__and3_1 _19001_ (.A(net3913),
    .B(net3889),
    .C(_02966_),
    .X(_02973_));
 sky130_fd_sc_hd__or2_1 _19002_ (.A(net3913),
    .B(_02970_),
    .X(_02974_));
 sky130_fd_sc_hd__and3b_1 _19003_ (.A_N(_02973_),
    .B(_02967_),
    .C(net3914),
    .X(_02975_));
 sky130_fd_sc_hd__clkbuf_1 _19004_ (.A(net3915),
    .X(_00623_));
 sky130_fd_sc_hd__and2_1 _19005_ (.A(net3904),
    .B(_02973_),
    .X(_02976_));
 sky130_fd_sc_hd__or2_1 _19006_ (.A(net3904),
    .B(_02973_),
    .X(_02977_));
 sky130_fd_sc_hd__and3b_1 _19007_ (.A_N(net7357),
    .B(_02967_),
    .C(net3905),
    .X(_02978_));
 sky130_fd_sc_hd__clkbuf_1 _19008_ (.A(net3906),
    .X(_00624_));
 sky130_fd_sc_hd__and3_1 _19009_ (.A(net3885),
    .B(net3904),
    .C(_02973_),
    .X(_02979_));
 sky130_fd_sc_hd__or2_1 _19010_ (.A(net3885),
    .B(_02976_),
    .X(_02980_));
 sky130_fd_sc_hd__and3b_1 _19011_ (.A_N(_02979_),
    .B(_02967_),
    .C(net3886),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_1 _19012_ (.A(net3887),
    .X(_00625_));
 sky130_fd_sc_hd__and2_1 _19013_ (.A(net3969),
    .B(_02979_),
    .X(_02982_));
 sky130_fd_sc_hd__or2_1 _19014_ (.A(net3374),
    .B(_02979_),
    .X(_02983_));
 sky130_fd_sc_hd__and3b_1 _19015_ (.A_N(_02982_),
    .B(_02523_),
    .C(net3375),
    .X(_02984_));
 sky130_fd_sc_hd__clkbuf_1 _19016_ (.A(net3376),
    .X(_00626_));
 sky130_fd_sc_hd__a21boi_1 _19017_ (.A1(net5619),
    .A2(_02982_),
    .B1_N(_02967_),
    .Y(_02985_));
 sky130_fd_sc_hd__o21a_1 _19018_ (.A1(net5619),
    .A2(_02982_),
    .B1(_02985_),
    .X(_00627_));
 sky130_fd_sc_hd__buf_1 _19019_ (.A(net6271),
    .X(_02986_));
 sky130_fd_sc_hd__nor3b_1 _19020_ (.A(net3945),
    .B(net88),
    .C_N(net2978),
    .Y(_02987_));
 sky130_fd_sc_hd__buf_2 _19021_ (.A(net2842),
    .X(_02988_));
 sky130_fd_sc_hd__or3b_1 _19022_ (.A(net3945),
    .B(net88),
    .C_N(net2978),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_2 _19023_ (.A(net2979),
    .X(_02990_));
 sky130_fd_sc_hd__or2_1 _19024_ (.A(net6307),
    .B(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_8 _19025_ (.A(_08274_),
    .X(_02992_));
 sky130_fd_sc_hd__buf_2 _19026_ (.A(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__o211a_1 _19027_ (.A1(net1572),
    .A2(_02988_),
    .B1(net1468),
    .C1(_02993_),
    .X(_00628_));
 sky130_fd_sc_hd__clkbuf_1 _19028_ (.A(net3949),
    .X(_02994_));
 sky130_fd_sc_hd__or2_1 _19029_ (.A(net1572),
    .B(_02990_),
    .X(_02995_));
 sky130_fd_sc_hd__o211a_1 _19030_ (.A1(net1608),
    .A2(_02988_),
    .B1(_02995_),
    .C1(_02993_),
    .X(_00629_));
 sky130_fd_sc_hd__buf_4 _19031_ (.A(net3957),
    .X(_02996_));
 sky130_fd_sc_hd__or2_1 _19032_ (.A(net1608),
    .B(_02990_),
    .X(_02997_));
 sky130_fd_sc_hd__o211a_1 _19033_ (.A1(net3958),
    .A2(_02988_),
    .B1(_02997_),
    .C1(_02993_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_4 _19034_ (.A(net3933),
    .X(_02998_));
 sky130_fd_sc_hd__or2_1 _19035_ (.A(_02996_),
    .B(_02990_),
    .X(_02999_));
 sky130_fd_sc_hd__o211a_1 _19036_ (.A1(net3934),
    .A2(_02988_),
    .B1(_02999_),
    .C1(_02993_),
    .X(_00631_));
 sky130_fd_sc_hd__buf_4 _19037_ (.A(net3940),
    .X(_03000_));
 sky130_fd_sc_hd__or2_1 _19038_ (.A(net3934),
    .B(_02990_),
    .X(_03001_));
 sky130_fd_sc_hd__o211a_1 _19039_ (.A1(net3941),
    .A2(_02988_),
    .B1(_03001_),
    .C1(_02993_),
    .X(_00632_));
 sky130_fd_sc_hd__clkbuf_1 _19040_ (.A(net6225),
    .X(_03002_));
 sky130_fd_sc_hd__or2_1 _19041_ (.A(net3941),
    .B(_02990_),
    .X(_03003_));
 sky130_fd_sc_hd__o211a_1 _19042_ (.A1(net1727),
    .A2(_02988_),
    .B1(net3942),
    .C1(_02993_),
    .X(_00633_));
 sky130_fd_sc_hd__or2_1 _19043_ (.A(net1727),
    .B(_02990_),
    .X(_03004_));
 sky130_fd_sc_hd__o211a_1 _19044_ (.A1(net3112),
    .A2(_02988_),
    .B1(_03004_),
    .C1(_02993_),
    .X(_00634_));
 sky130_fd_sc_hd__or2_1 _19045_ (.A(net3112),
    .B(_02990_),
    .X(_03005_));
 sky130_fd_sc_hd__o211a_1 _19046_ (.A1(net6164),
    .A2(_02988_),
    .B1(_03005_),
    .C1(_02993_),
    .X(_00635_));
 sky130_fd_sc_hd__or2_1 _19047_ (.A(net6164),
    .B(_02990_),
    .X(_03006_));
 sky130_fd_sc_hd__o211a_1 _19048_ (.A1(net6172),
    .A2(_02988_),
    .B1(_03006_),
    .C1(_02993_),
    .X(_00636_));
 sky130_fd_sc_hd__or2_1 _19049_ (.A(net6172),
    .B(_02990_),
    .X(_03007_));
 sky130_fd_sc_hd__o211a_1 _19050_ (.A1(net3096),
    .A2(_02988_),
    .B1(_03007_),
    .C1(_02993_),
    .X(_00637_));
 sky130_fd_sc_hd__clkbuf_1 _19051_ (.A(net2842),
    .X(_03008_));
 sky130_fd_sc_hd__buf_2 _19052_ (.A(net2979),
    .X(_03009_));
 sky130_fd_sc_hd__or2_1 _19053_ (.A(net3096),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_4 _19054_ (.A(_02992_),
    .X(_03011_));
 sky130_fd_sc_hd__o211a_1 _19055_ (.A1(net5838),
    .A2(net2843),
    .B1(net3097),
    .C1(_03011_),
    .X(_00638_));
 sky130_fd_sc_hd__or2_1 _19056_ (.A(net5838),
    .B(_03009_),
    .X(_03012_));
 sky130_fd_sc_hd__o211a_1 _19057_ (.A1(net3022),
    .A2(net2843),
    .B1(_03012_),
    .C1(_03011_),
    .X(_00639_));
 sky130_fd_sc_hd__or2_1 _19058_ (.A(net3022),
    .B(_03009_),
    .X(_03013_));
 sky130_fd_sc_hd__o211a_1 _19059_ (.A1(net3038),
    .A2(net2843),
    .B1(_03013_),
    .C1(_03011_),
    .X(_00640_));
 sky130_fd_sc_hd__or2_1 _19060_ (.A(net3038),
    .B(_03009_),
    .X(_03014_));
 sky130_fd_sc_hd__o211a_1 _19061_ (.A1(net3088),
    .A2(net2843),
    .B1(_03014_),
    .C1(_03011_),
    .X(_00641_));
 sky130_fd_sc_hd__or2_1 _19062_ (.A(net3088),
    .B(_03009_),
    .X(_03015_));
 sky130_fd_sc_hd__o211a_1 _19063_ (.A1(net3070),
    .A2(net2843),
    .B1(_03015_),
    .C1(_03011_),
    .X(_00642_));
 sky130_fd_sc_hd__or2_1 _19064_ (.A(net3070),
    .B(_03009_),
    .X(_03016_));
 sky130_fd_sc_hd__o211a_1 _19065_ (.A1(net3100),
    .A2(net2843),
    .B1(_03016_),
    .C1(_03011_),
    .X(_00643_));
 sky130_fd_sc_hd__or2_1 _19066_ (.A(net3100),
    .B(_03009_),
    .X(_03017_));
 sky130_fd_sc_hd__o211a_1 _19067_ (.A1(net6058),
    .A2(net2843),
    .B1(_03017_),
    .C1(_03011_),
    .X(_00644_));
 sky130_fd_sc_hd__or2_1 _19068_ (.A(net6058),
    .B(_03009_),
    .X(_03018_));
 sky130_fd_sc_hd__o211a_1 _19069_ (.A1(net6029),
    .A2(net2843),
    .B1(_03018_),
    .C1(_03011_),
    .X(_00645_));
 sky130_fd_sc_hd__or2_1 _19070_ (.A(net6029),
    .B(_03009_),
    .X(_03019_));
 sky130_fd_sc_hd__o211a_1 _19071_ (.A1(net3109),
    .A2(net2843),
    .B1(_03019_),
    .C1(_03011_),
    .X(_00646_));
 sky130_fd_sc_hd__or2_1 _19072_ (.A(net2970),
    .B(_03009_),
    .X(_03020_));
 sky130_fd_sc_hd__o211a_1 _19073_ (.A1(net6104),
    .A2(net2843),
    .B1(net2971),
    .C1(_03011_),
    .X(_00647_));
 sky130_fd_sc_hd__or2_1 _19074_ (.A(net642),
    .B(net2979),
    .X(_03021_));
 sky130_fd_sc_hd__buf_4 _19075_ (.A(_02992_),
    .X(_03022_));
 sky130_fd_sc_hd__o211a_1 _19076_ (.A1(net4318),
    .A2(net2842),
    .B1(net643),
    .C1(_03022_),
    .X(_00648_));
 sky130_fd_sc_hd__or2_1 _19077_ (.A(net4322),
    .B(net2979),
    .X(_03023_));
 sky130_fd_sc_hd__o211a_1 _19078_ (.A1(net4401),
    .A2(net2842),
    .B1(_03023_),
    .C1(_03022_),
    .X(_00649_));
 sky130_fd_sc_hd__or2_1 _19079_ (.A(net2962),
    .B(net2979),
    .X(_03024_));
 sky130_fd_sc_hd__o211a_1 _19080_ (.A1(net6047),
    .A2(net2842),
    .B1(net2980),
    .C1(_03022_),
    .X(_00650_));
 sky130_fd_sc_hd__or2_1 _19081_ (.A(net2948),
    .B(net2979),
    .X(_03025_));
 sky130_fd_sc_hd__o211a_1 _19082_ (.A1(net6033),
    .A2(net2842),
    .B1(net2949),
    .C1(_03022_),
    .X(_00651_));
 sky130_fd_sc_hd__buf_4 _19083_ (.A(_08274_),
    .X(_03026_));
 sky130_fd_sc_hd__and2_1 _19084_ (.A(net57),
    .B(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _19085_ (.A(_03027_),
    .X(_00652_));
 sky130_fd_sc_hd__and2_1 _19086_ (.A(net6324),
    .B(_03026_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _19087_ (.A(net622),
    .X(_00653_));
 sky130_fd_sc_hd__and2_1 _19088_ (.A(net4884),
    .B(_03026_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _19089_ (.A(net2123),
    .X(_00654_));
 sky130_fd_sc_hd__and3_1 _19090_ (.A(net4020),
    .B(net3897),
    .C(net3964),
    .X(_03030_));
 sky130_fd_sc_hd__nand2_1 _19091_ (.A(_05299_),
    .B(net3898),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2_2 _19092_ (.A(_09929_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__and4b_1 _19093_ (.A_N(net3937),
    .B(net3930),
    .C(net4002),
    .D(_04802_),
    .X(_03033_));
 sky130_fd_sc_hd__and4_2 _19094_ (.A(_04881_),
    .B(_05816_),
    .C(_03032_),
    .D(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_4 _19095_ (.A(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__buf_4 _19096_ (.A(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_4 _19097_ (.A(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__nand4_4 _19098_ (.A(_04881_),
    .B(_05816_),
    .C(_03032_),
    .D(_03033_),
    .Y(_03038_));
 sky130_fd_sc_hd__buf_4 _19099_ (.A(_03038_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_2 _19100_ (.A(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__or2_1 _19101_ (.A(net5255),
    .B(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__o211a_1 _19102_ (.A1(net5908),
    .A2(_03037_),
    .B1(_03041_),
    .C1(_03022_),
    .X(_00655_));
 sky130_fd_sc_hd__or2_1 _19103_ (.A(net5367),
    .B(_03040_),
    .X(_03042_));
 sky130_fd_sc_hd__o211a_1 _19104_ (.A1(net5944),
    .A2(_03037_),
    .B1(_03042_),
    .C1(_03022_),
    .X(_00656_));
 sky130_fd_sc_hd__or2_1 _19105_ (.A(net5562),
    .B(_03040_),
    .X(_03043_));
 sky130_fd_sc_hd__o211a_1 _19106_ (.A1(net6014),
    .A2(_03037_),
    .B1(_03043_),
    .C1(_03022_),
    .X(_00657_));
 sky130_fd_sc_hd__or2_1 _19107_ (.A(net5110),
    .B(_03040_),
    .X(_03044_));
 sky130_fd_sc_hd__o211a_1 _19108_ (.A1(net5808),
    .A2(_03037_),
    .B1(_03044_),
    .C1(_03022_),
    .X(_00658_));
 sky130_fd_sc_hd__or2_1 _19109_ (.A(net5402),
    .B(_03040_),
    .X(_03045_));
 sky130_fd_sc_hd__o211a_1 _19110_ (.A1(net5973),
    .A2(_03037_),
    .B1(_03045_),
    .C1(_03022_),
    .X(_00659_));
 sky130_fd_sc_hd__or2_1 _19111_ (.A(net5459),
    .B(_03040_),
    .X(_03046_));
 sky130_fd_sc_hd__o211a_1 _19112_ (.A1(net6017),
    .A2(_03037_),
    .B1(_03046_),
    .C1(_03022_),
    .X(_00660_));
 sky130_fd_sc_hd__or2_1 _19113_ (.A(net5406),
    .B(_03040_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_4 _19114_ (.A(_02992_),
    .X(_03048_));
 sky130_fd_sc_hd__o211a_1 _19115_ (.A1(net6005),
    .A2(_03037_),
    .B1(_03047_),
    .C1(_03048_),
    .X(_00661_));
 sky130_fd_sc_hd__or2_1 _19116_ (.A(net5124),
    .B(_03040_),
    .X(_03049_));
 sky130_fd_sc_hd__o211a_1 _19117_ (.A1(net5959),
    .A2(_03037_),
    .B1(_03049_),
    .C1(_03048_),
    .X(_00662_));
 sky130_fd_sc_hd__or2_1 _19118_ (.A(net5045),
    .B(_03040_),
    .X(_03050_));
 sky130_fd_sc_hd__o211a_1 _19119_ (.A1(net5876),
    .A2(_03037_),
    .B1(_03050_),
    .C1(_03048_),
    .X(_00663_));
 sky130_fd_sc_hd__or2_1 _19120_ (.A(net5375),
    .B(_03040_),
    .X(_03051_));
 sky130_fd_sc_hd__o211a_1 _19121_ (.A1(net5993),
    .A2(_03037_),
    .B1(_03051_),
    .C1(_03048_),
    .X(_00664_));
 sky130_fd_sc_hd__buf_2 _19122_ (.A(_03036_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_2 _19123_ (.A(_03039_),
    .X(_03053_));
 sky130_fd_sc_hd__or2_1 _19124_ (.A(net3864),
    .B(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__o211a_1 _19125_ (.A1(net4683),
    .A2(_03052_),
    .B1(_03054_),
    .C1(_03048_),
    .X(_00665_));
 sky130_fd_sc_hd__or2_1 _19126_ (.A(net5132),
    .B(_03053_),
    .X(_03055_));
 sky130_fd_sc_hd__o211a_1 _19127_ (.A1(net5966),
    .A2(_03052_),
    .B1(_03055_),
    .C1(_03048_),
    .X(_00666_));
 sky130_fd_sc_hd__or2_1 _19128_ (.A(net5190),
    .B(_03053_),
    .X(_03056_));
 sky130_fd_sc_hd__o211a_1 _19129_ (.A1(net5999),
    .A2(_03052_),
    .B1(_03056_),
    .C1(_03048_),
    .X(_00667_));
 sky130_fd_sc_hd__or2_1 _19130_ (.A(net5155),
    .B(_03053_),
    .X(_03057_));
 sky130_fd_sc_hd__o211a_1 _19131_ (.A1(net5950),
    .A2(_03052_),
    .B1(_03057_),
    .C1(_03048_),
    .X(_00668_));
 sky130_fd_sc_hd__or2_1 _19132_ (.A(net824),
    .B(_03053_),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _19133_ (.A1(net4345),
    .A2(_03052_),
    .B1(net631),
    .C1(_03048_),
    .X(_00669_));
 sky130_fd_sc_hd__or2_1 _19134_ (.A(net930),
    .B(_03053_),
    .X(_03059_));
 sky130_fd_sc_hd__o211a_1 _19135_ (.A1(net5699),
    .A2(_03052_),
    .B1(net637),
    .C1(_03048_),
    .X(_00670_));
 sky130_fd_sc_hd__or2_1 _19136_ (.A(net5099),
    .B(_03053_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_4 _19137_ (.A(_02992_),
    .X(_03061_));
 sky130_fd_sc_hd__o211a_1 _19138_ (.A1(net5559),
    .A2(_03052_),
    .B1(_03060_),
    .C1(_03061_),
    .X(_00671_));
 sky130_fd_sc_hd__or2_1 _19139_ (.A(net5065),
    .B(_03053_),
    .X(_03062_));
 sky130_fd_sc_hd__o211a_1 _19140_ (.A1(net5918),
    .A2(_03052_),
    .B1(_03062_),
    .C1(_03061_),
    .X(_00672_));
 sky130_fd_sc_hd__or2_1 _19141_ (.A(net5371),
    .B(_03053_),
    .X(_03063_));
 sky130_fd_sc_hd__o211a_1 _19142_ (.A1(net6002),
    .A2(_03052_),
    .B1(_03063_),
    .C1(_03061_),
    .X(_00673_));
 sky130_fd_sc_hd__or2_1 _19143_ (.A(net5216),
    .B(_03053_),
    .X(_03064_));
 sky130_fd_sc_hd__o211a_1 _19144_ (.A1(net5978),
    .A2(_03052_),
    .B1(_03064_),
    .C1(_03061_),
    .X(_00674_));
 sky130_fd_sc_hd__clkbuf_4 _19145_ (.A(_03036_),
    .X(_03065_));
 sky130_fd_sc_hd__buf_2 _19146_ (.A(_03039_),
    .X(_03066_));
 sky130_fd_sc_hd__or2_1 _19147_ (.A(net5014),
    .B(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__o211a_1 _19148_ (.A1(net5947),
    .A2(_03065_),
    .B1(_03067_),
    .C1(_03061_),
    .X(_00675_));
 sky130_fd_sc_hd__or2_1 _19149_ (.A(net5186),
    .B(_03066_),
    .X(_03068_));
 sky130_fd_sc_hd__o211a_1 _19150_ (.A1(net5939),
    .A2(_03065_),
    .B1(_03068_),
    .C1(_03061_),
    .X(_00676_));
 sky130_fd_sc_hd__or2_1 _19151_ (.A(net5079),
    .B(_03066_),
    .X(_03069_));
 sky130_fd_sc_hd__o211a_1 _19152_ (.A1(net5733),
    .A2(_03065_),
    .B1(_03069_),
    .C1(_03061_),
    .X(_00677_));
 sky130_fd_sc_hd__or2_1 _19153_ (.A(net5322),
    .B(_03066_),
    .X(_03070_));
 sky130_fd_sc_hd__o211a_1 _19154_ (.A1(net5497),
    .A2(_03065_),
    .B1(_03070_),
    .C1(_03061_),
    .X(_00678_));
 sky130_fd_sc_hd__or2_1 _19155_ (.A(net5283),
    .B(_03066_),
    .X(_03071_));
 sky130_fd_sc_hd__o211a_1 _19156_ (.A1(net5447),
    .A2(_03065_),
    .B1(_03071_),
    .C1(_03061_),
    .X(_00679_));
 sky130_fd_sc_hd__or2_1 _19157_ (.A(net5243),
    .B(_03066_),
    .X(_03072_));
 sky130_fd_sc_hd__o211a_1 _19158_ (.A1(net5442),
    .A2(_03065_),
    .B1(_03072_),
    .C1(_03061_),
    .X(_00680_));
 sky130_fd_sc_hd__or2_1 _19159_ (.A(net5279),
    .B(_03066_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_4 _19160_ (.A(_02992_),
    .X(_03074_));
 sky130_fd_sc_hd__o211a_1 _19161_ (.A1(net5678),
    .A2(_03065_),
    .B1(_03073_),
    .C1(_03074_),
    .X(_00681_));
 sky130_fd_sc_hd__or2_1 _19162_ (.A(net2541),
    .B(_03066_),
    .X(_03075_));
 sky130_fd_sc_hd__o211a_1 _19163_ (.A1(net5513),
    .A2(_03065_),
    .B1(_03075_),
    .C1(_03074_),
    .X(_00682_));
 sky130_fd_sc_hd__or2_1 _19164_ (.A(net1141),
    .B(_03066_),
    .X(_03076_));
 sky130_fd_sc_hd__o211a_1 _19165_ (.A1(net4197),
    .A2(_03065_),
    .B1(net1142),
    .C1(_03074_),
    .X(_00683_));
 sky130_fd_sc_hd__or2_1 _19166_ (.A(net2553),
    .B(_03066_),
    .X(_03077_));
 sky130_fd_sc_hd__o211a_1 _19167_ (.A1(net5710),
    .A2(_03065_),
    .B1(_03077_),
    .C1(_03074_),
    .X(_00684_));
 sky130_fd_sc_hd__clkbuf_4 _19168_ (.A(_03036_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_4 _19169_ (.A(_03039_),
    .X(_03079_));
 sky130_fd_sc_hd__or2_1 _19170_ (.A(net1735),
    .B(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__o211a_1 _19171_ (.A1(net5656),
    .A2(_03078_),
    .B1(_03080_),
    .C1(_03074_),
    .X(_00685_));
 sky130_fd_sc_hd__or2_1 _19172_ (.A(net2590),
    .B(_03079_),
    .X(_03081_));
 sky130_fd_sc_hd__o211a_1 _19173_ (.A1(net5702),
    .A2(_03078_),
    .B1(_03081_),
    .C1(_03074_),
    .X(_00686_));
 sky130_fd_sc_hd__or2_1 _19174_ (.A(net5783),
    .B(_03079_),
    .X(_03082_));
 sky130_fd_sc_hd__o211a_1 _19175_ (.A1(net5996),
    .A2(_03078_),
    .B1(net1635),
    .C1(_03074_),
    .X(_00687_));
 sky130_fd_sc_hd__clkbuf_8 _19176_ (.A(_04597_),
    .X(_03083_));
 sky130_fd_sc_hd__buf_4 _19177_ (.A(_03038_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _19178_ (.A0(net3254),
    .A1(net3144),
    .S(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__or2_1 _19179_ (.A(_03083_),
    .B(net3145),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _19180_ (.A(net3146),
    .X(_00688_));
 sky130_fd_sc_hd__or2_1 _19181_ (.A(net1595),
    .B(_03079_),
    .X(_03087_));
 sky130_fd_sc_hd__o211a_1 _19182_ (.A1(net5117),
    .A2(_03078_),
    .B1(_03087_),
    .C1(_03074_),
    .X(_00689_));
 sky130_fd_sc_hd__buf_2 _19183_ (.A(_04597_),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _19184_ (.A0(net2964),
    .A1(net7322),
    .S(_03084_),
    .X(_03089_));
 sky130_fd_sc_hd__or2_1 _19185_ (.A(_03088_),
    .B(net2965),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _19186_ (.A(net2966),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _19187_ (.A(net1531),
    .B(_03079_),
    .X(_03091_));
 sky130_fd_sc_hd__o211a_1 _19188_ (.A1(net5068),
    .A2(_03078_),
    .B1(_03091_),
    .C1(_03074_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _19189_ (.A0(net2995),
    .A1(net4081),
    .S(_03084_),
    .X(_03092_));
 sky130_fd_sc_hd__or2_1 _19190_ (.A(_03088_),
    .B(net2996),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _19191_ (.A(net2997),
    .X(_00692_));
 sky130_fd_sc_hd__or2_1 _19192_ (.A(net1790),
    .B(_03079_),
    .X(_03094_));
 sky130_fd_sc_hd__o211a_1 _19193_ (.A1(net5356),
    .A2(_03078_),
    .B1(_03094_),
    .C1(_03074_),
    .X(_00693_));
 sky130_fd_sc_hd__or2_1 _19194_ (.A(net1534),
    .B(_03079_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_4 _19195_ (.A(_02992_),
    .X(_03096_));
 sky130_fd_sc_hd__o211a_1 _19196_ (.A1(net5330),
    .A2(_03078_),
    .B1(_03095_),
    .C1(_03096_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _19197_ (.A0(net2973),
    .A1(net7325),
    .S(_03084_),
    .X(_03097_));
 sky130_fd_sc_hd__or2_1 _19198_ (.A(_03088_),
    .B(net2974),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _19199_ (.A(net2975),
    .X(_00695_));
 sky130_fd_sc_hd__or2_1 _19200_ (.A(net1615),
    .B(_03079_),
    .X(_03099_));
 sky130_fd_sc_hd__o211a_1 _19201_ (.A1(net5326),
    .A2(_03078_),
    .B1(_03099_),
    .C1(_03096_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _19202_ (.A0(net2951),
    .A1(net7327),
    .S(_03084_),
    .X(_03100_));
 sky130_fd_sc_hd__or2_1 _19203_ (.A(_03088_),
    .B(net2952),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _19204_ (.A(net2953),
    .X(_00697_));
 sky130_fd_sc_hd__or2_1 _19205_ (.A(net1540),
    .B(_03079_),
    .X(_03102_));
 sky130_fd_sc_hd__o211a_1 _19206_ (.A1(net5151),
    .A2(_03078_),
    .B1(_03102_),
    .C1(_03096_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _19207_ (.A0(net3116),
    .A1(net3128),
    .S(_03038_),
    .X(_03103_));
 sky130_fd_sc_hd__or2_1 _19208_ (.A(_03088_),
    .B(net3129),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _19209_ (.A(net3130),
    .X(_00699_));
 sky130_fd_sc_hd__or2_1 _19210_ (.A(net5247),
    .B(_03079_),
    .X(_03105_));
 sky130_fd_sc_hd__o211a_1 _19211_ (.A1(net5773),
    .A2(_03078_),
    .B1(_03105_),
    .C1(_03096_),
    .X(_00700_));
 sky130_fd_sc_hd__clkbuf_4 _19212_ (.A(_03036_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_4 _19213_ (.A(_03039_),
    .X(_03107_));
 sky130_fd_sc_hd__or2_1 _19214_ (.A(net5428),
    .B(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__o211a_1 _19215_ (.A1(net5721),
    .A2(_03106_),
    .B1(_03108_),
    .C1(_03096_),
    .X(_00701_));
 sky130_fd_sc_hd__or2_1 _19216_ (.A(net5547),
    .B(_03107_),
    .X(_03109_));
 sky130_fd_sc_hd__o211a_1 _19217_ (.A1(net5780),
    .A2(_03106_),
    .B1(_03109_),
    .C1(_03096_),
    .X(_00702_));
 sky130_fd_sc_hd__or2_1 _19218_ (.A(net5178),
    .B(_03107_),
    .X(_03110_));
 sky130_fd_sc_hd__o211a_1 _19219_ (.A1(net5852),
    .A2(_03106_),
    .B1(_03110_),
    .C1(_03096_),
    .X(_00703_));
 sky130_fd_sc_hd__or2_1 _19220_ (.A(net5302),
    .B(_03107_),
    .X(_03111_));
 sky130_fd_sc_hd__o211a_1 _19221_ (.A1(net5883),
    .A2(_03106_),
    .B1(_03111_),
    .C1(_03096_),
    .X(_00704_));
 sky130_fd_sc_hd__or2_1 _19222_ (.A(net5360),
    .B(_03107_),
    .X(_03112_));
 sky130_fd_sc_hd__o211a_1 _19223_ (.A1(net5802),
    .A2(_03106_),
    .B1(_03112_),
    .C1(_03096_),
    .X(_00705_));
 sky130_fd_sc_hd__or2_1 _19224_ (.A(net5087),
    .B(_03107_),
    .X(_03113_));
 sky130_fd_sc_hd__o211a_1 _19225_ (.A1(net5740),
    .A2(_03106_),
    .B1(_03113_),
    .C1(_03096_),
    .X(_00706_));
 sky130_fd_sc_hd__or2_1 _19226_ (.A(net5072),
    .B(_03107_),
    .X(_03114_));
 sky130_fd_sc_hd__clkbuf_4 _19227_ (.A(_02992_),
    .X(_03115_));
 sky130_fd_sc_hd__o211a_1 _19228_ (.A1(net5788),
    .A2(_03106_),
    .B1(_03114_),
    .C1(_03115_),
    .X(_00707_));
 sky130_fd_sc_hd__or2_1 _19229_ (.A(net5226),
    .B(_03107_),
    .X(_03116_));
 sky130_fd_sc_hd__o211a_1 _19230_ (.A1(net5669),
    .A2(_03106_),
    .B1(_03116_),
    .C1(_03115_),
    .X(_00708_));
 sky130_fd_sc_hd__or2_1 _19231_ (.A(net5236),
    .B(_03107_),
    .X(_03117_));
 sky130_fd_sc_hd__o211a_1 _19232_ (.A1(net5743),
    .A2(_03106_),
    .B1(_03117_),
    .C1(_03115_),
    .X(_00709_));
 sky130_fd_sc_hd__or2_1 _19233_ (.A(net5057),
    .B(_03107_),
    .X(_03118_));
 sky130_fd_sc_hd__o211a_1 _19234_ (.A1(net5609),
    .A2(_03106_),
    .B1(_03118_),
    .C1(_03115_),
    .X(_00710_));
 sky130_fd_sc_hd__clkbuf_4 _19235_ (.A(_03036_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_2 _19236_ (.A(_03039_),
    .X(_03120_));
 sky130_fd_sc_hd__or2_1 _19237_ (.A(net5318),
    .B(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__o211a_1 _19238_ (.A1(net5639),
    .A2(_03119_),
    .B1(_03121_),
    .C1(_03115_),
    .X(_00711_));
 sky130_fd_sc_hd__or2_1 _19239_ (.A(net809),
    .B(_03120_),
    .X(_03122_));
 sky130_fd_sc_hd__o211a_1 _19240_ (.A1(net5128),
    .A2(_03119_),
    .B1(_03122_),
    .C1(_03115_),
    .X(_00712_));
 sky130_fd_sc_hd__or2_1 _19241_ (.A(net5201),
    .B(_03120_),
    .X(_03123_));
 sky130_fd_sc_hd__o211a_1 _19242_ (.A1(net5230),
    .A2(_03119_),
    .B1(_03123_),
    .C1(_03115_),
    .X(_00713_));
 sky130_fd_sc_hd__or2_1 _19243_ (.A(net5222),
    .B(_03120_),
    .X(_03124_));
 sky130_fd_sc_hd__o211a_1 _19244_ (.A1(net5353),
    .A2(_03119_),
    .B1(_03124_),
    .C1(_03115_),
    .X(_00714_));
 sky130_fd_sc_hd__or2_1 _19245_ (.A(net5391),
    .B(_03120_),
    .X(_03125_));
 sky130_fd_sc_hd__o211a_1 _19246_ (.A1(net5649),
    .A2(_03119_),
    .B1(_03125_),
    .C1(_03115_),
    .X(_00715_));
 sky130_fd_sc_hd__or2_1 _19247_ (.A(net5030),
    .B(_03120_),
    .X(_03126_));
 sky130_fd_sc_hd__o211a_1 _19248_ (.A1(net5172),
    .A2(_03119_),
    .B1(_03126_),
    .C1(_03115_),
    .X(_00716_));
 sky130_fd_sc_hd__or2_1 _19249_ (.A(net603),
    .B(_03120_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_4 _19250_ (.A(_02992_),
    .X(_03128_));
 sky130_fd_sc_hd__o211a_1 _19251_ (.A1(net4121),
    .A2(_03119_),
    .B1(net604),
    .C1(_03128_),
    .X(_00717_));
 sky130_fd_sc_hd__or2_1 _19252_ (.A(net969),
    .B(_03120_),
    .X(_03129_));
 sky130_fd_sc_hd__o211a_1 _19253_ (.A1(net4149),
    .A2(_03119_),
    .B1(net610),
    .C1(_03128_),
    .X(_00718_));
 sky130_fd_sc_hd__or2_1 _19254_ (.A(net4115),
    .B(_03120_),
    .X(_03130_));
 sky130_fd_sc_hd__o211a_1 _19255_ (.A1(net4248),
    .A2(_03119_),
    .B1(_03130_),
    .C1(_03128_),
    .X(_00719_));
 sky130_fd_sc_hd__or2_1 _19256_ (.A(net606),
    .B(_03120_),
    .X(_03131_));
 sky130_fd_sc_hd__o211a_1 _19257_ (.A1(net4127),
    .A2(_03119_),
    .B1(net607),
    .C1(_03128_),
    .X(_00720_));
 sky130_fd_sc_hd__clkbuf_4 _19258_ (.A(_03036_),
    .X(_03132_));
 sky130_fd_sc_hd__clkbuf_4 _19259_ (.A(_03039_),
    .X(_03133_));
 sky130_fd_sc_hd__or2_1 _19260_ (.A(net5011),
    .B(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__o211a_1 _19261_ (.A1(net5395),
    .A2(_03132_),
    .B1(_03134_),
    .C1(_03128_),
    .X(_00721_));
 sky130_fd_sc_hd__or2_1 _19262_ (.A(net5061),
    .B(_03133_),
    .X(_03135_));
 sky130_fd_sc_hd__o211a_1 _19263_ (.A1(net5417),
    .A2(_03132_),
    .B1(_03135_),
    .C1(_03128_),
    .X(_00722_));
 sky130_fd_sc_hd__or2_1 _19264_ (.A(net4991),
    .B(_03133_),
    .X(_03136_));
 sky130_fd_sc_hd__o211a_1 _19265_ (.A1(net5165),
    .A2(_03132_),
    .B1(_03136_),
    .C1(_03128_),
    .X(_00723_));
 sky130_fd_sc_hd__or2_1 _19266_ (.A(net5140),
    .B(_03133_),
    .X(_03137_));
 sky130_fd_sc_hd__o211a_1 _19267_ (.A1(net5452),
    .A2(_03132_),
    .B1(_03137_),
    .C1(_03128_),
    .X(_00724_));
 sky130_fd_sc_hd__or2_1 _19268_ (.A(net5161),
    .B(_03133_),
    .X(_03138_));
 sky130_fd_sc_hd__o211a_1 _19269_ (.A1(net5681),
    .A2(_03132_),
    .B1(_03138_),
    .C1(_03128_),
    .X(_00725_));
 sky130_fd_sc_hd__or2_1 _19270_ (.A(net4607),
    .B(_03133_),
    .X(_03139_));
 sky130_fd_sc_hd__o211a_1 _19271_ (.A1(net5042),
    .A2(_03132_),
    .B1(_03139_),
    .C1(_03128_),
    .X(_00726_));
 sky130_fd_sc_hd__or2_1 _19272_ (.A(net5034),
    .B(_03133_),
    .X(_03140_));
 sky130_fd_sc_hd__buf_4 _19273_ (.A(_08274_),
    .X(_03141_));
 sky130_fd_sc_hd__buf_2 _19274_ (.A(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__o211a_1 _19275_ (.A1(net5076),
    .A2(_03132_),
    .B1(_03140_),
    .C1(_03142_),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _19276_ (.A(net5095),
    .B(_03133_),
    .X(_03143_));
 sky130_fd_sc_hd__o211a_1 _19277_ (.A1(net5295),
    .A2(_03132_),
    .B1(_03143_),
    .C1(_03142_),
    .X(_00728_));
 sky130_fd_sc_hd__or2_1 _19278_ (.A(net5038),
    .B(_03133_),
    .X(_03144_));
 sky130_fd_sc_hd__o211a_1 _19279_ (.A1(net5364),
    .A2(_03132_),
    .B1(_03144_),
    .C1(_03142_),
    .X(_00729_));
 sky130_fd_sc_hd__or2_1 _19280_ (.A(net1703),
    .B(_03133_),
    .X(_03145_));
 sky130_fd_sc_hd__o211a_1 _19281_ (.A1(net5298),
    .A2(_03132_),
    .B1(_03145_),
    .C1(_03142_),
    .X(_00730_));
 sky130_fd_sc_hd__clkbuf_4 _19282_ (.A(_03036_),
    .X(_03146_));
 sky130_fd_sc_hd__buf_2 _19283_ (.A(_03039_),
    .X(_03147_));
 sky130_fd_sc_hd__or2_1 _19284_ (.A(net1652),
    .B(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__o211a_1 _19285_ (.A1(net5306),
    .A2(_03146_),
    .B1(_03148_),
    .C1(_03142_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _19286_ (.A(net2076),
    .B(_03147_),
    .X(_03149_));
 sky130_fd_sc_hd__o211a_1 _19287_ (.A1(net5267),
    .A2(_03146_),
    .B1(_03149_),
    .C1(_03142_),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _19288_ (.A(net1667),
    .B(_03147_),
    .X(_03150_));
 sky130_fd_sc_hd__o211a_1 _19289_ (.A1(net5477),
    .A2(_03146_),
    .B1(_03150_),
    .C1(_03142_),
    .X(_00733_));
 sky130_fd_sc_hd__or2_1 _19290_ (.A(net1829),
    .B(_03147_),
    .X(_03151_));
 sky130_fd_sc_hd__o211a_1 _19291_ (.A1(net5342),
    .A2(_03146_),
    .B1(_03151_),
    .C1(_03142_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _19292_ (.A(net1604),
    .B(_03147_),
    .X(_03152_));
 sky130_fd_sc_hd__o211a_1 _19293_ (.A1(net5136),
    .A2(_03146_),
    .B1(_03152_),
    .C1(_03142_),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _19294_ (.A(net2274),
    .B(_03147_),
    .X(_03153_));
 sky130_fd_sc_hd__o211a_1 _19295_ (.A1(net5026),
    .A2(_03146_),
    .B1(_03153_),
    .C1(_03142_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _19296_ (.A(net2090),
    .B(_03147_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_4 _19297_ (.A(_03141_),
    .X(_03155_));
 sky130_fd_sc_hd__o211a_1 _19298_ (.A1(net5022),
    .A2(_03146_),
    .B1(_03154_),
    .C1(_03155_),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _19299_ (.A(net2256),
    .B(_03147_),
    .X(_03156_));
 sky130_fd_sc_hd__o211a_1 _19300_ (.A1(net4995),
    .A2(_03146_),
    .B1(_03156_),
    .C1(_03155_),
    .X(_00738_));
 sky130_fd_sc_hd__or2_1 _19301_ (.A(net1912),
    .B(_03147_),
    .X(_03157_));
 sky130_fd_sc_hd__o211a_1 _19302_ (.A1(net4983),
    .A2(_03146_),
    .B1(_03157_),
    .C1(_03155_),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _19303_ (.A(net3011),
    .B(_03147_),
    .X(_03158_));
 sky130_fd_sc_hd__o211a_1 _19304_ (.A1(net4124),
    .A2(_03146_),
    .B1(net619),
    .C1(_03155_),
    .X(_00740_));
 sky130_fd_sc_hd__clkbuf_4 _19305_ (.A(_03036_),
    .X(_03159_));
 sky130_fd_sc_hd__buf_2 _19306_ (.A(_03039_),
    .X(_03160_));
 sky130_fd_sc_hd__or2_1 _19307_ (.A(net1647),
    .B(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__o211a_1 _19308_ (.A1(net5259),
    .A2(_03159_),
    .B1(_03161_),
    .C1(_03155_),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _19309_ (.A(net1625),
    .B(_03160_),
    .X(_03162_));
 sky130_fd_sc_hd__o211a_1 _19310_ (.A1(net5182),
    .A2(_03159_),
    .B1(_03162_),
    .C1(_03155_),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _19311_ (.A(net1692),
    .B(_03160_),
    .X(_03163_));
 sky130_fd_sc_hd__o211a_1 _19312_ (.A1(net5614),
    .A2(_03159_),
    .B1(_03163_),
    .C1(_03155_),
    .X(_00743_));
 sky130_fd_sc_hd__or2_1 _19313_ (.A(net2593),
    .B(_03160_),
    .X(_03164_));
 sky130_fd_sc_hd__o211a_1 _19314_ (.A1(net5083),
    .A2(_03159_),
    .B1(_03164_),
    .C1(_03155_),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _19315_ (.A(net2487),
    .B(_03160_),
    .X(_03165_));
 sky130_fd_sc_hd__o211a_1 _19316_ (.A1(net5053),
    .A2(_03159_),
    .B1(_03165_),
    .C1(_03155_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _19317_ (.A(net4214),
    .B(_03160_),
    .X(_03166_));
 sky130_fd_sc_hd__o211a_1 _19318_ (.A1(net794),
    .A2(_03159_),
    .B1(net4215),
    .C1(_03155_),
    .X(_00746_));
 sky130_fd_sc_hd__or2_1 _19319_ (.A(net1859),
    .B(_03160_),
    .X(_03167_));
 sky130_fd_sc_hd__clkbuf_4 _19320_ (.A(_03141_),
    .X(_03168_));
 sky130_fd_sc_hd__o211a_1 _19321_ (.A1(net5314),
    .A2(_03159_),
    .B1(_03167_),
    .C1(_03168_),
    .X(_00747_));
 sky130_fd_sc_hd__or2_1 _19322_ (.A(net1729),
    .B(_03160_),
    .X(_03169_));
 sky130_fd_sc_hd__o211a_1 _19323_ (.A1(net5007),
    .A2(_03159_),
    .B1(_03169_),
    .C1(_03168_),
    .X(_00748_));
 sky130_fd_sc_hd__or2_1 _19324_ (.A(net1768),
    .B(_03160_),
    .X(_03170_));
 sky130_fd_sc_hd__o211a_1 _19325_ (.A1(net5275),
    .A2(_03159_),
    .B1(_03170_),
    .C1(_03168_),
    .X(_00749_));
 sky130_fd_sc_hd__or2_1 _19326_ (.A(net4672),
    .B(_03160_),
    .X(_03171_));
 sky130_fd_sc_hd__o211a_1 _19327_ (.A1(net5158),
    .A2(_03159_),
    .B1(_03171_),
    .C1(_03168_),
    .X(_00750_));
 sky130_fd_sc_hd__clkbuf_4 _19328_ (.A(_03035_),
    .X(_03172_));
 sky130_fd_sc_hd__buf_2 _19329_ (.A(_03084_),
    .X(_03173_));
 sky130_fd_sc_hd__or2_1 _19330_ (.A(net1712),
    .B(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__o211a_1 _19331_ (.A1(net5660),
    .A2(_03172_),
    .B1(_03174_),
    .C1(_03168_),
    .X(_00751_));
 sky130_fd_sc_hd__or2_1 _19332_ (.A(net1670),
    .B(_03173_),
    .X(_03175_));
 sky130_fd_sc_hd__o211a_1 _19333_ (.A1(net5714),
    .A2(_03172_),
    .B1(_03175_),
    .C1(_03168_),
    .X(_00752_));
 sky130_fd_sc_hd__or2_1 _19334_ (.A(net1548),
    .B(_03173_),
    .X(_03176_));
 sky130_fd_sc_hd__o211a_1 _19335_ (.A1(net5724),
    .A2(_03172_),
    .B1(_03176_),
    .C1(_03168_),
    .X(_00753_));
 sky130_fd_sc_hd__or2_1 _19336_ (.A(net1083),
    .B(_03173_),
    .X(_03177_));
 sky130_fd_sc_hd__o211a_1 _19337_ (.A1(net4191),
    .A2(_03172_),
    .B1(net1084),
    .C1(_03168_),
    .X(_00754_));
 sky130_fd_sc_hd__or2_1 _19338_ (.A(net1909),
    .B(_03173_),
    .X(_03178_));
 sky130_fd_sc_hd__o211a_1 _19339_ (.A1(net5594),
    .A2(_03172_),
    .B1(_03178_),
    .C1(_03168_),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _19340_ (.A(net1787),
    .B(_03173_),
    .X(_03179_));
 sky130_fd_sc_hd__o211a_1 _19341_ (.A1(net5642),
    .A2(_03172_),
    .B1(_03179_),
    .C1(_03168_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _19342_ (.A(net1868),
    .B(_03173_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_4 _19343_ (.A(_03141_),
    .X(_03181_));
 sky130_fd_sc_hd__o211a_1 _19344_ (.A1(net5652),
    .A2(_03172_),
    .B1(_03180_),
    .C1(_03181_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _19345_ (.A(net2113),
    .B(_03173_),
    .X(_03182_));
 sky130_fd_sc_hd__o211a_1 _19346_ (.A1(net5633),
    .A2(_03172_),
    .B1(_03182_),
    .C1(_03181_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _19347_ (.A(net1883),
    .B(_03173_),
    .X(_03183_));
 sky130_fd_sc_hd__o211a_1 _19348_ (.A1(net5674),
    .A2(_03172_),
    .B1(_03183_),
    .C1(_03181_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _19349_ (.A(net1217),
    .B(_03173_),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _19350_ (.A1(net4211),
    .A2(_03172_),
    .B1(net1218),
    .C1(_03181_),
    .X(_00760_));
 sky130_fd_sc_hd__clkbuf_4 _19351_ (.A(_03035_),
    .X(_03185_));
 sky130_fd_sc_hd__buf_2 _19352_ (.A(_03084_),
    .X(_03186_));
 sky130_fd_sc_hd__or2_1 _19353_ (.A(net2455),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__o211a_1 _19354_ (.A1(net5736),
    .A2(_03185_),
    .B1(_03187_),
    .C1(_03181_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19355_ (.A(net2533),
    .B(_03186_),
    .X(_03188_));
 sky130_fd_sc_hd__o211a_1 _19356_ (.A1(net5758),
    .A2(_03185_),
    .B1(_03188_),
    .C1(_03181_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19357_ (.A(net1806),
    .B(_03186_),
    .X(_03189_));
 sky130_fd_sc_hd__o211a_1 _19358_ (.A1(net5750),
    .A2(_03185_),
    .B1(_03189_),
    .C1(_03181_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _19359_ (.A(net4257),
    .B(_03186_),
    .X(_03190_));
 sky130_fd_sc_hd__o211a_1 _19360_ (.A1(net4268),
    .A2(_03185_),
    .B1(_03190_),
    .C1(_03181_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _19361_ (.A(net4243),
    .B(_03186_),
    .X(_03191_));
 sky130_fd_sc_hd__o211a_1 _19362_ (.A1(net1959),
    .A2(_03185_),
    .B1(net4244),
    .C1(_03181_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _19363_ (.A(net1655),
    .B(_03186_),
    .X(_03192_));
 sky130_fd_sc_hd__o211a_1 _19364_ (.A1(net4227),
    .A2(_03185_),
    .B1(net1656),
    .C1(_03181_),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _19365_ (.A(net2094),
    .B(_03186_),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_4 _19366_ (.A(_03141_),
    .X(_03194_));
 sky130_fd_sc_hd__o211a_1 _19367_ (.A1(net4261),
    .A2(_03185_),
    .B1(net592),
    .C1(_03194_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _19368_ (.A(net1563),
    .B(_03186_),
    .X(_03195_));
 sky130_fd_sc_hd__o211a_1 _19369_ (.A1(net4291),
    .A2(_03185_),
    .B1(net595),
    .C1(_03194_),
    .X(_00768_));
 sky130_fd_sc_hd__or2_1 _19370_ (.A(net1214),
    .B(_03186_),
    .X(_03196_));
 sky130_fd_sc_hd__o211a_1 _19371_ (.A1(net4208),
    .A2(_03185_),
    .B1(net1215),
    .C1(_03194_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _19372_ (.A(net1784),
    .B(_03186_),
    .X(_03197_));
 sky130_fd_sc_hd__o211a_1 _19373_ (.A1(net4205),
    .A2(_03185_),
    .B1(net1407),
    .C1(_03194_),
    .X(_00770_));
 sky130_fd_sc_hd__clkbuf_4 _19374_ (.A(_03035_),
    .X(_03198_));
 sky130_fd_sc_hd__buf_2 _19375_ (.A(_03084_),
    .X(_03199_));
 sky130_fd_sc_hd__or2_1 _19376_ (.A(net1644),
    .B(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__o211a_1 _19377_ (.A1(net5504),
    .A2(_03198_),
    .B1(_03200_),
    .C1(_03194_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _19378_ (.A(net2020),
    .B(_03199_),
    .X(_03201_));
 sky130_fd_sc_hd__o211a_1 _19379_ (.A1(net5527),
    .A2(_03198_),
    .B1(_03201_),
    .C1(_03194_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _19380_ (.A(net1638),
    .B(_03199_),
    .X(_03202_));
 sky130_fd_sc_hd__o211a_1 _19381_ (.A1(net4170),
    .A2(_03198_),
    .B1(net1133),
    .C1(_03194_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _19382_ (.A(net1537),
    .B(_03199_),
    .X(_03203_));
 sky130_fd_sc_hd__o211a_1 _19383_ (.A1(net5523),
    .A2(_03198_),
    .B1(_03203_),
    .C1(_03194_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _19384_ (.A(net1574),
    .B(_03199_),
    .X(_03204_));
 sky130_fd_sc_hd__o211a_1 _19385_ (.A1(net5487),
    .A2(_03198_),
    .B1(_03204_),
    .C1(_03194_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _19386_ (.A(net2354),
    .B(_03199_),
    .X(_03205_));
 sky130_fd_sc_hd__o211a_1 _19387_ (.A1(net5629),
    .A2(_03198_),
    .B1(_03205_),
    .C1(_03194_),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _19388_ (.A(net1115),
    .B(_03199_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_4 _19389_ (.A(_03141_),
    .X(_03207_));
 sky130_fd_sc_hd__o211a_1 _19390_ (.A1(net4194),
    .A2(_03198_),
    .B1(net1116),
    .C1(_03207_),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _19391_ (.A(net1559),
    .B(_03199_),
    .X(_03208_));
 sky130_fd_sc_hd__o211a_1 _19392_ (.A1(net5263),
    .A2(_03198_),
    .B1(_03208_),
    .C1(_03207_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _19393_ (.A(net1903),
    .B(_03199_),
    .X(_03209_));
 sky130_fd_sc_hd__o211a_1 _19394_ (.A1(net5147),
    .A2(_03198_),
    .B1(_03209_),
    .C1(_03207_),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _19395_ (.A(net1709),
    .B(_03199_),
    .X(_03210_));
 sky130_fd_sc_hd__o211a_1 _19396_ (.A1(net5398),
    .A2(_03198_),
    .B1(_03210_),
    .C1(_03207_),
    .X(_00780_));
 sky130_fd_sc_hd__clkbuf_4 _19397_ (.A(_03035_),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_4 _19398_ (.A(_03084_),
    .X(_03212_));
 sky130_fd_sc_hd__or2_1 _19399_ (.A(net1686),
    .B(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__o211a_1 _19400_ (.A1(net5435),
    .A2(_03211_),
    .B1(_03213_),
    .C1(_03207_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _19401_ (.A(net1871),
    .B(_03212_),
    .X(_03214_));
 sky130_fd_sc_hd__o211a_1 _19402_ (.A1(net5338),
    .A2(_03211_),
    .B1(_03214_),
    .C1(_03207_),
    .X(_00782_));
 sky130_fd_sc_hd__or2_1 _19403_ (.A(net1661),
    .B(_03212_),
    .X(_03215_));
 sky130_fd_sc_hd__o211a_1 _19404_ (.A1(net5346),
    .A2(_03211_),
    .B1(_03215_),
    .C1(_03207_),
    .X(_00783_));
 sky130_fd_sc_hd__or2_1 _19405_ (.A(net1964),
    .B(_03212_),
    .X(_03216_));
 sky130_fd_sc_hd__o211a_1 _19406_ (.A1(net5536),
    .A2(_03211_),
    .B1(_03216_),
    .C1(_03207_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _19407_ (.A(net2070),
    .B(_03212_),
    .X(_03217_));
 sky130_fd_sc_hd__o211a_1 _19408_ (.A1(net5605),
    .A2(_03211_),
    .B1(_03217_),
    .C1(_03207_),
    .X(_00785_));
 sky130_fd_sc_hd__or2_1 _19409_ (.A(net1689),
    .B(_03212_),
    .X(_03218_));
 sky130_fd_sc_hd__o211a_1 _19410_ (.A1(net5690),
    .A2(_03211_),
    .B1(_03218_),
    .C1(_03207_),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _19411_ (.A(net1744),
    .B(_03212_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_4 _19412_ (.A(_03141_),
    .X(_03220_));
 sky130_fd_sc_hd__o211a_1 _19413_ (.A1(net5102),
    .A2(_03211_),
    .B1(_03219_),
    .C1(_03220_),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _19414_ (.A(net647),
    .B(_03212_),
    .X(_03221_));
 sky130_fd_sc_hd__o211a_1 _19415_ (.A1(net4999),
    .A2(_03211_),
    .B1(_03221_),
    .C1(_03220_),
    .X(_00788_));
 sky130_fd_sc_hd__or2_1 _19416_ (.A(net2014),
    .B(_03212_),
    .X(_03222_));
 sky130_fd_sc_hd__o211a_1 _19417_ (.A1(net4118),
    .A2(_03211_),
    .B1(net598),
    .C1(_03220_),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _19418_ (.A(net1989),
    .B(_03212_),
    .X(_03223_));
 sky130_fd_sc_hd__o211a_1 _19419_ (.A1(net4112),
    .A2(_03211_),
    .B1(net601),
    .C1(_03220_),
    .X(_00790_));
 sky130_fd_sc_hd__clkbuf_4 _19420_ (.A(_03035_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_4 _19421_ (.A(_03084_),
    .X(_03225_));
 sky130_fd_sc_hd__or2_1 _19422_ (.A(net1718),
    .B(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__o211a_1 _19423_ (.A1(net5578),
    .A2(_03224_),
    .B1(_03226_),
    .C1(_03220_),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _19424_ (.A(net5861),
    .B(_03225_),
    .X(_03227_));
 sky130_fd_sc_hd__o211a_1 _19425_ (.A1(net2352),
    .A2(_03224_),
    .B1(net5862),
    .C1(_03220_),
    .X(_00792_));
 sky130_fd_sc_hd__or2_1 _19426_ (.A(net1543),
    .B(_03225_),
    .X(_03228_));
 sky130_fd_sc_hd__o211a_1 _19427_ (.A1(net5143),
    .A2(_03224_),
    .B1(_03228_),
    .C1(_03220_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _19428_ (.A(net1566),
    .B(_03225_),
    .X(_03229_));
 sky130_fd_sc_hd__o211a_1 _19429_ (.A1(net5018),
    .A2(_03224_),
    .B1(_03229_),
    .C1(_03220_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _19430_ (.A(net1844),
    .B(_03225_),
    .X(_03230_));
 sky130_fd_sc_hd__o211a_1 _19431_ (.A1(net5003),
    .A2(_03224_),
    .B1(_03230_),
    .C1(_03220_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _19432_ (.A(net1847),
    .B(_03225_),
    .X(_03231_));
 sky130_fd_sc_hd__o211a_1 _19433_ (.A1(net5413),
    .A2(_03224_),
    .B1(_03231_),
    .C1(_03220_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _19434_ (.A(net1631),
    .B(_03225_),
    .X(_03232_));
 sky130_fd_sc_hd__clkbuf_4 _19435_ (.A(_03141_),
    .X(_03233_));
 sky130_fd_sc_hd__o211a_1 _19436_ (.A1(net5287),
    .A2(_03224_),
    .B1(_03232_),
    .C1(_03233_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _19437_ (.A(net1862),
    .B(_03225_),
    .X(_03234_));
 sky130_fd_sc_hd__o211a_1 _19438_ (.A1(net5106),
    .A2(_03224_),
    .B1(_03234_),
    .C1(_03233_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _19439_ (.A(net2230),
    .B(_03225_),
    .X(_03235_));
 sky130_fd_sc_hd__o211a_1 _19440_ (.A1(net4979),
    .A2(_03224_),
    .B1(_03235_),
    .C1(_03233_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _19441_ (.A(net2282),
    .B(_03225_),
    .X(_03236_));
 sky130_fd_sc_hd__o211a_1 _19442_ (.A1(net5291),
    .A2(_03224_),
    .B1(_03236_),
    .C1(_03233_),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _19443_ (.A(net2873),
    .B(_03039_),
    .X(_03237_));
 sky130_fd_sc_hd__o211a_1 _19444_ (.A1(net5091),
    .A2(_03036_),
    .B1(_03237_),
    .C1(_03233_),
    .X(_00801_));
 sky130_fd_sc_hd__clkbuf_4 _19445_ (.A(_02507_),
    .X(_03238_));
 sky130_fd_sc_hd__nand2_1 _19446_ (.A(net4326),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__or3_1 _19447_ (.A(net3075),
    .B(net3151),
    .C(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__clkbuf_2 _19448_ (.A(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__mux2_1 _19449_ (.A0(net1571),
    .A1(net3254),
    .S(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__or2_1 _19450_ (.A(_03088_),
    .B(net3255),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_1 _19451_ (.A(net3256),
    .X(_00802_));
 sky130_fd_sc_hd__a31o_1 _19452_ (.A1(_02492_),
    .A2(_02498_),
    .A3(_03238_),
    .B1(net6245),
    .X(_03244_));
 sky130_fd_sc_hd__o211a_1 _19453_ (.A1(net1608),
    .A2(_03241_),
    .B1(net1596),
    .C1(_03233_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _19454_ (.A0(net3180),
    .A1(net2964),
    .S(_03241_),
    .X(_03245_));
 sky130_fd_sc_hd__or2_1 _19455_ (.A(_03088_),
    .B(net3181),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_1 _19456_ (.A(net3182),
    .X(_00804_));
 sky130_fd_sc_hd__a31o_1 _19457_ (.A1(_02492_),
    .A2(_02498_),
    .A3(_03238_),
    .B1(net6229),
    .X(_03247_));
 sky130_fd_sc_hd__o211a_1 _19458_ (.A1(_02998_),
    .A2(_03241_),
    .B1(net1532),
    .C1(_03233_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _19459_ (.A0(net3104),
    .A1(net2995),
    .S(_03241_),
    .X(_03248_));
 sky130_fd_sc_hd__or2_1 _19460_ (.A(_03088_),
    .B(net3105),
    .X(_03249_));
 sky130_fd_sc_hd__clkbuf_1 _19461_ (.A(net3106),
    .X(_00806_));
 sky130_fd_sc_hd__a31o_1 _19462_ (.A1(_02492_),
    .A2(_02498_),
    .A3(_03238_),
    .B1(net1790),
    .X(_03250_));
 sky130_fd_sc_hd__o211a_1 _19463_ (.A1(net1727),
    .A2(_03241_),
    .B1(net1791),
    .C1(_03233_),
    .X(_00807_));
 sky130_fd_sc_hd__nor2b_1 _19464_ (.A(net3075),
    .B_N(net3151),
    .Y(_03251_));
 sky130_fd_sc_hd__nand2b_1 _19465_ (.A_N(_03239_),
    .B(net3076),
    .Y(_03252_));
 sky130_fd_sc_hd__a31o_1 _19466_ (.A1(_02492_),
    .A2(_03238_),
    .A3(net3076),
    .B1(net6302),
    .X(_03253_));
 sky130_fd_sc_hd__o211a_1 _19467_ (.A1(net1572),
    .A2(net3077),
    .B1(net1535),
    .C1(_03233_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _19468_ (.A0(net1607),
    .A1(net2973),
    .S(net3077),
    .X(_03254_));
 sky130_fd_sc_hd__or2_1 _19469_ (.A(_03088_),
    .B(net3078),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_1 _19470_ (.A(net3079),
    .X(_00809_));
 sky130_fd_sc_hd__a31o_1 _19471_ (.A1(_02492_),
    .A2(_03238_),
    .A3(net3076),
    .B1(net6559),
    .X(_03256_));
 sky130_fd_sc_hd__o211a_1 _19472_ (.A1(_02996_),
    .A2(net3077),
    .B1(net1616),
    .C1(_03233_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _19473_ (.A0(net3123),
    .A1(net2951),
    .S(net3077),
    .X(_03257_));
 sky130_fd_sc_hd__or2_1 _19474_ (.A(_03088_),
    .B(net3124),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_1 _19475_ (.A(net3125),
    .X(_00811_));
 sky130_fd_sc_hd__a31o_1 _19476_ (.A1(_02492_),
    .A2(_03238_),
    .A3(net3076),
    .B1(net6524),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_4 _19477_ (.A(_03141_),
    .X(_03260_));
 sky130_fd_sc_hd__o211a_1 _19478_ (.A1(_03000_),
    .A2(net3077),
    .B1(net1541),
    .C1(_03260_),
    .X(_00812_));
 sky130_fd_sc_hd__buf_4 _19479_ (.A(_04597_),
    .X(_03261_));
 sky130_fd_sc_hd__mux2_1 _19480_ (.A0(net1726),
    .A1(net3116),
    .S(net3077),
    .X(_03262_));
 sky130_fd_sc_hd__or2_1 _19481_ (.A(_03261_),
    .B(net3117),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_1 _19482_ (.A(net3118),
    .X(_00813_));
 sky130_fd_sc_hd__or3b_1 _19483_ (.A(net3151),
    .B(_03239_),
    .C_N(net3075),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_2 _19484_ (.A(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__and3_2 _19485_ (.A(_02491_),
    .B(_02500_),
    .C(_03238_),
    .X(_03266_));
 sky130_fd_sc_hd__or2_1 _19486_ (.A(net2541),
    .B(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__o211a_1 _19487_ (.A1(net1572),
    .A2(_03265_),
    .B1(net2542),
    .C1(_03260_),
    .X(_00814_));
 sky130_fd_sc_hd__or2_1 _19488_ (.A(net5754),
    .B(_03266_),
    .X(_03268_));
 sky130_fd_sc_hd__o211a_1 _19489_ (.A1(net1608),
    .A2(_03265_),
    .B1(net5755),
    .C1(_03260_),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _19490_ (.A(net6275),
    .B(_03266_),
    .X(_03269_));
 sky130_fd_sc_hd__o211a_1 _19491_ (.A1(_02996_),
    .A2(_03265_),
    .B1(net2554),
    .C1(_03260_),
    .X(_00816_));
 sky130_fd_sc_hd__or2_1 _19492_ (.A(net6290),
    .B(_03266_),
    .X(_03270_));
 sky130_fd_sc_hd__o211a_1 _19493_ (.A1(_02998_),
    .A2(_03265_),
    .B1(net1736),
    .C1(_03260_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _19494_ (.A(net6294),
    .B(_03266_),
    .X(_03271_));
 sky130_fd_sc_hd__o211a_1 _19495_ (.A1(_03000_),
    .A2(_03265_),
    .B1(net2591),
    .C1(_03260_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _19496_ (.A(net5783),
    .B(_03266_),
    .X(_03272_));
 sky130_fd_sc_hd__o211a_1 _19497_ (.A1(net1727),
    .A2(_03265_),
    .B1(net5784),
    .C1(_03260_),
    .X(_00819_));
 sky130_fd_sc_hd__and3_1 _19498_ (.A(_02491_),
    .B(_02495_),
    .C(_03238_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_4 _19499_ (.A(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__nand3_4 _19500_ (.A(_02492_),
    .B(_02495_),
    .C(_03238_),
    .Y(_03275_));
 sky130_fd_sc_hd__or2_1 _19501_ (.A(net3112),
    .B(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__o211a_1 _19502_ (.A1(net5255),
    .A2(_03274_),
    .B1(_03276_),
    .C1(_03260_),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _19503_ (.A(net3050),
    .B(_03275_),
    .X(_03277_));
 sky130_fd_sc_hd__o211a_1 _19504_ (.A1(net5367),
    .A2(_03274_),
    .B1(_03277_),
    .C1(_03260_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _19505_ (.A(net3093),
    .B(_03275_),
    .X(_03278_));
 sky130_fd_sc_hd__o211a_1 _19506_ (.A1(net5562),
    .A2(_03274_),
    .B1(_03278_),
    .C1(_03260_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _19507_ (.A(net3096),
    .B(_03275_),
    .X(_03279_));
 sky130_fd_sc_hd__clkbuf_4 _19508_ (.A(_03141_),
    .X(_03280_));
 sky130_fd_sc_hd__o211a_1 _19509_ (.A1(net5110),
    .A2(_03274_),
    .B1(_03279_),
    .C1(_03280_),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _19510_ (.A(net614),
    .B(_03275_),
    .X(_03281_));
 sky130_fd_sc_hd__o211a_1 _19511_ (.A1(net5402),
    .A2(_03274_),
    .B1(_03281_),
    .C1(_03280_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _19512_ (.A(net1572),
    .B(_03275_),
    .X(_03282_));
 sky130_fd_sc_hd__o211a_1 _19513_ (.A1(net5459),
    .A2(_03274_),
    .B1(_03282_),
    .C1(_03280_),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _19514_ (.A(net1608),
    .B(_03275_),
    .X(_03283_));
 sky130_fd_sc_hd__o211a_1 _19515_ (.A1(net5406),
    .A2(_03274_),
    .B1(_03283_),
    .C1(_03280_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _19516_ (.A(_02996_),
    .B(_03275_),
    .X(_03284_));
 sky130_fd_sc_hd__o211a_1 _19517_ (.A1(net5124),
    .A2(_03274_),
    .B1(_03284_),
    .C1(_03280_),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _19518_ (.A(_02998_),
    .B(_03275_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _19519_ (.A1(net5045),
    .A2(_03274_),
    .B1(_03285_),
    .C1(_03280_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _19520_ (.A(_03000_),
    .B(_03275_),
    .X(_03286_));
 sky130_fd_sc_hd__o211a_1 _19521_ (.A1(net5375),
    .A2(_03274_),
    .B1(_03286_),
    .C1(_03280_),
    .X(_00829_));
 sky130_fd_sc_hd__and3_1 _19522_ (.A(_02492_),
    .B(_02497_),
    .C(_02498_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_2 _19523_ (.A(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__nand3_2 _19524_ (.A(_02492_),
    .B(_02497_),
    .C(_02498_),
    .Y(_03289_));
 sky130_fd_sc_hd__or2_1 _19525_ (.A(net1572),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__o211a_1 _19526_ (.A1(net5247),
    .A2(_03288_),
    .B1(_03290_),
    .C1(_03280_),
    .X(_00830_));
 sky130_fd_sc_hd__or2_1 _19527_ (.A(net1608),
    .B(_03289_),
    .X(_03291_));
 sky130_fd_sc_hd__o211a_1 _19528_ (.A1(net5428),
    .A2(_03288_),
    .B1(_03291_),
    .C1(_03280_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _19529_ (.A(_02996_),
    .B(_03289_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_1 _19530_ (.A1(net5547),
    .A2(_03288_),
    .B1(_03292_),
    .C1(_03280_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _19531_ (.A(_02998_),
    .B(_03289_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_4 _19532_ (.A(_08274_),
    .X(_03294_));
 sky130_fd_sc_hd__clkbuf_4 _19533_ (.A(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__o211a_1 _19534_ (.A1(net5178),
    .A2(_03288_),
    .B1(_03293_),
    .C1(_03295_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_1 _19535_ (.A(_03000_),
    .B(_03289_),
    .X(_03296_));
 sky130_fd_sc_hd__o211a_1 _19536_ (.A1(net5302),
    .A2(_03288_),
    .B1(_03296_),
    .C1(_03295_),
    .X(_00834_));
 sky130_fd_sc_hd__or2_1 _19537_ (.A(net1727),
    .B(_03289_),
    .X(_03297_));
 sky130_fd_sc_hd__o211a_1 _19538_ (.A1(net5360),
    .A2(_03288_),
    .B1(_03297_),
    .C1(_03295_),
    .X(_00835_));
 sky130_fd_sc_hd__and3_1 _19539_ (.A(_02491_),
    .B(_02497_),
    .C(net3076),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _19540_ (.A0(net3864),
    .A1(net1571),
    .S(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__and2_1 _19541_ (.A(_08279_),
    .B(net3865),
    .X(_03300_));
 sky130_fd_sc_hd__clkbuf_1 _19542_ (.A(net3866),
    .X(_00836_));
 sky130_fd_sc_hd__and3_1 _19543_ (.A(_02491_),
    .B(_02497_),
    .C(_02500_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_2 _19544_ (.A(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_4 _19545_ (.A(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__nand3_2 _19546_ (.A(_02491_),
    .B(_02497_),
    .C(_02500_),
    .Y(_03304_));
 sky130_fd_sc_hd__buf_2 _19547_ (.A(net7312),
    .X(_03305_));
 sky130_fd_sc_hd__or2_1 _19548_ (.A(net614),
    .B(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__o211a_1 _19549_ (.A1(net5132),
    .A2(_03303_),
    .B1(_03306_),
    .C1(_03295_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _19550_ (.A(net3022),
    .B(_03305_),
    .X(_03307_));
 sky130_fd_sc_hd__o211a_1 _19551_ (.A1(net5190),
    .A2(_03303_),
    .B1(_03307_),
    .C1(_03295_),
    .X(_00838_));
 sky130_fd_sc_hd__or2_1 _19552_ (.A(net3038),
    .B(_03305_),
    .X(_03308_));
 sky130_fd_sc_hd__o211a_1 _19553_ (.A1(net5155),
    .A2(_03303_),
    .B1(_03308_),
    .C1(_03295_),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _19554_ (.A(net3088),
    .B(_03305_),
    .X(_03309_));
 sky130_fd_sc_hd__o211a_1 _19555_ (.A1(net824),
    .A2(_03303_),
    .B1(_03309_),
    .C1(_03295_),
    .X(_00840_));
 sky130_fd_sc_hd__or2_1 _19556_ (.A(net3070),
    .B(_03305_),
    .X(_03310_));
 sky130_fd_sc_hd__o211a_1 _19557_ (.A1(net930),
    .A2(_03303_),
    .B1(_03310_),
    .C1(_03295_),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _19558_ (.A(net3100),
    .B(_03305_),
    .X(_03311_));
 sky130_fd_sc_hd__o211a_1 _19559_ (.A1(net5099),
    .A2(_03303_),
    .B1(_03311_),
    .C1(_03295_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _19560_ (.A(_03000_),
    .B(_03305_),
    .X(_03312_));
 sky130_fd_sc_hd__o211a_1 _19561_ (.A1(net5065),
    .A2(_03303_),
    .B1(_03312_),
    .C1(_03295_),
    .X(_00843_));
 sky130_fd_sc_hd__or2_1 _19562_ (.A(net1727),
    .B(_03305_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_4 _19563_ (.A(_03294_),
    .X(_03314_));
 sky130_fd_sc_hd__o211a_1 _19564_ (.A1(net5371),
    .A2(_03303_),
    .B1(_03313_),
    .C1(_03314_),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _19565_ (.A(net3112),
    .B(_03305_),
    .X(_03315_));
 sky130_fd_sc_hd__o211a_1 _19566_ (.A1(net5216),
    .A2(_03303_),
    .B1(_03315_),
    .C1(_03314_),
    .X(_00845_));
 sky130_fd_sc_hd__or2_1 _19567_ (.A(net3050),
    .B(_03305_),
    .X(_03316_));
 sky130_fd_sc_hd__o211a_1 _19568_ (.A1(net5014),
    .A2(_03303_),
    .B1(_03316_),
    .C1(_03314_),
    .X(_00846_));
 sky130_fd_sc_hd__or2_1 _19569_ (.A(net3093),
    .B(_03304_),
    .X(_03317_));
 sky130_fd_sc_hd__o211a_1 _19570_ (.A1(net5186),
    .A2(_03302_),
    .B1(_03317_),
    .C1(_03314_),
    .X(_00847_));
 sky130_fd_sc_hd__or2_1 _19571_ (.A(net3096),
    .B(_03304_),
    .X(_03318_));
 sky130_fd_sc_hd__o211a_1 _19572_ (.A1(net5079),
    .A2(_03302_),
    .B1(_03318_),
    .C1(_03314_),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _19573_ (.A(_02996_),
    .B(_03304_),
    .X(_03319_));
 sky130_fd_sc_hd__o211a_1 _19574_ (.A1(net5322),
    .A2(_03302_),
    .B1(_03319_),
    .C1(_03314_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_1 _19575_ (.A(_02998_),
    .B(_03304_),
    .X(_03320_));
 sky130_fd_sc_hd__o211a_1 _19576_ (.A1(net5283),
    .A2(_03302_),
    .B1(_03320_),
    .C1(_03314_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _19577_ (.A(net1572),
    .B(_03304_),
    .X(_03321_));
 sky130_fd_sc_hd__o211a_1 _19578_ (.A1(net5243),
    .A2(_03302_),
    .B1(_03321_),
    .C1(_03314_),
    .X(_00851_));
 sky130_fd_sc_hd__or2_1 _19579_ (.A(net1608),
    .B(_03304_),
    .X(_03322_));
 sky130_fd_sc_hd__o211a_1 _19580_ (.A1(net5279),
    .A2(_03302_),
    .B1(_03322_),
    .C1(_03314_),
    .X(_00852_));
 sky130_fd_sc_hd__nand2_1 _19581_ (.A(net796),
    .B(_02497_),
    .Y(_03323_));
 sky130_fd_sc_hd__nor2_1 _19582_ (.A(_02501_),
    .B(net797),
    .Y(_03324_));
 sky130_fd_sc_hd__clkbuf_4 _19583_ (.A(net798),
    .X(_03325_));
 sky130_fd_sc_hd__or2_4 _19584_ (.A(_02501_),
    .B(net797),
    .X(_03326_));
 sky130_fd_sc_hd__buf_2 _19585_ (.A(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__or2_1 _19586_ (.A(net1571),
    .B(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__o211a_1 _19587_ (.A1(net5087),
    .A2(_03325_),
    .B1(_03328_),
    .C1(_03314_),
    .X(_00853_));
 sky130_fd_sc_hd__or2_1 _19588_ (.A(net3949),
    .B(_03327_),
    .X(_03329_));
 sky130_fd_sc_hd__clkbuf_4 _19589_ (.A(_03294_),
    .X(_03330_));
 sky130_fd_sc_hd__o211a_1 _19590_ (.A1(net5072),
    .A2(_03325_),
    .B1(_03329_),
    .C1(_03330_),
    .X(_00854_));
 sky130_fd_sc_hd__or2_1 _19591_ (.A(net3957),
    .B(_03327_),
    .X(_03331_));
 sky130_fd_sc_hd__o211a_1 _19592_ (.A1(net5226),
    .A2(_03325_),
    .B1(_03331_),
    .C1(_03330_),
    .X(_00855_));
 sky130_fd_sc_hd__or2_1 _19593_ (.A(net3933),
    .B(_03327_),
    .X(_03332_));
 sky130_fd_sc_hd__o211a_1 _19594_ (.A1(net5236),
    .A2(_03325_),
    .B1(_03332_),
    .C1(_03330_),
    .X(_00856_));
 sky130_fd_sc_hd__or2_1 _19595_ (.A(net3940),
    .B(_03327_),
    .X(_03333_));
 sky130_fd_sc_hd__o211a_1 _19596_ (.A1(net5057),
    .A2(_03325_),
    .B1(_03333_),
    .C1(_03330_),
    .X(_00857_));
 sky130_fd_sc_hd__or2_1 _19597_ (.A(net1727),
    .B(_03327_),
    .X(_03334_));
 sky130_fd_sc_hd__o211a_1 _19598_ (.A1(net5318),
    .A2(_03325_),
    .B1(_03334_),
    .C1(_03330_),
    .X(_00858_));
 sky130_fd_sc_hd__or2_1 _19599_ (.A(net3112),
    .B(_03327_),
    .X(_03335_));
 sky130_fd_sc_hd__o211a_1 _19600_ (.A1(net5197),
    .A2(_03325_),
    .B1(_03335_),
    .C1(_03330_),
    .X(_00859_));
 sky130_fd_sc_hd__or2_1 _19601_ (.A(net3050),
    .B(_03327_),
    .X(_03336_));
 sky130_fd_sc_hd__o211a_1 _19602_ (.A1(net5201),
    .A2(_03325_),
    .B1(_03336_),
    .C1(_03330_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_1 _19603_ (.A(net3093),
    .B(_03327_),
    .X(_03337_));
 sky130_fd_sc_hd__o211a_1 _19604_ (.A1(net5222),
    .A2(_03325_),
    .B1(_03337_),
    .C1(_03330_),
    .X(_00861_));
 sky130_fd_sc_hd__or2_1 _19605_ (.A(net3096),
    .B(_03327_),
    .X(_03338_));
 sky130_fd_sc_hd__o211a_1 _19606_ (.A1(net5391),
    .A2(_03325_),
    .B1(_03338_),
    .C1(_03330_),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_1 _19607_ (.A(net798),
    .X(_03339_));
 sky130_fd_sc_hd__buf_2 _19608_ (.A(_03326_),
    .X(_03340_));
 sky130_fd_sc_hd__or2_1 _19609_ (.A(net614),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__o211a_1 _19610_ (.A1(net5030),
    .A2(net799),
    .B1(_03341_),
    .C1(_03330_),
    .X(_00863_));
 sky130_fd_sc_hd__or2_1 _19611_ (.A(net3022),
    .B(_03340_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_4 _19612_ (.A(_03294_),
    .X(_03343_));
 sky130_fd_sc_hd__o211a_1 _19613_ (.A1(net5121),
    .A2(net799),
    .B1(_03342_),
    .C1(_03343_),
    .X(_00864_));
 sky130_fd_sc_hd__or2_1 _19614_ (.A(net3038),
    .B(_03340_),
    .X(_03344_));
 sky130_fd_sc_hd__o211a_1 _19615_ (.A1(net969),
    .A2(net799),
    .B1(_03344_),
    .C1(_03343_),
    .X(_00865_));
 sky130_fd_sc_hd__or2_1 _19616_ (.A(net3088),
    .B(_03340_),
    .X(_03345_));
 sky130_fd_sc_hd__o211a_1 _19617_ (.A1(net4115),
    .A2(net799),
    .B1(net698),
    .C1(_03343_),
    .X(_00866_));
 sky130_fd_sc_hd__or2_1 _19618_ (.A(net910),
    .B(_03340_),
    .X(_03346_));
 sky130_fd_sc_hd__o211a_1 _19619_ (.A1(net5350),
    .A2(net799),
    .B1(net911),
    .C1(_03343_),
    .X(_00867_));
 sky130_fd_sc_hd__or2_1 _19620_ (.A(net3100),
    .B(_03340_),
    .X(_03347_));
 sky130_fd_sc_hd__o211a_1 _19621_ (.A1(net5011),
    .A2(net799),
    .B1(_03347_),
    .C1(_03343_),
    .X(_00868_));
 sky130_fd_sc_hd__or2_1 _19622_ (.A(net1591),
    .B(_03340_),
    .X(_03348_));
 sky130_fd_sc_hd__o211a_1 _19623_ (.A1(net5061),
    .A2(net799),
    .B1(_03348_),
    .C1(_03343_),
    .X(_00869_));
 sky130_fd_sc_hd__or2_1 _19624_ (.A(net3072),
    .B(_03340_),
    .X(_03349_));
 sky130_fd_sc_hd__o211a_1 _19625_ (.A1(net4991),
    .A2(net799),
    .B1(_03349_),
    .C1(_03343_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _19626_ (.A(net3109),
    .B(_03340_),
    .X(_03350_));
 sky130_fd_sc_hd__o211a_1 _19627_ (.A1(net5140),
    .A2(net799),
    .B1(_03350_),
    .C1(_03343_),
    .X(_00871_));
 sky130_fd_sc_hd__or2_1 _19628_ (.A(net642),
    .B(_03340_),
    .X(_03351_));
 sky130_fd_sc_hd__o211a_1 _19629_ (.A1(net5161),
    .A2(net799),
    .B1(_03351_),
    .C1(_03343_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _19630_ (.A(net4322),
    .B(_03326_),
    .X(_03352_));
 sky130_fd_sc_hd__o211a_1 _19631_ (.A1(net4607),
    .A2(net798),
    .B1(_03352_),
    .C1(_03343_),
    .X(_00873_));
 sky130_fd_sc_hd__or2_1 _19632_ (.A(net4401),
    .B(_03326_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_4 _19633_ (.A(_03294_),
    .X(_03354_));
 sky130_fd_sc_hd__o211a_1 _19634_ (.A1(net5034),
    .A2(net798),
    .B1(_03353_),
    .C1(_03354_),
    .X(_00874_));
 sky130_fd_sc_hd__or2_1 _19635_ (.A(net2948),
    .B(_03326_),
    .X(_03355_));
 sky130_fd_sc_hd__o211a_1 _19636_ (.A1(net5095),
    .A2(net798),
    .B1(_03355_),
    .C1(_03354_),
    .X(_00875_));
 sky130_fd_sc_hd__or2_1 _19637_ (.A(net1613),
    .B(_03326_),
    .X(_03356_));
 sky130_fd_sc_hd__o211a_1 _19638_ (.A1(net5038),
    .A2(net798),
    .B1(_03356_),
    .C1(_03354_),
    .X(_00876_));
 sky130_fd_sc_hd__nand2_1 _19639_ (.A(_02491_),
    .B(_02514_),
    .Y(_03357_));
 sky130_fd_sc_hd__or3_1 _19640_ (.A(net3075),
    .B(net3151),
    .C(net4327),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_4 _19641_ (.A(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_4 _19642_ (.A(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__and3_2 _19643_ (.A(_02491_),
    .B(_02514_),
    .C(_02498_),
    .X(_03361_));
 sky130_fd_sc_hd__buf_2 _19644_ (.A(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__or2_1 _19645_ (.A(net6300),
    .B(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__o211a_1 _19646_ (.A1(net1572),
    .A2(_03360_),
    .B1(net1704),
    .C1(_03354_),
    .X(_00877_));
 sky130_fd_sc_hd__or2_1 _19647_ (.A(net6602),
    .B(_03362_),
    .X(_03364_));
 sky130_fd_sc_hd__o211a_1 _19648_ (.A1(net1608),
    .A2(_03360_),
    .B1(net1653),
    .C1(_03354_),
    .X(_00878_));
 sky130_fd_sc_hd__or2_1 _19649_ (.A(net6854),
    .B(_03362_),
    .X(_03365_));
 sky130_fd_sc_hd__o211a_1 _19650_ (.A1(_02996_),
    .A2(_03360_),
    .B1(net2077),
    .C1(_03354_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _19651_ (.A(net6608),
    .B(_03362_),
    .X(_03366_));
 sky130_fd_sc_hd__o211a_1 _19652_ (.A1(_02998_),
    .A2(_03360_),
    .B1(net1668),
    .C1(_03354_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _19653_ (.A(net6630),
    .B(_03362_),
    .X(_03367_));
 sky130_fd_sc_hd__o211a_1 _19654_ (.A1(_03000_),
    .A2(_03360_),
    .B1(net1830),
    .C1(_03354_),
    .X(_00881_));
 sky130_fd_sc_hd__or2_1 _19655_ (.A(net6258),
    .B(_03362_),
    .X(_03368_));
 sky130_fd_sc_hd__o211a_1 _19656_ (.A1(net1727),
    .A2(_03360_),
    .B1(net1605),
    .C1(_03354_),
    .X(_00882_));
 sky130_fd_sc_hd__or2_1 _19657_ (.A(net6730),
    .B(_03362_),
    .X(_03369_));
 sky130_fd_sc_hd__o211a_1 _19658_ (.A1(net3112),
    .A2(_03360_),
    .B1(net2275),
    .C1(_03354_),
    .X(_00883_));
 sky130_fd_sc_hd__or2_1 _19659_ (.A(net6170),
    .B(_03362_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_4 _19660_ (.A(_03294_),
    .X(_03371_));
 sky130_fd_sc_hd__o211a_1 _19661_ (.A1(net6164),
    .A2(_03360_),
    .B1(net2091),
    .C1(_03371_),
    .X(_00884_));
 sky130_fd_sc_hd__or2_1 _19662_ (.A(net6180),
    .B(_03362_),
    .X(_03372_));
 sky130_fd_sc_hd__o211a_1 _19663_ (.A1(net6172),
    .A2(_03360_),
    .B1(net2257),
    .C1(_03371_),
    .X(_00885_));
 sky130_fd_sc_hd__or2_1 _19664_ (.A(net6285),
    .B(_03362_),
    .X(_03373_));
 sky130_fd_sc_hd__o211a_1 _19665_ (.A1(net3096),
    .A2(_03360_),
    .B1(net1913),
    .C1(_03371_),
    .X(_00886_));
 sky130_fd_sc_hd__clkbuf_4 _19666_ (.A(_03359_),
    .X(_03374_));
 sky130_fd_sc_hd__buf_2 _19667_ (.A(_03361_),
    .X(_03375_));
 sky130_fd_sc_hd__or2_1 _19668_ (.A(net3011),
    .B(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__o211a_1 _19669_ (.A1(net5838),
    .A2(_03374_),
    .B1(net3012),
    .C1(_03371_),
    .X(_00887_));
 sky130_fd_sc_hd__or2_1 _19670_ (.A(net6586),
    .B(_03375_),
    .X(_03377_));
 sky130_fd_sc_hd__o211a_1 _19671_ (.A1(net3022),
    .A2(_03374_),
    .B1(net1648),
    .C1(_03371_),
    .X(_00888_));
 sky130_fd_sc_hd__or2_1 _19672_ (.A(net6562),
    .B(_03375_),
    .X(_03378_));
 sky130_fd_sc_hd__o211a_1 _19673_ (.A1(net3038),
    .A2(_03374_),
    .B1(net1626),
    .C1(_03371_),
    .X(_00889_));
 sky130_fd_sc_hd__or2_1 _19674_ (.A(net6588),
    .B(_03375_),
    .X(_03379_));
 sky130_fd_sc_hd__o211a_1 _19675_ (.A1(net3088),
    .A2(_03374_),
    .B1(net1693),
    .C1(_03371_),
    .X(_00890_));
 sky130_fd_sc_hd__or2_1 _19676_ (.A(net6928),
    .B(_03375_),
    .X(_03380_));
 sky130_fd_sc_hd__o211a_1 _19677_ (.A1(net3070),
    .A2(_03374_),
    .B1(net2594),
    .C1(_03371_),
    .X(_00891_));
 sky130_fd_sc_hd__or2_1 _19678_ (.A(net7195),
    .B(_03375_),
    .X(_03381_));
 sky130_fd_sc_hd__o211a_1 _19679_ (.A1(net3100),
    .A2(_03374_),
    .B1(net2488),
    .C1(_03371_),
    .X(_00892_));
 sky130_fd_sc_hd__or2_1 _19680_ (.A(net4223),
    .B(_03375_),
    .X(_03382_));
 sky130_fd_sc_hd__o211a_1 _19681_ (.A1(net1591),
    .A2(_03374_),
    .B1(net4224),
    .C1(_03371_),
    .X(_00893_));
 sky130_fd_sc_hd__or2_1 _19682_ (.A(net1859),
    .B(_03375_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_4 _19683_ (.A(_03294_),
    .X(_03384_));
 sky130_fd_sc_hd__o211a_1 _19684_ (.A1(net6029),
    .A2(_03374_),
    .B1(net1860),
    .C1(_03384_),
    .X(_00894_));
 sky130_fd_sc_hd__or2_1 _19685_ (.A(net6622),
    .B(_03375_),
    .X(_03385_));
 sky130_fd_sc_hd__o211a_1 _19686_ (.A1(net3109),
    .A2(_03374_),
    .B1(net1730),
    .C1(_03384_),
    .X(_00895_));
 sky130_fd_sc_hd__or2_1 _19687_ (.A(net1768),
    .B(_03375_),
    .X(_03386_));
 sky130_fd_sc_hd__o211a_1 _19688_ (.A1(net6104),
    .A2(_03374_),
    .B1(net1769),
    .C1(_03384_),
    .X(_00896_));
 sky130_fd_sc_hd__or2_1 _19689_ (.A(net4672),
    .B(_03361_),
    .X(_03387_));
 sky130_fd_sc_hd__o211a_1 _19690_ (.A1(net4322),
    .A2(_03359_),
    .B1(net1701),
    .C1(_03384_),
    .X(_00897_));
 sky130_fd_sc_hd__or2_1 _19691_ (.A(net6062),
    .B(_03361_),
    .X(_03388_));
 sky130_fd_sc_hd__o211a_1 _19692_ (.A1(net4401),
    .A2(_03359_),
    .B1(net1713),
    .C1(_03384_),
    .X(_00898_));
 sky130_fd_sc_hd__or2_1 _19693_ (.A(net6071),
    .B(_03361_),
    .X(_03389_));
 sky130_fd_sc_hd__o211a_1 _19694_ (.A1(net6047),
    .A2(_03359_),
    .B1(net1671),
    .C1(_03384_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _19695_ (.A(net6043),
    .B(_03361_),
    .X(_03390_));
 sky130_fd_sc_hd__o211a_1 _19696_ (.A1(net6033),
    .A2(_03359_),
    .B1(net1549),
    .C1(_03384_),
    .X(_00900_));
 sky130_fd_sc_hd__or3b_1 _19697_ (.A(net4327),
    .B(net3075),
    .C_N(net3151),
    .X(_03391_));
 sky130_fd_sc_hd__buf_2 _19698_ (.A(net4328),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_4 _19699_ (.A(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__and3_2 _19700_ (.A(_02491_),
    .B(_02514_),
    .C(net3076),
    .X(_03394_));
 sky130_fd_sc_hd__buf_2 _19701_ (.A(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__or2_1 _19702_ (.A(net5728),
    .B(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__o211a_1 _19703_ (.A1(net1572),
    .A2(_03393_),
    .B1(net5729),
    .C1(_03384_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _19704_ (.A(net6568),
    .B(_03395_),
    .X(_03397_));
 sky130_fd_sc_hd__o211a_1 _19705_ (.A1(net1608),
    .A2(_03393_),
    .B1(net1910),
    .C1(_03384_),
    .X(_00902_));
 sky130_fd_sc_hd__or2_1 _19706_ (.A(net6682),
    .B(_03395_),
    .X(_03398_));
 sky130_fd_sc_hd__o211a_1 _19707_ (.A1(_02996_),
    .A2(_03393_),
    .B1(net1788),
    .C1(_03384_),
    .X(_00903_));
 sky130_fd_sc_hd__or2_1 _19708_ (.A(net6740),
    .B(_03395_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_4 _19709_ (.A(_03294_),
    .X(_03400_));
 sky130_fd_sc_hd__o211a_1 _19710_ (.A1(_02998_),
    .A2(_03393_),
    .B1(net1869),
    .C1(_03400_),
    .X(_00904_));
 sky130_fd_sc_hd__or2_1 _19711_ (.A(net6662),
    .B(_03395_),
    .X(_03401_));
 sky130_fd_sc_hd__o211a_1 _19712_ (.A1(_03000_),
    .A2(_03393_),
    .B1(net2114),
    .C1(_03400_),
    .X(_00905_));
 sky130_fd_sc_hd__or2_1 _19713_ (.A(net6236),
    .B(_03395_),
    .X(_03402_));
 sky130_fd_sc_hd__o211a_1 _19714_ (.A1(net1727),
    .A2(_03393_),
    .B1(net1884),
    .C1(_03400_),
    .X(_00906_));
 sky130_fd_sc_hd__or2_1 _19715_ (.A(net5792),
    .B(_03395_),
    .X(_03403_));
 sky130_fd_sc_hd__o211a_1 _19716_ (.A1(net3112),
    .A2(_03393_),
    .B1(net5793),
    .C1(_03400_),
    .X(_00907_));
 sky130_fd_sc_hd__or2_1 _19717_ (.A(net6195),
    .B(_03395_),
    .X(_03404_));
 sky130_fd_sc_hd__o211a_1 _19718_ (.A1(net6164),
    .A2(_03393_),
    .B1(net2456),
    .C1(_03400_),
    .X(_00908_));
 sky130_fd_sc_hd__or2_1 _19719_ (.A(net6202),
    .B(_03395_),
    .X(_03405_));
 sky130_fd_sc_hd__o211a_1 _19720_ (.A1(net6172),
    .A2(_03393_),
    .B1(net2534),
    .C1(_03400_),
    .X(_00909_));
 sky130_fd_sc_hd__or2_1 _19721_ (.A(net6256),
    .B(_03395_),
    .X(_03406_));
 sky130_fd_sc_hd__o211a_1 _19722_ (.A1(net3096),
    .A2(_03393_),
    .B1(net1807),
    .C1(_03400_),
    .X(_00910_));
 sky130_fd_sc_hd__clkbuf_4 _19723_ (.A(_03392_),
    .X(_03407_));
 sky130_fd_sc_hd__buf_2 _19724_ (.A(_03394_),
    .X(_03408_));
 sky130_fd_sc_hd__or2_1 _19725_ (.A(net4257),
    .B(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__o211a_1 _19726_ (.A1(net614),
    .A2(_03407_),
    .B1(net4258),
    .C1(_03400_),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _19727_ (.A(net4235),
    .B(_03408_),
    .X(_03410_));
 sky130_fd_sc_hd__o211a_1 _19728_ (.A1(net3022),
    .A2(_03407_),
    .B1(net4236),
    .C1(_03400_),
    .X(_00912_));
 sky130_fd_sc_hd__or2_1 _19729_ (.A(net5795),
    .B(_03408_),
    .X(_03411_));
 sky130_fd_sc_hd__o211a_1 _19730_ (.A1(net3038),
    .A2(_03407_),
    .B1(net5796),
    .C1(_03400_),
    .X(_00913_));
 sky130_fd_sc_hd__or2_1 _19731_ (.A(net2094),
    .B(_03408_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_4 _19732_ (.A(_03294_),
    .X(_03413_));
 sky130_fd_sc_hd__o211a_1 _19733_ (.A1(net3088),
    .A2(_03407_),
    .B1(net2095),
    .C1(_03413_),
    .X(_00914_));
 sky130_fd_sc_hd__or2_1 _19734_ (.A(net1563),
    .B(_03408_),
    .X(_03414_));
 sky130_fd_sc_hd__o211a_1 _19735_ (.A1(net3070),
    .A2(_03407_),
    .B1(net1564),
    .C1(_03413_),
    .X(_00915_));
 sky130_fd_sc_hd__or2_1 _19736_ (.A(net5718),
    .B(_03408_),
    .X(_03415_));
 sky130_fd_sc_hd__o211a_1 _19737_ (.A1(net3100),
    .A2(_03407_),
    .B1(net5719),
    .C1(_03413_),
    .X(_00916_));
 sky130_fd_sc_hd__or2_1 _19738_ (.A(net1784),
    .B(_03408_),
    .X(_03416_));
 sky130_fd_sc_hd__o211a_1 _19739_ (.A1(net6058),
    .A2(_03407_),
    .B1(net1785),
    .C1(_03413_),
    .X(_00917_));
 sky130_fd_sc_hd__or2_1 _19740_ (.A(net6066),
    .B(_03408_),
    .X(_03417_));
 sky130_fd_sc_hd__o211a_1 _19741_ (.A1(net6029),
    .A2(_03407_),
    .B1(net1645),
    .C1(_03413_),
    .X(_00918_));
 sky130_fd_sc_hd__or2_1 _19742_ (.A(net6784),
    .B(_03408_),
    .X(_03418_));
 sky130_fd_sc_hd__o211a_1 _19743_ (.A1(net3109),
    .A2(_03407_),
    .B1(net2021),
    .C1(_03413_),
    .X(_00919_));
 sky130_fd_sc_hd__or2_1 _19744_ (.A(net1638),
    .B(_03408_),
    .X(_03419_));
 sky130_fd_sc_hd__o211a_1 _19745_ (.A1(net6104),
    .A2(_03407_),
    .B1(net1639),
    .C1(_03413_),
    .X(_00920_));
 sky130_fd_sc_hd__or2_1 _19746_ (.A(net1537),
    .B(_03394_),
    .X(_03420_));
 sky130_fd_sc_hd__o211a_1 _19747_ (.A1(net4322),
    .A2(_03392_),
    .B1(net1538),
    .C1(_03413_),
    .X(_00921_));
 sky130_fd_sc_hd__or2_1 _19748_ (.A(net6055),
    .B(_03394_),
    .X(_03421_));
 sky130_fd_sc_hd__o211a_1 _19749_ (.A1(net4401),
    .A2(_03392_),
    .B1(net1575),
    .C1(_03413_),
    .X(_00922_));
 sky130_fd_sc_hd__or2_1 _19750_ (.A(net6076),
    .B(_03394_),
    .X(_03422_));
 sky130_fd_sc_hd__o211a_1 _19751_ (.A1(net6047),
    .A2(_03392_),
    .B1(net2355),
    .C1(_03413_),
    .X(_00923_));
 sky130_fd_sc_hd__or2_1 _19752_ (.A(net5762),
    .B(_03394_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_4 _19753_ (.A(_03294_),
    .X(_03424_));
 sky130_fd_sc_hd__o211a_1 _19754_ (.A1(net1613),
    .A2(_03392_),
    .B1(net5763),
    .C1(_03424_),
    .X(_00924_));
 sky130_fd_sc_hd__or3b_1 _19755_ (.A(net3151),
    .B(net4327),
    .C_N(net3075),
    .X(_03425_));
 sky130_fd_sc_hd__buf_2 _19756_ (.A(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__clkbuf_4 _19757_ (.A(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__and3_2 _19758_ (.A(_02491_),
    .B(_02500_),
    .C(_02514_),
    .X(_03428_));
 sky130_fd_sc_hd__buf_2 _19759_ (.A(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__or2_1 _19760_ (.A(net6298),
    .B(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__o211a_1 _19761_ (.A1(net1572),
    .A2(_03427_),
    .B1(net1560),
    .C1(_03424_),
    .X(_00925_));
 sky130_fd_sc_hd__or2_1 _19762_ (.A(net6624),
    .B(_03429_),
    .X(_03431_));
 sky130_fd_sc_hd__o211a_1 _19763_ (.A1(net1608),
    .A2(_03427_),
    .B1(net1904),
    .C1(_03424_),
    .X(_00926_));
 sky130_fd_sc_hd__or2_1 _19764_ (.A(net6694),
    .B(_03429_),
    .X(_03432_));
 sky130_fd_sc_hd__o211a_1 _19765_ (.A1(_02996_),
    .A2(_03427_),
    .B1(net1710),
    .C1(_03424_),
    .X(_00927_));
 sky130_fd_sc_hd__or2_1 _19766_ (.A(net6590),
    .B(_03429_),
    .X(_03433_));
 sky130_fd_sc_hd__o211a_1 _19767_ (.A1(_02998_),
    .A2(_03427_),
    .B1(net1687),
    .C1(_03424_),
    .X(_00928_));
 sky130_fd_sc_hd__or2_1 _19768_ (.A(net6720),
    .B(_03429_),
    .X(_03434_));
 sky130_fd_sc_hd__o211a_1 _19769_ (.A1(_03000_),
    .A2(_03427_),
    .B1(net1872),
    .C1(_03424_),
    .X(_00929_));
 sky130_fd_sc_hd__or2_1 _19770_ (.A(net6233),
    .B(_03429_),
    .X(_03435_));
 sky130_fd_sc_hd__o211a_1 _19771_ (.A1(net1727),
    .A2(_03427_),
    .B1(net1662),
    .C1(_03424_),
    .X(_00930_));
 sky130_fd_sc_hd__or2_1 _19772_ (.A(net6660),
    .B(_03429_),
    .X(_03436_));
 sky130_fd_sc_hd__o211a_1 _19773_ (.A1(net3112),
    .A2(_03427_),
    .B1(net1965),
    .C1(_03424_),
    .X(_00931_));
 sky130_fd_sc_hd__or2_1 _19774_ (.A(net2070),
    .B(_03429_),
    .X(_03437_));
 sky130_fd_sc_hd__o211a_1 _19775_ (.A1(net6164),
    .A2(_03427_),
    .B1(net2071),
    .C1(_03424_),
    .X(_00932_));
 sky130_fd_sc_hd__or2_1 _19776_ (.A(net1689),
    .B(_03429_),
    .X(_03438_));
 sky130_fd_sc_hd__o211a_1 _19777_ (.A1(net6172),
    .A2(_03427_),
    .B1(net1690),
    .C1(_03424_),
    .X(_00933_));
 sky130_fd_sc_hd__or2_1 _19778_ (.A(net6263),
    .B(_03429_),
    .X(_03439_));
 sky130_fd_sc_hd__buf_4 _19779_ (.A(_08274_),
    .X(_03440_));
 sky130_fd_sc_hd__buf_4 _19780_ (.A(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__o211a_1 _19781_ (.A1(net3096),
    .A2(_03427_),
    .B1(net1745),
    .C1(_03441_),
    .X(_00934_));
 sky130_fd_sc_hd__buf_4 _19782_ (.A(_03426_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_4 _19783_ (.A(_03428_),
    .X(_03443_));
 sky130_fd_sc_hd__or2_1 _19784_ (.A(net647),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__o211a_1 _19785_ (.A1(net5838),
    .A2(_03442_),
    .B1(net648),
    .C1(_03441_),
    .X(_00935_));
 sky130_fd_sc_hd__or2_1 _19786_ (.A(net2014),
    .B(_03443_),
    .X(_03445_));
 sky130_fd_sc_hd__o211a_1 _19787_ (.A1(net3022),
    .A2(_03442_),
    .B1(net2015),
    .C1(_03441_),
    .X(_00936_));
 sky130_fd_sc_hd__or2_1 _19788_ (.A(net1989),
    .B(_03443_),
    .X(_03446_));
 sky130_fd_sc_hd__o211a_1 _19789_ (.A1(net3038),
    .A2(_03442_),
    .B1(net1990),
    .C1(_03441_),
    .X(_00937_));
 sky130_fd_sc_hd__or2_1 _19790_ (.A(net6650),
    .B(_03443_),
    .X(_03447_));
 sky130_fd_sc_hd__o211a_1 _19791_ (.A1(net3088),
    .A2(_03442_),
    .B1(net1719),
    .C1(_03441_),
    .X(_00938_));
 sky130_fd_sc_hd__or2_1 _19792_ (.A(net5861),
    .B(_03443_),
    .X(_03448_));
 sky130_fd_sc_hd__o211a_1 _19793_ (.A1(net3070),
    .A2(_03442_),
    .B1(net2156),
    .C1(_03441_),
    .X(_00939_));
 sky130_fd_sc_hd__or2_1 _19794_ (.A(net6549),
    .B(_03443_),
    .X(_03449_));
 sky130_fd_sc_hd__o211a_1 _19795_ (.A1(net3100),
    .A2(_03442_),
    .B1(net1544),
    .C1(_03441_),
    .X(_00940_));
 sky130_fd_sc_hd__or2_1 _19796_ (.A(net6114),
    .B(_03443_),
    .X(_03450_));
 sky130_fd_sc_hd__o211a_1 _19797_ (.A1(net6058),
    .A2(_03442_),
    .B1(net1567),
    .C1(_03441_),
    .X(_00941_));
 sky130_fd_sc_hd__or2_1 _19798_ (.A(net6060),
    .B(_03443_),
    .X(_03451_));
 sky130_fd_sc_hd__o211a_1 _19799_ (.A1(net6029),
    .A2(_03442_),
    .B1(net1845),
    .C1(_03441_),
    .X(_00942_));
 sky130_fd_sc_hd__or2_1 _19800_ (.A(net6722),
    .B(_03443_),
    .X(_03452_));
 sky130_fd_sc_hd__o211a_1 _19801_ (.A1(net3109),
    .A2(_03442_),
    .B1(net1848),
    .C1(_03441_),
    .X(_00943_));
 sky130_fd_sc_hd__or2_1 _19802_ (.A(net6111),
    .B(_03443_),
    .X(_03453_));
 sky130_fd_sc_hd__buf_4 _19803_ (.A(_03440_),
    .X(_03454_));
 sky130_fd_sc_hd__o211a_1 _19804_ (.A1(net6104),
    .A2(_03442_),
    .B1(net1632),
    .C1(_03454_),
    .X(_00944_));
 sky130_fd_sc_hd__or2_1 _19805_ (.A(net1862),
    .B(_03428_),
    .X(_03455_));
 sky130_fd_sc_hd__o211a_1 _19806_ (.A1(net4322),
    .A2(_03426_),
    .B1(net1863),
    .C1(_03454_),
    .X(_00945_));
 sky130_fd_sc_hd__or2_1 _19807_ (.A(net6037),
    .B(_03428_),
    .X(_03456_));
 sky130_fd_sc_hd__o211a_1 _19808_ (.A1(net4401),
    .A2(_03426_),
    .B1(net2231),
    .C1(_03454_),
    .X(_00946_));
 sky130_fd_sc_hd__or2_1 _19809_ (.A(net6051),
    .B(_03428_),
    .X(_03457_));
 sky130_fd_sc_hd__o211a_1 _19810_ (.A1(net6047),
    .A2(_03426_),
    .B1(net2283),
    .C1(_03454_),
    .X(_00947_));
 sky130_fd_sc_hd__or2_1 _19811_ (.A(net2873),
    .B(_03428_),
    .X(_03458_));
 sky130_fd_sc_hd__o211a_1 _19812_ (.A1(net6033),
    .A2(_03426_),
    .B1(net2874),
    .C1(_03454_),
    .X(_00948_));
 sky130_fd_sc_hd__nand2_2 _19813_ (.A(net3971),
    .B(net2978),
    .Y(_03459_));
 sky130_fd_sc_hd__mux2_1 _19814_ (.A0(net1467),
    .A1(net3151),
    .S(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__and2_1 _19815_ (.A(_02967_),
    .B(net3152),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_1 _19816_ (.A(net3153),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _19817_ (.A0(net3151),
    .A1(net3075),
    .S(net3972),
    .X(_03462_));
 sky130_fd_sc_hd__and2_1 _19818_ (.A(_02967_),
    .B(net3973),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _19819_ (.A(net3974),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _19820_ (.A0(net3075),
    .A1(net3960),
    .S(_03459_),
    .X(_03464_));
 sky130_fd_sc_hd__and2_1 _19821_ (.A(_02967_),
    .B(net3961),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_1 _19822_ (.A(net3962),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _19823_ (.A0(net3960),
    .A1(net3925),
    .S(_03459_),
    .X(_03466_));
 sky130_fd_sc_hd__and2_1 _19824_ (.A(_02967_),
    .B(net3926),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_1 _19825_ (.A(net3927),
    .X(_00952_));
 sky130_fd_sc_hd__and2_1 _19826_ (.A(net55),
    .B(_03026_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_1 _19827_ (.A(_03468_),
    .X(_00953_));
 sky130_fd_sc_hd__and2_1 _19828_ (.A(net6322),
    .B(_03026_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _19829_ (.A(net625),
    .X(_00954_));
 sky130_fd_sc_hd__or2_2 _19830_ (.A(net41),
    .B(net40),
    .X(_03470_));
 sky130_fd_sc_hd__nand2_2 _19831_ (.A(_03034_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__and2_1 _19832_ (.A(net5467),
    .B(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__buf_2 _19833_ (.A(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__o21a_2 _19834_ (.A1(net40),
    .A2(_03473_),
    .B1(_03034_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_4 _19835_ (.A(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_4 _19836_ (.A(_03471_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_4 _19837_ (.A(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__o21ai_2 _19838_ (.A1(net40),
    .A2(_03473_),
    .B1(_03035_),
    .Y(_03478_));
 sky130_fd_sc_hd__buf_2 _19839_ (.A(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_4 _19840_ (.A(_03476_),
    .X(_03480_));
 sky130_fd_sc_hd__nor2_1 _19841_ (.A(net4335),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__a211o_1 _19842_ (.A1(net733),
    .A2(_03477_),
    .B1(_03479_),
    .C1(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__o211a_1 _19843_ (.A1(net4335),
    .A2(_03475_),
    .B1(net734),
    .C1(_03454_),
    .X(_00955_));
 sky130_fd_sc_hd__nor2_2 _19844_ (.A(net41),
    .B(net40),
    .Y(_03483_));
 sky130_fd_sc_hd__nor2_4 _19845_ (.A(_03038_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__clkbuf_4 _19846_ (.A(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__o21a_1 _19847_ (.A1(_08342_),
    .A2(_08343_),
    .B1(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__a211o_1 _19848_ (.A1(net1156),
    .A2(_03477_),
    .B1(_03479_),
    .C1(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__o211a_1 _19849_ (.A1(net4306),
    .A2(_03475_),
    .B1(net1157),
    .C1(_03454_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _19850_ (.A0(net3258),
    .A1(_08364_),
    .S(_03484_),
    .X(_03488_));
 sky130_fd_sc_hd__or2_1 _19851_ (.A(_03479_),
    .B(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__o211a_1 _19852_ (.A1(net5463),
    .A2(_03475_),
    .B1(_03489_),
    .C1(_03454_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19853_ (.A0(net3030),
    .A1(_08385_),
    .S(_03484_),
    .X(_03490_));
 sky130_fd_sc_hd__or2_1 _19854_ (.A(_03479_),
    .B(net3031),
    .X(_03491_));
 sky130_fd_sc_hd__o211a_1 _19855_ (.A1(net4338),
    .A2(_03475_),
    .B1(net3032),
    .C1(_03454_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19856_ (.A0(net6008),
    .A1(_08402_),
    .S(_03484_),
    .X(_03492_));
 sky130_fd_sc_hd__or2_1 _19857_ (.A(_03479_),
    .B(net6009),
    .X(_03493_));
 sky130_fd_sc_hd__o211a_1 _19858_ (.A1(net2935),
    .A2(_03475_),
    .B1(net6010),
    .C1(_03454_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19859_ (.A0(net2944),
    .A1(_08420_),
    .S(_03484_),
    .X(_03494_));
 sky130_fd_sc_hd__or2_1 _19860_ (.A(_03479_),
    .B(net2945),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_4 _19861_ (.A(_03440_),
    .X(_03496_));
 sky130_fd_sc_hd__o211a_1 _19862_ (.A1(net4300),
    .A2(_03475_),
    .B1(net2946),
    .C1(_03496_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _19863_ (.A0(net2927),
    .A1(_08441_),
    .S(_03484_),
    .X(_03497_));
 sky130_fd_sc_hd__or2_1 _19864_ (.A(_03478_),
    .B(net2928),
    .X(_03498_));
 sky130_fd_sc_hd__o211a_1 _19865_ (.A1(net6130),
    .A2(_03475_),
    .B1(net2929),
    .C1(_03496_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _19866_ (.A0(net2999),
    .A1(_08467_),
    .S(_03484_),
    .X(_03499_));
 sky130_fd_sc_hd__or2_1 _19867_ (.A(_03478_),
    .B(net3000),
    .X(_03500_));
 sky130_fd_sc_hd__o211a_1 _19868_ (.A1(net6199),
    .A2(_03475_),
    .B1(net3001),
    .C1(_03496_),
    .X(_00962_));
 sky130_fd_sc_hd__o221a_1 _19869_ (.A1(net1013),
    .A2(_03470_),
    .B1(_03480_),
    .B2(_08481_),
    .C1(_03475_),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_8 _19870_ (.A(_04597_),
    .X(_03502_));
 sky130_fd_sc_hd__a211o_1 _19871_ (.A1(net4219),
    .A2(_03479_),
    .B1(net1014),
    .C1(_03502_),
    .X(_00963_));
 sky130_fd_sc_hd__or2_1 _19872_ (.A(net3821),
    .B(_08479_),
    .X(_03503_));
 sky130_fd_sc_hd__nand2_1 _19873_ (.A(_03485_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21o_1 _19874_ (.A1(net3821),
    .A2(_08479_),
    .B1(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__o211a_1 _19875_ (.A1(net744),
    .A2(_03485_),
    .B1(_03474_),
    .C1(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__a211o_1 _19876_ (.A1(net6155),
    .A2(_03479_),
    .B1(net745),
    .C1(_03502_),
    .X(_00964_));
 sky130_fd_sc_hd__o21ai_1 _19877_ (.A1(net3995),
    .A2(_03503_),
    .B1(_03484_),
    .Y(_03507_));
 sky130_fd_sc_hd__o211a_1 _19878_ (.A1(net2812),
    .A2(_03485_),
    .B1(_03474_),
    .C1(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__a21oi_1 _19879_ (.A1(_03474_),
    .A2(_03504_),
    .B1(net3996),
    .Y(_03509_));
 sky130_fd_sc_hd__or3_1 _19880_ (.A(_04597_),
    .B(net2813),
    .C(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_1 _19881_ (.A(net2814),
    .X(_00965_));
 sky130_fd_sc_hd__or3_1 _19882_ (.A(net4090),
    .B(net3995),
    .C(_03503_),
    .X(_03511_));
 sky130_fd_sc_hd__o21ai_1 _19883_ (.A1(net3995),
    .A2(_03503_),
    .B1(net4090),
    .Y(_03512_));
 sky130_fd_sc_hd__a21oi_1 _19884_ (.A1(_03511_),
    .A2(_03512_),
    .B1(_03476_),
    .Y(_03513_));
 sky130_fd_sc_hd__a211o_1 _19885_ (.A1(net675),
    .A2(_03477_),
    .B1(_03479_),
    .C1(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__o211a_1 _19886_ (.A1(net6182),
    .A2(_03475_),
    .B1(net676),
    .C1(_03496_),
    .X(_00966_));
 sky130_fd_sc_hd__or2_1 _19887_ (.A(net3921),
    .B(_03511_),
    .X(_03515_));
 sky130_fd_sc_hd__inv_2 _19888_ (.A(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__a21o_1 _19889_ (.A1(net3921),
    .A2(_03511_),
    .B1(_03476_),
    .X(_03517_));
 sky130_fd_sc_hd__o221a_1 _19890_ (.A1(net3524),
    .A2(_03485_),
    .B1(_03516_),
    .B2(_03517_),
    .C1(_03474_),
    .X(_03518_));
 sky130_fd_sc_hd__buf_4 _19891_ (.A(_04597_),
    .X(_03519_));
 sky130_fd_sc_hd__a211o_1 _19892_ (.A1(net6210),
    .A2(_03479_),
    .B1(net726),
    .C1(_03519_),
    .X(_00967_));
 sky130_fd_sc_hd__nor2_1 _19893_ (.A(net3853),
    .B(_03515_),
    .Y(_03520_));
 sky130_fd_sc_hd__o21ai_1 _19894_ (.A1(_03483_),
    .A2(_03520_),
    .B1(_03474_),
    .Y(_03521_));
 sky130_fd_sc_hd__nor2_1 _19895_ (.A(net1034),
    .B(_03485_),
    .Y(_03522_));
 sky130_fd_sc_hd__a21oi_1 _19896_ (.A1(_03470_),
    .A2(_03515_),
    .B1(_03478_),
    .Y(_03523_));
 sky130_fd_sc_hd__o22a_1 _19897_ (.A1(_03521_),
    .A2(net1035),
    .B1(_03523_),
    .B2(_06226_),
    .X(_03524_));
 sky130_fd_sc_hd__nor2_1 _19898_ (.A(_03502_),
    .B(net1036),
    .Y(_00968_));
 sky130_fd_sc_hd__nor2_1 _19899_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(_03471_),
    .Y(_03525_));
 sky130_fd_sc_hd__a22o_1 _19900_ (.A1(net3156),
    .A2(_03471_),
    .B1(_03520_),
    .B2(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__a22o_1 _19901_ (.A1(net6140),
    .A2(_03521_),
    .B1(net3157),
    .B2(_03474_),
    .X(_03527_));
 sky130_fd_sc_hd__and2_1 _19902_ (.A(_08279_),
    .B(net3158),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _19903_ (.A(net3159),
    .X(_00969_));
 sky130_fd_sc_hd__o21a_2 _19904_ (.A1(net41),
    .A2(_03473_),
    .B1(_03035_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_4 _19905_ (.A(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__o21ai_2 _19906_ (.A1(net41),
    .A2(_03473_),
    .B1(_03035_),
    .Y(_03531_));
 sky130_fd_sc_hd__clkbuf_4 _19907_ (.A(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__nor2_1 _19908_ (.A(net4355),
    .B(_03480_),
    .Y(_03533_));
 sky130_fd_sc_hd__a211o_1 _19909_ (.A1(net3365),
    .A2(_03477_),
    .B1(_03532_),
    .C1(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__o211a_1 _19910_ (.A1(net4355),
    .A2(_03530_),
    .B1(net2912),
    .C1(_03496_),
    .X(_00970_));
 sky130_fd_sc_hd__nand2_1 _19911_ (.A(net2835),
    .B(_03480_),
    .Y(_03535_));
 sky130_fd_sc_hd__o211a_1 _19912_ (.A1(_08333_),
    .A2(_03480_),
    .B1(_03529_),
    .C1(net2836),
    .X(_03536_));
 sky130_fd_sc_hd__o21ai_1 _19913_ (.A1(net6082),
    .A2(_03530_),
    .B1(_08276_),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_1 _19914_ (.A(net2837),
    .B(_03537_),
    .Y(_00971_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(net3713),
    .A1(_08356_),
    .S(_03484_),
    .X(_03538_));
 sky130_fd_sc_hd__or2_1 _19916_ (.A(_03531_),
    .B(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__o211a_1 _19917_ (.A1(net4893),
    .A2(_03530_),
    .B1(_03539_),
    .C1(_03496_),
    .X(_00972_));
 sky130_fd_sc_hd__nor2_1 _19918_ (.A(_08377_),
    .B(_03480_),
    .Y(_03540_));
 sky130_fd_sc_hd__a211o_1 _19919_ (.A1(net3611),
    .A2(_03477_),
    .B1(_03532_),
    .C1(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__o211a_1 _19920_ (.A1(net6097),
    .A2(_03530_),
    .B1(net2923),
    .C1(_03496_),
    .X(_00973_));
 sky130_fd_sc_hd__nor2_1 _19921_ (.A(_08398_),
    .B(_03480_),
    .Y(_03542_));
 sky130_fd_sc_hd__a211o_1 _19922_ (.A1(net2990),
    .A2(_03477_),
    .B1(_03532_),
    .C1(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__o211a_1 _19923_ (.A1(net4294),
    .A2(_03530_),
    .B1(net2991),
    .C1(_03496_),
    .X(_00974_));
 sky130_fd_sc_hd__nor2_1 _19924_ (.A(_08414_),
    .B(_03476_),
    .Y(_03544_));
 sky130_fd_sc_hd__a211o_1 _19925_ (.A1(net3580),
    .A2(_03477_),
    .B1(_03532_),
    .C1(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__o211a_1 _19926_ (.A1(net6127),
    .A2(_03530_),
    .B1(net2890),
    .C1(_03496_),
    .X(_00975_));
 sky130_fd_sc_hd__nor2_1 _19927_ (.A(_08436_),
    .B(_03476_),
    .Y(_03546_));
 sky130_fd_sc_hd__a211o_1 _19928_ (.A1(net2956),
    .A2(_03477_),
    .B1(_03532_),
    .C1(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__o211a_1 _19929_ (.A1(net6191),
    .A2(_03530_),
    .B1(net2957),
    .C1(_03496_),
    .X(_00976_));
 sky130_fd_sc_hd__nor2_1 _19930_ (.A(_08464_),
    .B(_03476_),
    .Y(_03548_));
 sky130_fd_sc_hd__a211o_1 _19931_ (.A1(net2914),
    .A2(_03477_),
    .B1(_03532_),
    .C1(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_4 _19932_ (.A(_03440_),
    .X(_03550_));
 sky130_fd_sc_hd__o211a_1 _19933_ (.A1(net4358),
    .A2(_03530_),
    .B1(net2915),
    .C1(_03550_),
    .X(_00977_));
 sky130_fd_sc_hd__inv_2 _19934_ (.A(_08475_),
    .Y(_03551_));
 sky130_fd_sc_hd__o221a_1 _19935_ (.A1(net1018),
    .A2(_03470_),
    .B1(_03480_),
    .B2(_03551_),
    .C1(_03529_),
    .X(_03552_));
 sky130_fd_sc_hd__a211o_1 _19936_ (.A1(net4288),
    .A2(_03532_),
    .B1(net1019),
    .C1(_03519_),
    .X(_00978_));
 sky130_fd_sc_hd__or2_2 _19937_ (.A(net3917),
    .B(_08473_),
    .X(_03553_));
 sky130_fd_sc_hd__nand2_1 _19938_ (.A(net3917),
    .B(_08473_),
    .Y(_03554_));
 sky130_fd_sc_hd__a21oi_1 _19939_ (.A1(_03553_),
    .A2(_03554_),
    .B1(_03476_),
    .Y(_03555_));
 sky130_fd_sc_hd__a211o_1 _19940_ (.A1(net3360),
    .A2(_03480_),
    .B1(_03532_),
    .C1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__o211a_1 _19941_ (.A1(net6207),
    .A2(_03530_),
    .B1(net2893),
    .C1(_03550_),
    .X(_00979_));
 sky130_fd_sc_hd__or2_1 _19942_ (.A(net3286),
    .B(_03485_),
    .X(_03557_));
 sky130_fd_sc_hd__o21ai_1 _19943_ (.A1(net4675),
    .A2(_03553_),
    .B1(_03485_),
    .Y(_03558_));
 sky130_fd_sc_hd__a22o_1 _19944_ (.A1(net4675),
    .A2(_03553_),
    .B1(_03558_),
    .B2(_03529_),
    .X(_03559_));
 sky130_fd_sc_hd__a221o_1 _19945_ (.A1(net4675),
    .A2(_03532_),
    .B1(net640),
    .B2(_03559_),
    .C1(_03083_),
    .X(_00980_));
 sky130_fd_sc_hd__or3_1 _19946_ (.A(net4387),
    .B(net4675),
    .C(_03553_),
    .X(_03560_));
 sky130_fd_sc_hd__o21ai_1 _19947_ (.A1(net3880),
    .A2(_03553_),
    .B1(net4387),
    .Y(_03561_));
 sky130_fd_sc_hd__a21oi_1 _19948_ (.A1(_03560_),
    .A2(_03561_),
    .B1(_03476_),
    .Y(_03562_));
 sky130_fd_sc_hd__a211o_1 _19949_ (.A1(net668),
    .A2(_03480_),
    .B1(_03531_),
    .C1(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__o211a_1 _19950_ (.A1(net4387),
    .A2(_03530_),
    .B1(net669),
    .C1(_03550_),
    .X(_00981_));
 sky130_fd_sc_hd__or2_1 _19951_ (.A(net3893),
    .B(_03560_),
    .X(_03564_));
 sky130_fd_sc_hd__inv_2 _19952_ (.A(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a21o_1 _19953_ (.A1(net3893),
    .A2(_03560_),
    .B1(_03476_),
    .X(_03566_));
 sky130_fd_sc_hd__o221a_1 _19954_ (.A1(net747),
    .A2(_03485_),
    .B1(_03565_),
    .B2(_03566_),
    .C1(_03529_),
    .X(_03567_));
 sky130_fd_sc_hd__a211o_1 _19955_ (.A1(net6213),
    .A2(_03532_),
    .B1(net748),
    .C1(_03519_),
    .X(_00982_));
 sky130_fd_sc_hd__nor2_1 _19956_ (.A(net3279),
    .B(_03564_),
    .Y(_03568_));
 sky130_fd_sc_hd__o21ai_1 _19957_ (.A1(_03483_),
    .A2(_03568_),
    .B1(_03529_),
    .Y(_03569_));
 sky130_fd_sc_hd__nor2_1 _19958_ (.A(net3081),
    .B(_03485_),
    .Y(_03570_));
 sky130_fd_sc_hd__a21oi_1 _19959_ (.A1(_03470_),
    .A2(_03564_),
    .B1(_03531_),
    .Y(_03571_));
 sky130_fd_sc_hd__o22a_1 _19960_ (.A1(_03569_),
    .A2(net3082),
    .B1(_03571_),
    .B2(_04827_),
    .X(_03572_));
 sky130_fd_sc_hd__nor2_1 _19961_ (.A(_03502_),
    .B(net3083),
    .Y(_00983_));
 sky130_fd_sc_hd__nor2_1 _19962_ (.A(net3952),
    .B(_03471_),
    .Y(_03573_));
 sky130_fd_sc_hd__a22o_1 _19963_ (.A1(net3483),
    .A2(_03471_),
    .B1(_03568_),
    .B2(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__a22o_1 _19964_ (.A1(net3952),
    .A2(_03569_),
    .B1(_03574_),
    .B2(_03529_),
    .X(_03575_));
 sky130_fd_sc_hd__and2_1 _19965_ (.A(_08279_),
    .B(net3953),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _19966_ (.A(net3954),
    .X(_00984_));
 sky130_fd_sc_hd__nand2_4 _19967_ (.A(_03035_),
    .B(_03473_),
    .Y(_03577_));
 sky130_fd_sc_hd__clkbuf_4 _19968_ (.A(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__and3_1 _19969_ (.A(net1070),
    .B(_03034_),
    .C(_03483_),
    .X(_03579_));
 sky130_fd_sc_hd__buf_2 _19970_ (.A(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_4 _19971_ (.A(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__buf_2 _19972_ (.A(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__or2_1 _19973_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__o211a_1 _19974_ (.A1(net3695),
    .A2(_03578_),
    .B1(net4631),
    .C1(_03550_),
    .X(_00985_));
 sky130_fd_sc_hd__or2_1 _19975_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_03582_),
    .X(_03584_));
 sky130_fd_sc_hd__o211a_1 _19976_ (.A1(net3422),
    .A2(_03578_),
    .B1(net4364),
    .C1(_03550_),
    .X(_00986_));
 sky130_fd_sc_hd__or2_1 _19977_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_03582_),
    .X(_03585_));
 sky130_fd_sc_hd__o211a_1 _19978_ (.A1(net951),
    .A2(_03578_),
    .B1(net4443),
    .C1(_03550_),
    .X(_00987_));
 sky130_fd_sc_hd__or2_1 _19979_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(_03582_),
    .X(_03586_));
 sky130_fd_sc_hd__o211a_1 _19980_ (.A1(net721),
    .A2(_03578_),
    .B1(net4521),
    .C1(_03550_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _19981_ (.A0(\rbzero.debug_overlay.facingX[-5] ),
    .A1(net3519),
    .S(_03581_),
    .X(_03587_));
 sky130_fd_sc_hd__or2_1 _19982_ (.A(_03261_),
    .B(net3873),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _19983_ (.A(net3874),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _19984_ (.A0(\rbzero.debug_overlay.facingX[-4] ),
    .A1(net3775),
    .S(_03581_),
    .X(_03589_));
 sky130_fd_sc_hd__or2_1 _19985_ (.A(_03261_),
    .B(net3848),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _19986_ (.A(net3849),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _19987_ (.A0(\rbzero.debug_overlay.facingX[-3] ),
    .A1(net3139),
    .S(_03581_),
    .X(_03591_));
 sky130_fd_sc_hd__or2_1 _19988_ (.A(_03261_),
    .B(net3140),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _19989_ (.A(net3141),
    .X(_00991_));
 sky130_fd_sc_hd__or2_1 _19990_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_03582_),
    .X(_03593_));
 sky130_fd_sc_hd__o211a_1 _19991_ (.A1(net3337),
    .A2(_03578_),
    .B1(net4645),
    .C1(_03550_),
    .X(_00992_));
 sky130_fd_sc_hd__buf_4 _19992_ (.A(_03580_),
    .X(_03594_));
 sky130_fd_sc_hd__mux2_1 _19993_ (.A0(net3786),
    .A1(net3305),
    .S(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__or2_1 _19994_ (.A(_03261_),
    .B(net3787),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _19995_ (.A(net3788),
    .X(_00993_));
 sky130_fd_sc_hd__or2_1 _19996_ (.A(net4561),
    .B(_03582_),
    .X(_03597_));
 sky130_fd_sc_hd__o211a_1 _19997_ (.A1(net3301),
    .A2(_03578_),
    .B1(net4562),
    .C1(_03550_),
    .X(_00994_));
 sky130_fd_sc_hd__or2_1 _19998_ (.A(net4406),
    .B(_03582_),
    .X(_03598_));
 sky130_fd_sc_hd__o211a_1 _19999_ (.A1(net3440),
    .A2(_03578_),
    .B1(net4407),
    .C1(_03550_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _20000_ (.A0(\rbzero.debug_overlay.facingY[-9] ),
    .A1(net3756),
    .S(_03594_),
    .X(_03599_));
 sky130_fd_sc_hd__or2_1 _20001_ (.A(_03261_),
    .B(net3901),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _20002_ (.A(net3902),
    .X(_00996_));
 sky130_fd_sc_hd__or2_1 _20003_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_03582_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_4 _20004_ (.A(_03440_),
    .X(_03602_));
 sky130_fd_sc_hd__o211a_1 _20005_ (.A1(net3296),
    .A2(_03578_),
    .B1(net4515),
    .C1(_03602_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _20006_ (.A0(\rbzero.debug_overlay.facingY[-7] ),
    .A1(net3728),
    .S(_03594_),
    .X(_03603_));
 sky130_fd_sc_hd__or2_1 _20007_ (.A(_03261_),
    .B(net3830),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_1 _20008_ (.A(net3831),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _20009_ (.A0(\rbzero.debug_overlay.facingY[-6] ),
    .A1(net3743),
    .S(_03594_),
    .X(_03605_));
 sky130_fd_sc_hd__or2_1 _20010_ (.A(_03261_),
    .B(net3744),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_1 _20011_ (.A(net3745),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _20012_ (.A0(\rbzero.debug_overlay.facingY[-5] ),
    .A1(net3547),
    .S(_03594_),
    .X(_03607_));
 sky130_fd_sc_hd__or2_1 _20013_ (.A(_03261_),
    .B(net3656),
    .X(_03608_));
 sky130_fd_sc_hd__clkbuf_1 _20014_ (.A(net3657),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _20015_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_03582_),
    .X(_03609_));
 sky130_fd_sc_hd__o211a_1 _20016_ (.A1(net1098),
    .A2(_03578_),
    .B1(net4413),
    .C1(_03602_),
    .X(_01001_));
 sky130_fd_sc_hd__or2_1 _20017_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_03582_),
    .X(_03610_));
 sky130_fd_sc_hd__o211a_1 _20018_ (.A1(net888),
    .A2(_03578_),
    .B1(net4419),
    .C1(_03602_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _20019_ (.A0(\rbzero.debug_overlay.facingY[-2] ),
    .A1(net3833),
    .S(_03594_),
    .X(_03611_));
 sky130_fd_sc_hd__or2_1 _20020_ (.A(_03261_),
    .B(net3769),
    .X(_03612_));
 sky130_fd_sc_hd__clkbuf_1 _20021_ (.A(net3770),
    .X(_01003_));
 sky130_fd_sc_hd__clkbuf_4 _20022_ (.A(_03577_),
    .X(_03613_));
 sky130_fd_sc_hd__buf_2 _20023_ (.A(_03581_),
    .X(_03614_));
 sky130_fd_sc_hd__or2_1 _20024_ (.A(net4600),
    .B(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__o211a_1 _20025_ (.A1(net2887),
    .A2(_03613_),
    .B1(net4601),
    .C1(_03602_),
    .X(_01004_));
 sky130_fd_sc_hd__buf_2 _20026_ (.A(_04241_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _20027_ (.A0(net3857),
    .A1(net3764),
    .S(_03594_),
    .X(_03617_));
 sky130_fd_sc_hd__or2_1 _20028_ (.A(_03616_),
    .B(net3858),
    .X(_03618_));
 sky130_fd_sc_hd__clkbuf_1 _20029_ (.A(net3859),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _20030_ (.A0(net3876),
    .A1(net3709),
    .S(_03594_),
    .X(_03619_));
 sky130_fd_sc_hd__or2_1 _20031_ (.A(_03616_),
    .B(net3877),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _20032_ (.A(net3878),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _20033_ (.A0(net4424),
    .A1(net3543),
    .S(_03594_),
    .X(_03621_));
 sky130_fd_sc_hd__or2_1 _20034_ (.A(_03616_),
    .B(net3544),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_1 _20035_ (.A(net3545),
    .X(_01007_));
 sky130_fd_sc_hd__or2_1 _20036_ (.A(_05403_),
    .B(_03614_),
    .X(_03623_));
 sky130_fd_sc_hd__o211a_1 _20037_ (.A1(net4776),
    .A2(_03613_),
    .B1(_03623_),
    .C1(_03602_),
    .X(_01008_));
 sky130_fd_sc_hd__or2_1 _20038_ (.A(net4446),
    .B(_03614_),
    .X(_03624_));
 sky130_fd_sc_hd__o211a_1 _20039_ (.A1(net1298),
    .A2(_03613_),
    .B1(net4447),
    .C1(_03602_),
    .X(_01009_));
 sky130_fd_sc_hd__or2_1 _20040_ (.A(net4493),
    .B(_03614_),
    .X(_03625_));
 sky130_fd_sc_hd__o211a_1 _20041_ (.A1(net3388),
    .A2(_03613_),
    .B1(net4494),
    .C1(_03602_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _20042_ (.A0(net3838),
    .A1(net3453),
    .S(_03594_),
    .X(_03626_));
 sky130_fd_sc_hd__or2_1 _20043_ (.A(_03616_),
    .B(net3839),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_1 _20044_ (.A(net3840),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _20045_ (.A0(net6237),
    .A1(net3175),
    .S(_03580_),
    .X(_03628_));
 sky130_fd_sc_hd__or2_1 _20046_ (.A(_03616_),
    .B(net3176),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _20047_ (.A(net3177),
    .X(_01012_));
 sky130_fd_sc_hd__or2_1 _20048_ (.A(net4463),
    .B(_03614_),
    .X(_03630_));
 sky130_fd_sc_hd__o211a_1 _20049_ (.A1(net3323),
    .A2(_03613_),
    .B1(net4464),
    .C1(_03602_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _20050_ (.A0(net3242),
    .A1(net3229),
    .S(_03580_),
    .X(_03631_));
 sky130_fd_sc_hd__or2_1 _20051_ (.A(_03616_),
    .B(net3243),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _20052_ (.A(net3244),
    .X(_01014_));
 sky130_fd_sc_hd__or2_1 _20053_ (.A(_05401_),
    .B(_03614_),
    .X(_03633_));
 sky130_fd_sc_hd__o211a_1 _20054_ (.A1(net3449),
    .A2(_03613_),
    .B1(net4773),
    .C1(_03602_),
    .X(_01015_));
 sky130_fd_sc_hd__or2_1 _20055_ (.A(net4587),
    .B(_03614_),
    .X(_03634_));
 sky130_fd_sc_hd__o211a_1 _20056_ (.A1(net3352),
    .A2(_03613_),
    .B1(net4588),
    .C1(_03602_),
    .X(_01016_));
 sky130_fd_sc_hd__or2_1 _20057_ (.A(_02647_),
    .B(_03614_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_4 _20058_ (.A(_03440_),
    .X(_03636_));
 sky130_fd_sc_hd__o211a_1 _20059_ (.A1(net5696),
    .A2(_03613_),
    .B1(_03635_),
    .C1(_03636_),
    .X(_01017_));
 sky130_fd_sc_hd__or2_1 _20060_ (.A(net4438),
    .B(_03614_),
    .X(_03637_));
 sky130_fd_sc_hd__o211a_1 _20061_ (.A1(net4615),
    .A2(_03613_),
    .B1(_03637_),
    .C1(_03636_),
    .X(_01018_));
 sky130_fd_sc_hd__or2_1 _20062_ (.A(_05393_),
    .B(_03614_),
    .X(_03638_));
 sky130_fd_sc_hd__o211a_1 _20063_ (.A1(net4729),
    .A2(_03613_),
    .B1(_03638_),
    .C1(_03636_),
    .X(_01019_));
 sky130_fd_sc_hd__or2_1 _20064_ (.A(net4640),
    .B(_03581_),
    .X(_03639_));
 sky130_fd_sc_hd__o211a_1 _20065_ (.A1(net719),
    .A2(_03577_),
    .B1(net4641),
    .C1(_03636_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _20066_ (.A0(net4799),
    .A1(net3674),
    .S(_03580_),
    .X(_03640_));
 sky130_fd_sc_hd__or2_1 _20067_ (.A(_03616_),
    .B(net3675),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _20068_ (.A(net3676),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _20069_ (.A0(_05396_),
    .A1(net3615),
    .S(_03580_),
    .X(_03642_));
 sky130_fd_sc_hd__or2_1 _20070_ (.A(_03616_),
    .B(net3616),
    .X(_03643_));
 sky130_fd_sc_hd__clkbuf_1 _20071_ (.A(net3617),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _20072_ (.A0(net3807),
    .A1(net3189),
    .S(_03580_),
    .X(_03644_));
 sky130_fd_sc_hd__or2_1 _20073_ (.A(_03616_),
    .B(net3808),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _20074_ (.A(net3809),
    .X(_01023_));
 sky130_fd_sc_hd__or2_1 _20075_ (.A(net4459),
    .B(_03581_),
    .X(_03646_));
 sky130_fd_sc_hd__o211a_1 _20076_ (.A1(net3428),
    .A2(_03577_),
    .B1(net4460),
    .C1(_03636_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _20077_ (.A0(net3700),
    .A1(net3636),
    .S(_03580_),
    .X(_03647_));
 sky130_fd_sc_hd__or2_1 _20078_ (.A(_03616_),
    .B(net3701),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_1 _20079_ (.A(net3702),
    .X(_01025_));
 sky130_fd_sc_hd__or2_1 _20080_ (.A(_05391_),
    .B(_03581_),
    .X(_03649_));
 sky130_fd_sc_hd__o211a_1 _20081_ (.A1(net4748),
    .A2(_03577_),
    .B1(_03649_),
    .C1(_03636_),
    .X(_01026_));
 sky130_fd_sc_hd__or2_1 _20082_ (.A(net4634),
    .B(_03581_),
    .X(_03650_));
 sky130_fd_sc_hd__o211a_1 _20083_ (.A1(net3317),
    .A2(_03577_),
    .B1(net4635),
    .C1(_03636_),
    .X(_01027_));
 sky130_fd_sc_hd__or2_1 _20084_ (.A(_02864_),
    .B(_03581_),
    .X(_03651_));
 sky130_fd_sc_hd__o211a_1 _20085_ (.A1(net6020),
    .A2(_03577_),
    .B1(_03651_),
    .C1(_03636_),
    .X(_01028_));
 sky130_fd_sc_hd__nor2_1 _20086_ (.A(net3561),
    .B(_04241_),
    .Y(_03652_));
 sky130_fd_sc_hd__and2b_1 _20087_ (.A_N(net4794),
    .B(net2122),
    .X(_03653_));
 sky130_fd_sc_hd__or2_1 _20088_ (.A(net3225),
    .B(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__nand2_1 _20089_ (.A(net3225),
    .B(net4795),
    .Y(_03655_));
 sky130_fd_sc_hd__and3_1 _20090_ (.A(net3562),
    .B(net3226),
    .C(net4796),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _20091_ (.A(net3227),
    .X(_01029_));
 sky130_fd_sc_hd__inv_2 _20092_ (.A(net2628),
    .Y(_03657_));
 sky130_fd_sc_hd__nor2_1 _20093_ (.A(net2629),
    .B(net4796),
    .Y(_03658_));
 sky130_fd_sc_hd__or4b_1 _20094_ (.A(net3825),
    .B(net1601),
    .C(net2628),
    .D_N(net3328),
    .X(_03659_));
 sky130_fd_sc_hd__or4b_1 _20095_ (.A(net2937),
    .B(net4796),
    .C(_03659_),
    .D_N(net4968),
    .X(_03660_));
 sky130_fd_sc_hd__and2_1 _20096_ (.A(net3562),
    .B(net2938),
    .X(_03661_));
 sky130_fd_sc_hd__a21bo_1 _20097_ (.A1(net2629),
    .A2(net4796),
    .B1_N(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__nor2_1 _20098_ (.A(net4797),
    .B(net2630),
    .Y(_01030_));
 sky130_fd_sc_hd__a21boi_1 _20099_ (.A1(net4865),
    .A2(net4797),
    .B1_N(net3562),
    .Y(_03663_));
 sky130_fd_sc_hd__o21a_1 _20100_ (.A1(net4865),
    .A2(net4797),
    .B1(_03663_),
    .X(_01031_));
 sky130_fd_sc_hd__and3_1 _20101_ (.A(net3328),
    .B(net4865),
    .C(net4797),
    .X(_03664_));
 sky130_fd_sc_hd__a21o_1 _20102_ (.A1(net1601),
    .A2(_03658_),
    .B1(net3328),
    .X(_03665_));
 sky130_fd_sc_hd__and3b_1 _20103_ (.A_N(_03664_),
    .B(_03661_),
    .C(net3329),
    .X(_03666_));
 sky130_fd_sc_hd__clkbuf_1 _20104_ (.A(net3330),
    .X(_01032_));
 sky130_fd_sc_hd__and2_1 _20105_ (.A(net3825),
    .B(_03664_),
    .X(_03667_));
 sky130_fd_sc_hd__or2_1 _20106_ (.A(net3825),
    .B(_03664_),
    .X(_03668_));
 sky130_fd_sc_hd__and3b_1 _20107_ (.A_N(_03667_),
    .B(net3562),
    .C(net3826),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _20108_ (.A(net3827),
    .X(_01033_));
 sky130_fd_sc_hd__and3_1 _20109_ (.A(net2937),
    .B(net3825),
    .C(_03664_),
    .X(_03670_));
 sky130_fd_sc_hd__or2_1 _20110_ (.A(net2937),
    .B(_03667_),
    .X(_03671_));
 sky130_fd_sc_hd__and3b_1 _20111_ (.A_N(_03670_),
    .B(net3562),
    .C(net7330),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_1 _20112_ (.A(net3563),
    .X(_01034_));
 sky130_fd_sc_hd__o21ai_1 _20113_ (.A1(net4968),
    .A2(_03670_),
    .B1(_03661_),
    .Y(_03673_));
 sky130_fd_sc_hd__a21oi_1 _20114_ (.A1(net4968),
    .A2(_03670_),
    .B1(_03673_),
    .Y(_01035_));
 sky130_fd_sc_hd__and2b_1 _20115_ (.A_N(net4844),
    .B(net4795),
    .X(_03674_));
 sky130_fd_sc_hd__buf_4 _20116_ (.A(net4845),
    .X(_03675_));
 sky130_fd_sc_hd__buf_2 _20117_ (.A(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__or3b_1 _20118_ (.A(net3561),
    .B(net4837),
    .C_N(net2122),
    .X(_03677_));
 sky130_fd_sc_hd__clkbuf_4 _20119_ (.A(net4838),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_2 _20120_ (.A(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__or2_1 _20121_ (.A(net5598),
    .B(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__o211a_1 _20122_ (.A1(net5571),
    .A2(_03676_),
    .B1(net954),
    .C1(_03636_),
    .X(_01036_));
 sky130_fd_sc_hd__or2_1 _20123_ (.A(net5571),
    .B(_03679_),
    .X(_03681_));
 sky130_fd_sc_hd__o211a_1 _20124_ (.A1(net3641),
    .A2(_03676_),
    .B1(net5572),
    .C1(_03636_),
    .X(_01037_));
 sky130_fd_sc_hd__or2_1 _20125_ (.A(net3641),
    .B(_03679_),
    .X(_03682_));
 sky130_fd_sc_hd__clkbuf_4 _20126_ (.A(_03440_),
    .X(_03683_));
 sky130_fd_sc_hd__o211a_1 _20127_ (.A1(net3590),
    .A2(_03676_),
    .B1(_03682_),
    .C1(_03683_),
    .X(_01038_));
 sky130_fd_sc_hd__or2_1 _20128_ (.A(net3590),
    .B(_03679_),
    .X(_03684_));
 sky130_fd_sc_hd__o211a_1 _20129_ (.A1(net3817),
    .A2(_03676_),
    .B1(_03684_),
    .C1(_03683_),
    .X(_01039_));
 sky130_fd_sc_hd__or2_1 _20130_ (.A(net3817),
    .B(_03679_),
    .X(_03685_));
 sky130_fd_sc_hd__o211a_1 _20131_ (.A1(net3737),
    .A2(_03676_),
    .B1(_03685_),
    .C1(_03683_),
    .X(_01040_));
 sky130_fd_sc_hd__or2_1 _20132_ (.A(net3737),
    .B(_03679_),
    .X(_03686_));
 sky130_fd_sc_hd__o211a_1 _20133_ (.A1(net5551),
    .A2(_03676_),
    .B1(_03686_),
    .C1(_03683_),
    .X(_01041_));
 sky130_fd_sc_hd__or2_1 _20134_ (.A(net1204),
    .B(_03679_),
    .X(_03687_));
 sky130_fd_sc_hd__o211a_1 _20135_ (.A1(net5251),
    .A2(_03676_),
    .B1(_03687_),
    .C1(_03683_),
    .X(_01042_));
 sky130_fd_sc_hd__or2_1 _20136_ (.A(net5251),
    .B(_03679_),
    .X(_03688_));
 sky130_fd_sc_hd__o211a_1 _20137_ (.A1(net5410),
    .A2(_03676_),
    .B1(_03688_),
    .C1(_03683_),
    .X(_01043_));
 sky130_fd_sc_hd__or2_1 _20138_ (.A(net5410),
    .B(_03679_),
    .X(_03689_));
 sky130_fd_sc_hd__o211a_1 _20139_ (.A1(net3585),
    .A2(_03676_),
    .B1(_03689_),
    .C1(_03683_),
    .X(_01044_));
 sky130_fd_sc_hd__or2_1 _20140_ (.A(net3585),
    .B(_03679_),
    .X(_03690_));
 sky130_fd_sc_hd__o211a_1 _20141_ (.A1(net5209),
    .A2(_03676_),
    .B1(_03690_),
    .C1(_03683_),
    .X(_01045_));
 sky130_fd_sc_hd__clkbuf_4 _20142_ (.A(_03675_),
    .X(_03691_));
 sky130_fd_sc_hd__clkbuf_2 _20143_ (.A(_03678_),
    .X(_03692_));
 sky130_fd_sc_hd__or2_1 _20144_ (.A(net5209),
    .B(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__o211a_1 _20145_ (.A1(net3684),
    .A2(_03691_),
    .B1(_03693_),
    .C1(_03683_),
    .X(_01046_));
 sky130_fd_sc_hd__or2_1 _20146_ (.A(net3684),
    .B(_03692_),
    .X(_03694_));
 sky130_fd_sc_hd__o211a_1 _20147_ (.A1(net5554),
    .A2(_03691_),
    .B1(_03694_),
    .C1(_03683_),
    .X(_01047_));
 sky130_fd_sc_hd__or2_1 _20148_ (.A(net5554),
    .B(_03692_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_4 _20149_ (.A(_03440_),
    .X(_03696_));
 sky130_fd_sc_hd__o211a_1 _20150_ (.A1(net3660),
    .A2(_03691_),
    .B1(_03695_),
    .C1(_03696_),
    .X(_01048_));
 sky130_fd_sc_hd__or2_1 _20151_ (.A(net3660),
    .B(_03692_),
    .X(_03697_));
 sky130_fd_sc_hd__o211a_1 _20152_ (.A1(net3466),
    .A2(_03691_),
    .B1(_03697_),
    .C1(_03696_),
    .X(_01049_));
 sky130_fd_sc_hd__or2_1 _20153_ (.A(net3466),
    .B(_03692_),
    .X(_03698_));
 sky130_fd_sc_hd__o211a_1 _20154_ (.A1(net5566),
    .A2(_03691_),
    .B1(_03698_),
    .C1(_03696_),
    .X(_01050_));
 sky130_fd_sc_hd__or2_1 _20155_ (.A(net5566),
    .B(_03692_),
    .X(_03699_));
 sky130_fd_sc_hd__o211a_1 _20156_ (.A1(net5585),
    .A2(_03691_),
    .B1(_03699_),
    .C1(_03696_),
    .X(_01051_));
 sky130_fd_sc_hd__or2_1 _20157_ (.A(net1162),
    .B(_03692_),
    .X(_03700_));
 sky130_fd_sc_hd__o211a_1 _20158_ (.A1(net5500),
    .A2(_03691_),
    .B1(_03700_),
    .C1(_03696_),
    .X(_01052_));
 sky130_fd_sc_hd__or2_1 _20159_ (.A(net5500),
    .B(_03692_),
    .X(_03701_));
 sky130_fd_sc_hd__o211a_1 _20160_ (.A1(net5582),
    .A2(_03691_),
    .B1(_03701_),
    .C1(_03696_),
    .X(_01053_));
 sky130_fd_sc_hd__or2_1 _20161_ (.A(net1276),
    .B(_03692_),
    .X(_03702_));
 sky130_fd_sc_hd__o211a_1 _20162_ (.A1(net5540),
    .A2(_03691_),
    .B1(_03702_),
    .C1(_03696_),
    .X(_01054_));
 sky130_fd_sc_hd__or2_1 _20163_ (.A(net5540),
    .B(_03692_),
    .X(_03703_));
 sky130_fd_sc_hd__o211a_1 _20164_ (.A1(net5575),
    .A2(_03691_),
    .B1(_03703_),
    .C1(_03696_),
    .X(_01055_));
 sky130_fd_sc_hd__clkbuf_4 _20165_ (.A(_03675_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_2 _20166_ (.A(_03678_),
    .X(_03705_));
 sky130_fd_sc_hd__or2_1 _20167_ (.A(net5575),
    .B(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__o211a_1 _20168_ (.A1(net5591),
    .A2(_03704_),
    .B1(_03706_),
    .C1(_03696_),
    .X(_01056_));
 sky130_fd_sc_hd__or2_1 _20169_ (.A(net5591),
    .B(_03705_),
    .X(_03707_));
 sky130_fd_sc_hd__o211a_1 _20170_ (.A1(net3291),
    .A2(_03704_),
    .B1(_03707_),
    .C1(_03696_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_1 _20171_ (.A(net3291),
    .B(_03705_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_4 _20172_ (.A(_03440_),
    .X(_03709_));
 sky130_fd_sc_hd__o211a_1 _20173_ (.A1(net5517),
    .A2(_03704_),
    .B1(_03708_),
    .C1(_03709_),
    .X(_01058_));
 sky130_fd_sc_hd__or2_1 _20174_ (.A(net5517),
    .B(_03705_),
    .X(_03710_));
 sky130_fd_sc_hd__o211a_1 _20175_ (.A1(net5520),
    .A2(_03704_),
    .B1(_03710_),
    .C1(_03709_),
    .X(_01059_));
 sky130_fd_sc_hd__or2_1 _20176_ (.A(net5520),
    .B(_03705_),
    .X(_03711_));
 sky130_fd_sc_hd__o211a_1 _20177_ (.A1(net5544),
    .A2(_03704_),
    .B1(_03711_),
    .C1(_03709_),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _20178_ (.A(net5544),
    .B(_03705_),
    .X(_03712_));
 sky130_fd_sc_hd__o211a_1 _20179_ (.A1(net3843),
    .A2(_03704_),
    .B1(_03712_),
    .C1(_03709_),
    .X(_01061_));
 sky130_fd_sc_hd__or2_1 _20180_ (.A(net3843),
    .B(_03705_),
    .X(_03713_));
 sky130_fd_sc_hd__o211a_1 _20181_ (.A1(net5481),
    .A2(_03704_),
    .B1(_03713_),
    .C1(_03709_),
    .X(_01062_));
 sky130_fd_sc_hd__or2_1 _20182_ (.A(net5481),
    .B(_03705_),
    .X(_03714_));
 sky130_fd_sc_hd__o211a_1 _20183_ (.A1(net3557),
    .A2(_03704_),
    .B1(net5482),
    .C1(_03709_),
    .X(_01063_));
 sky130_fd_sc_hd__or2_1 _20184_ (.A(net3557),
    .B(_03705_),
    .X(_03715_));
 sky130_fd_sc_hd__o211a_1 _20185_ (.A1(net3651),
    .A2(_03704_),
    .B1(_03715_),
    .C1(_03709_),
    .X(_01064_));
 sky130_fd_sc_hd__or2_1 _20186_ (.A(net3651),
    .B(_03705_),
    .X(_03716_));
 sky130_fd_sc_hd__o211a_1 _20187_ (.A1(net5175),
    .A2(_03704_),
    .B1(_03716_),
    .C1(_03709_),
    .X(_01065_));
 sky130_fd_sc_hd__clkbuf_4 _20188_ (.A(_03675_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_2 _20189_ (.A(_03678_),
    .X(_03718_));
 sky130_fd_sc_hd__or2_1 _20190_ (.A(net5175),
    .B(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__o211a_1 _20191_ (.A1(net3782),
    .A2(_03717_),
    .B1(_03719_),
    .C1(_03709_),
    .X(_01066_));
 sky130_fd_sc_hd__or2_1 _20192_ (.A(net3782),
    .B(_03718_),
    .X(_03720_));
 sky130_fd_sc_hd__o211a_1 _20193_ (.A1(net5114),
    .A2(_03717_),
    .B1(_03720_),
    .C1(_03709_),
    .X(_01067_));
 sky130_fd_sc_hd__or2_1 _20194_ (.A(net1278),
    .B(_03718_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_4 _20195_ (.A(_03440_),
    .X(_03722_));
 sky130_fd_sc_hd__o211a_1 _20196_ (.A1(net5049),
    .A2(_03717_),
    .B1(_03721_),
    .C1(_03722_),
    .X(_01068_));
 sky130_fd_sc_hd__or2_1 _20197_ (.A(net5049),
    .B(_03718_),
    .X(_03723_));
 sky130_fd_sc_hd__o211a_1 _20198_ (.A1(net5233),
    .A2(_03717_),
    .B1(_03723_),
    .C1(_03722_),
    .X(_01069_));
 sky130_fd_sc_hd__or2_1 _20199_ (.A(net5233),
    .B(_03718_),
    .X(_03724_));
 sky130_fd_sc_hd__o211a_1 _20200_ (.A1(net5533),
    .A2(_03717_),
    .B1(_03724_),
    .C1(_03722_),
    .X(_01070_));
 sky130_fd_sc_hd__or2_1 _20201_ (.A(net5533),
    .B(_03718_),
    .X(_03725_));
 sky130_fd_sc_hd__o211a_1 _20202_ (.A1(net3412),
    .A2(_03717_),
    .B1(_03725_),
    .C1(_03722_),
    .X(_01071_));
 sky130_fd_sc_hd__or2_1 _20203_ (.A(net3412),
    .B(_03718_),
    .X(_03726_));
 sky130_fd_sc_hd__o211a_1 _20204_ (.A1(net3665),
    .A2(_03717_),
    .B1(_03726_),
    .C1(_03722_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_1 _20205_ (.A(net3665),
    .B(_03718_),
    .X(_03727_));
 sky130_fd_sc_hd__o211a_1 _20206_ (.A1(net5626),
    .A2(_03717_),
    .B1(_03727_),
    .C1(_03722_),
    .X(_01073_));
 sky130_fd_sc_hd__or2_1 _20207_ (.A(net5626),
    .B(_03718_),
    .X(_03728_));
 sky130_fd_sc_hd__o211a_1 _20208_ (.A1(net5646),
    .A2(_03717_),
    .B1(_03728_),
    .C1(_03722_),
    .X(_01074_));
 sky130_fd_sc_hd__or2_1 _20209_ (.A(net5646),
    .B(_03718_),
    .X(_03729_));
 sky130_fd_sc_hd__o211a_1 _20210_ (.A1(net3530),
    .A2(_03717_),
    .B1(_03729_),
    .C1(_03722_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_2 _20211_ (.A(_03675_),
    .X(_03730_));
 sky130_fd_sc_hd__buf_2 _20212_ (.A(_03678_),
    .X(_03731_));
 sky130_fd_sc_hd__or2_1 _20213_ (.A(net3530),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__o211a_1 _20214_ (.A1(net5439),
    .A2(_03730_),
    .B1(_03732_),
    .C1(_03722_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_1 _20215_ (.A(net1491),
    .B(_03731_),
    .X(_03733_));
 sky130_fd_sc_hd__o211a_1 _20216_ (.A1(net5387),
    .A2(_03730_),
    .B1(_03733_),
    .C1(_03722_),
    .X(_01077_));
 sky130_fd_sc_hd__or2_1 _20217_ (.A(net1318),
    .B(_03731_),
    .X(_03734_));
 sky130_fd_sc_hd__buf_2 _20218_ (.A(_08275_),
    .X(_03735_));
 sky130_fd_sc_hd__o211a_1 _20219_ (.A1(net5383),
    .A2(_03730_),
    .B1(_03734_),
    .C1(_03735_),
    .X(_01078_));
 sky130_fd_sc_hd__or2_1 _20220_ (.A(net1284),
    .B(_03731_),
    .X(_03736_));
 sky130_fd_sc_hd__o211a_1 _20221_ (.A1(net5212),
    .A2(_03730_),
    .B1(_03736_),
    .C1(_03735_),
    .X(_01079_));
 sky130_fd_sc_hd__or2_1 _20222_ (.A(net1228),
    .B(_03731_),
    .X(_03737_));
 sky130_fd_sc_hd__o211a_1 _20223_ (.A1(net5193),
    .A2(_03730_),
    .B1(_03737_),
    .C1(_03735_),
    .X(_01080_));
 sky130_fd_sc_hd__or2_1 _20224_ (.A(net5193),
    .B(_03731_),
    .X(_03738_));
 sky130_fd_sc_hd__o211a_1 _20225_ (.A1(net5240),
    .A2(_03730_),
    .B1(_03738_),
    .C1(_03735_),
    .X(_01081_));
 sky130_fd_sc_hd__or2_1 _20226_ (.A(net1270),
    .B(_03731_),
    .X(_03739_));
 sky130_fd_sc_hd__o211a_1 _20227_ (.A1(net5205),
    .A2(_03730_),
    .B1(_03739_),
    .C1(_03735_),
    .X(_01082_));
 sky130_fd_sc_hd__or2_1 _20228_ (.A(net5205),
    .B(_03731_),
    .X(_03740_));
 sky130_fd_sc_hd__o211a_1 _20229_ (.A1(net5219),
    .A2(_03730_),
    .B1(_03740_),
    .C1(_03735_),
    .X(_01083_));
 sky130_fd_sc_hd__or2_1 _20230_ (.A(net5219),
    .B(_03731_),
    .X(_03741_));
 sky130_fd_sc_hd__o211a_1 _20231_ (.A1(net3275),
    .A2(_03730_),
    .B1(_03741_),
    .C1(_03735_),
    .X(_01084_));
 sky130_fd_sc_hd__or2_1 _20232_ (.A(net3275),
    .B(_03731_),
    .X(_03742_));
 sky130_fd_sc_hd__o211a_1 _20233_ (.A1(net5432),
    .A2(_03730_),
    .B1(_03742_),
    .C1(_03735_),
    .X(_01085_));
 sky130_fd_sc_hd__clkbuf_4 _20234_ (.A(_03675_),
    .X(_03743_));
 sky130_fd_sc_hd__buf_2 _20235_ (.A(_03678_),
    .X(_03744_));
 sky130_fd_sc_hd__or2_1 _20236_ (.A(net5432),
    .B(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__o211a_1 _20237_ (.A1(net3342),
    .A2(_03743_),
    .B1(_03745_),
    .C1(_03735_),
    .X(_01086_));
 sky130_fd_sc_hd__or2_1 _20238_ (.A(net3342),
    .B(_03744_),
    .X(_03746_));
 sky130_fd_sc_hd__o211a_1 _20239_ (.A1(net3435),
    .A2(_03743_),
    .B1(_03746_),
    .C1(_03735_),
    .X(_01087_));
 sky130_fd_sc_hd__or2_1 _20240_ (.A(net3435),
    .B(_03744_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_4 _20241_ (.A(_08275_),
    .X(_03748_));
 sky130_fd_sc_hd__o211a_1 _20242_ (.A1(net3800),
    .A2(_03743_),
    .B1(_03747_),
    .C1(_03748_),
    .X(_01088_));
 sky130_fd_sc_hd__or2_1 _20243_ (.A(net3800),
    .B(_03744_),
    .X(_03749_));
 sky130_fd_sc_hd__o211a_1 _20244_ (.A1(net5623),
    .A2(_03743_),
    .B1(_03749_),
    .C1(_03748_),
    .X(_01089_));
 sky130_fd_sc_hd__or2_1 _20245_ (.A(net5623),
    .B(_03744_),
    .X(_03750_));
 sky130_fd_sc_hd__o211a_1 _20246_ (.A1(net5665),
    .A2(_03743_),
    .B1(_03750_),
    .C1(_03748_),
    .X(_01090_));
 sky130_fd_sc_hd__or2_1 _20247_ (.A(net5665),
    .B(_03744_),
    .X(_03751_));
 sky130_fd_sc_hd__o211a_1 _20248_ (.A1(net3598),
    .A2(_03743_),
    .B1(_03751_),
    .C1(_03748_),
    .X(_01091_));
 sky130_fd_sc_hd__or2_1 _20249_ (.A(net3598),
    .B(_03744_),
    .X(_03752_));
 sky130_fd_sc_hd__o211a_1 _20250_ (.A1(net3646),
    .A2(_03743_),
    .B1(_03752_),
    .C1(_03748_),
    .X(_01092_));
 sky130_fd_sc_hd__or2_1 _20251_ (.A(net3646),
    .B(_03744_),
    .X(_03753_));
 sky130_fd_sc_hd__o211a_1 _20252_ (.A1(net3568),
    .A2(_03743_),
    .B1(_03753_),
    .C1(_03748_),
    .X(_01093_));
 sky130_fd_sc_hd__or2_1 _20253_ (.A(net3568),
    .B(_03744_),
    .X(_03754_));
 sky130_fd_sc_hd__o211a_1 _20254_ (.A1(net5588),
    .A2(_03743_),
    .B1(_03754_),
    .C1(_03748_),
    .X(_01094_));
 sky130_fd_sc_hd__or2_1 _20255_ (.A(net5588),
    .B(_03744_),
    .X(_03755_));
 sky130_fd_sc_hd__o211a_1 _20256_ (.A1(net3488),
    .A2(_03743_),
    .B1(_03755_),
    .C1(_03748_),
    .X(_01095_));
 sky130_fd_sc_hd__clkbuf_4 _20257_ (.A(net4845),
    .X(_03756_));
 sky130_fd_sc_hd__buf_1 _20258_ (.A(net4838),
    .X(_03757_));
 sky130_fd_sc_hd__or2_1 _20259_ (.A(net3488),
    .B(net4839),
    .X(_03758_));
 sky130_fd_sc_hd__o211a_1 _20260_ (.A1(net3476),
    .A2(_03756_),
    .B1(_03758_),
    .C1(_03748_),
    .X(_01096_));
 sky130_fd_sc_hd__or2_1 _20261_ (.A(net3476),
    .B(net4839),
    .X(_03759_));
 sky130_fd_sc_hd__o211a_1 _20262_ (.A1(net4850),
    .A2(_03756_),
    .B1(_03759_),
    .C1(_03748_),
    .X(_01097_));
 sky130_fd_sc_hd__or2_1 _20263_ (.A(net4850),
    .B(net4839),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_4 _20264_ (.A(_08275_),
    .X(_03761_));
 sky130_fd_sc_hd__o211a_1 _20265_ (.A1(net3705),
    .A2(_03756_),
    .B1(net4851),
    .C1(_03761_),
    .X(_01098_));
 sky130_fd_sc_hd__or2_1 _20266_ (.A(net3705),
    .B(_03757_),
    .X(_03762_));
 sky130_fd_sc_hd__o211a_1 _20267_ (.A1(net4833),
    .A2(_03756_),
    .B1(_03762_),
    .C1(_03761_),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _20268_ (.A(net4833),
    .B(net4839),
    .X(_03763_));
 sky130_fd_sc_hd__o211a_1 _20269_ (.A1(net3812),
    .A2(_03756_),
    .B1(_03763_),
    .C1(_03761_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _20270_ (.A(net3812),
    .B(net4839),
    .X(_03764_));
 sky130_fd_sc_hd__o211a_1 _20271_ (.A1(net3752),
    .A2(_03756_),
    .B1(net4840),
    .C1(_03761_),
    .X(_01101_));
 sky130_fd_sc_hd__or2_1 _20272_ (.A(net3752),
    .B(net4839),
    .X(_03765_));
 sky130_fd_sc_hd__o211a_1 _20273_ (.A1(net3670),
    .A2(_03756_),
    .B1(_03765_),
    .C1(_03761_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _20274_ (.A(net3670),
    .B(net4839),
    .X(_03766_));
 sky130_fd_sc_hd__o211a_1 _20275_ (.A1(net3679),
    .A2(_03756_),
    .B1(_03766_),
    .C1(_03761_),
    .X(_01103_));
 sky130_fd_sc_hd__or2_1 _20276_ (.A(net3679),
    .B(net4839),
    .X(_03767_));
 sky130_fd_sc_hd__o211a_1 _20277_ (.A1(net3514),
    .A2(_03756_),
    .B1(_03767_),
    .C1(_03761_),
    .X(_01104_));
 sky130_fd_sc_hd__or2_1 _20278_ (.A(net3514),
    .B(net4839),
    .X(_03768_));
 sky130_fd_sc_hd__o211a_1 _20279_ (.A1(net3496),
    .A2(_03756_),
    .B1(_03768_),
    .C1(_03761_),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _20280_ (.A(net3496),
    .B(_03678_),
    .X(_03769_));
 sky130_fd_sc_hd__o211a_1 _20281_ (.A1(net3383),
    .A2(_03675_),
    .B1(_03769_),
    .C1(_03761_),
    .X(_01106_));
 sky130_fd_sc_hd__or2_1 _20282_ (.A(net3383),
    .B(_03678_),
    .X(_03770_));
 sky130_fd_sc_hd__o211a_1 _20283_ (.A1(net4881),
    .A2(_03675_),
    .B1(_03770_),
    .C1(_03761_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _20284_ (.A(net1302),
    .B(_03678_),
    .X(_03771_));
 sky130_fd_sc_hd__o211a_1 _20285_ (.A1(net4868),
    .A2(_03675_),
    .B1(_03771_),
    .C1(_08276_),
    .X(_01108_));
 sky130_fd_sc_hd__or2_1 _20286_ (.A(net1508),
    .B(_03678_),
    .X(_03772_));
 sky130_fd_sc_hd__o211a_1 _20287_ (.A1(net4861),
    .A2(_03675_),
    .B1(_03772_),
    .C1(_08276_),
    .X(_01109_));
 sky130_fd_sc_hd__buf_1 _20288_ (.A(clknet_1_0__leaf__04800_),
    .X(_03773_));
 sky130_fd_sc_hd__buf_1 _20289_ (.A(clknet_1_0__leaf__03773_),
    .X(_03774_));
 sky130_fd_sc_hd__inv_2 _20290__27 (.A(clknet_1_1__leaf__03774_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _20291__28 (.A(clknet_1_1__leaf__03774_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _20292__29 (.A(clknet_1_1__leaf__03774_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _20293__30 (.A(clknet_1_1__leaf__03774_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _20294__31 (.A(clknet_1_1__leaf__03774_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _20295__32 (.A(clknet_1_1__leaf__03774_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _20296__33 (.A(clknet_1_0__leaf__03774_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _20297__34 (.A(clknet_1_0__leaf__03774_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _20298__35 (.A(clknet_1_0__leaf__03774_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _20299__36 (.A(clknet_1_0__leaf__03774_),
    .Y(net175));
 sky130_fd_sc_hd__buf_1 _20300_ (.A(clknet_1_1__leaf__03773_),
    .X(_03775_));
 sky130_fd_sc_hd__inv_2 _20301__37 (.A(clknet_1_1__leaf__03775_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _20302__38 (.A(clknet_1_1__leaf__03775_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _20303__39 (.A(clknet_1_1__leaf__03775_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _20304__40 (.A(clknet_1_1__leaf__03775_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _20305__41 (.A(clknet_1_0__leaf__03775_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _20306__42 (.A(clknet_1_0__leaf__03775_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _20307__43 (.A(clknet_1_0__leaf__03775_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _20308__44 (.A(clknet_1_0__leaf__03775_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _20309__45 (.A(clknet_1_0__leaf__03775_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _20310__46 (.A(clknet_1_0__leaf__03775_),
    .Y(net185));
 sky130_fd_sc_hd__buf_1 _20311_ (.A(clknet_1_1__leaf__03773_),
    .X(_03776_));
 sky130_fd_sc_hd__inv_2 _20312__47 (.A(clknet_1_0__leaf__03776_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _20313__48 (.A(clknet_1_0__leaf__03776_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _20314__49 (.A(clknet_1_0__leaf__03776_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _20315__50 (.A(clknet_1_0__leaf__03776_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _20316__51 (.A(clknet_1_0__leaf__03776_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _20317__52 (.A(clknet_1_0__leaf__03776_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _20318__53 (.A(clknet_1_1__leaf__03776_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _20319__54 (.A(clknet_1_1__leaf__03776_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _20320__55 (.A(clknet_1_1__leaf__03776_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _20321__56 (.A(clknet_1_1__leaf__03776_),
    .Y(net195));
 sky130_fd_sc_hd__buf_1 _20322_ (.A(clknet_1_1__leaf__03773_),
    .X(_03777_));
 sky130_fd_sc_hd__inv_2 _20323__57 (.A(clknet_1_0__leaf__03777_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _20324__58 (.A(clknet_1_0__leaf__03777_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _20325__59 (.A(clknet_1_0__leaf__03777_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _20326__60 (.A(clknet_1_0__leaf__03777_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _20327__61 (.A(clknet_1_0__leaf__03777_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _20328__62 (.A(clknet_1_1__leaf__03777_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _20329__63 (.A(clknet_1_1__leaf__03777_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _20330__64 (.A(clknet_1_1__leaf__03777_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _20331__65 (.A(clknet_1_1__leaf__03777_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _20332__66 (.A(clknet_1_1__leaf__03777_),
    .Y(net205));
 sky130_fd_sc_hd__buf_1 _20333_ (.A(clknet_1_1__leaf__03773_),
    .X(_03778_));
 sky130_fd_sc_hd__inv_2 _20334__67 (.A(clknet_1_1__leaf__03778_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _20335__68 (.A(clknet_1_1__leaf__03778_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _20336__69 (.A(clknet_1_1__leaf__03778_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _20337__70 (.A(clknet_1_1__leaf__03778_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _20338__71 (.A(clknet_1_1__leaf__03778_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _20339__72 (.A(clknet_1_1__leaf__03778_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _20340__73 (.A(clknet_1_0__leaf__03778_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _20341__74 (.A(clknet_1_0__leaf__03778_),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _20342__75 (.A(clknet_1_0__leaf__03778_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _20343__76 (.A(clknet_1_0__leaf__03778_),
    .Y(net215));
 sky130_fd_sc_hd__buf_1 _20344_ (.A(clknet_1_1__leaf__03773_),
    .X(_03779_));
 sky130_fd_sc_hd__inv_2 _20345__77 (.A(clknet_1_1__leaf__03779_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _20346__78 (.A(clknet_1_1__leaf__03779_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _20347__79 (.A(clknet_1_1__leaf__03779_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _20348__80 (.A(clknet_1_1__leaf__03779_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _20349__81 (.A(clknet_1_1__leaf__03779_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _20350__82 (.A(clknet_1_0__leaf__03779_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _20351__83 (.A(clknet_1_0__leaf__03779_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _20352__84 (.A(clknet_1_0__leaf__03779_),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _20353__85 (.A(clknet_1_0__leaf__03779_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _20354__86 (.A(clknet_1_0__leaf__03779_),
    .Y(net225));
 sky130_fd_sc_hd__buf_1 _20355_ (.A(clknet_1_0__leaf__04800_),
    .X(_03780_));
 sky130_fd_sc_hd__buf_1 _20356_ (.A(clknet_1_1__leaf__03780_),
    .X(_03781_));
 sky130_fd_sc_hd__inv_2 _20357__87 (.A(clknet_1_0__leaf__03781_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _20358__88 (.A(clknet_1_0__leaf__03781_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _20359__89 (.A(clknet_1_0__leaf__03781_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _20360__90 (.A(clknet_1_0__leaf__03781_),
    .Y(net229));
 sky130_fd_sc_hd__buf_4 _20361_ (.A(net6176),
    .X(_03782_));
 sky130_fd_sc_hd__o211a_1 _20362_ (.A1(_03782_),
    .A2(net5467),
    .B1(_08276_),
    .C1(_03477_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _20363_ (.A0(net1587),
    .A1(net3268),
    .S(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__and2_1 _20364_ (.A(_08279_),
    .B(net3269),
    .X(_03784_));
 sky130_fd_sc_hd__clkbuf_1 _20365_ (.A(net3270),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _20366_ (.A0(net1623),
    .A1(net3641),
    .S(_03782_),
    .X(_03785_));
 sky130_fd_sc_hd__and2_1 _20367_ (.A(_08279_),
    .B(net3642),
    .X(_03786_));
 sky130_fd_sc_hd__clkbuf_1 _20368_ (.A(net3643),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _20369_ (.A0(net719),
    .A1(net3590),
    .S(_03782_),
    .X(_03787_));
 sky130_fd_sc_hd__and2_1 _20370_ (.A(_08279_),
    .B(net3591),
    .X(_03788_));
 sky130_fd_sc_hd__clkbuf_1 _20371_ (.A(net3592),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _20372_ (.A0(net3674),
    .A1(net3817),
    .S(_03782_),
    .X(_03789_));
 sky130_fd_sc_hd__and2_1 _20373_ (.A(_08279_),
    .B(net3818),
    .X(_03790_));
 sky130_fd_sc_hd__clkbuf_1 _20374_ (.A(net3819),
    .X(_01178_));
 sky130_fd_sc_hd__buf_2 _20375_ (.A(_08275_),
    .X(_03791_));
 sky130_fd_sc_hd__mux2_1 _20376_ (.A0(net3615),
    .A1(net3737),
    .S(_03782_),
    .X(_03792_));
 sky130_fd_sc_hd__and2_1 _20377_ (.A(_03791_),
    .B(net3738),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_1 _20378_ (.A(net3739),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _20379_ (.A0(net3189),
    .A1(net1204),
    .S(_03782_),
    .X(_03794_));
 sky130_fd_sc_hd__and2_1 _20380_ (.A(_03791_),
    .B(net3190),
    .X(_03795_));
 sky130_fd_sc_hd__clkbuf_1 _20381_ (.A(net3191),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _20382_ (.A0(net3428),
    .A1(net1232),
    .S(_03782_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _20383_ (.A(_03791_),
    .B(net3429),
    .X(_03797_));
 sky130_fd_sc_hd__clkbuf_1 _20384_ (.A(net3430),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _20385_ (.A0(net3636),
    .A1(net1222),
    .S(_03782_),
    .X(_03798_));
 sky130_fd_sc_hd__and2_1 _20386_ (.A(_03791_),
    .B(net3637),
    .X(_03799_));
 sky130_fd_sc_hd__clkbuf_1 _20387_ (.A(net3638),
    .X(_01182_));
 sky130_fd_sc_hd__buf_1 _20388_ (.A(net3249),
    .X(_03800_));
 sky130_fd_sc_hd__buf_4 _20389_ (.A(net3250),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _20390_ (.A0(net1598),
    .A1(net3585),
    .S(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_1 _20391_ (.A(_03791_),
    .B(net3586),
    .X(_03803_));
 sky130_fd_sc_hd__clkbuf_1 _20392_ (.A(net3587),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _20393_ (.A0(net3317),
    .A1(net1245),
    .S(_03801_),
    .X(_03804_));
 sky130_fd_sc_hd__and2_1 _20394_ (.A(_03791_),
    .B(net3318),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _20395_ (.A(net3319),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _20396_ (.A0(net2900),
    .A1(net3684),
    .S(_03801_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_1 _20397_ (.A(_03791_),
    .B(net3685),
    .X(_03807_));
 sky130_fd_sc_hd__clkbuf_1 _20398_ (.A(net3686),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _20399_ (.A0(net3606),
    .A1(net1286),
    .S(_03801_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_1 _20400_ (.A(_03791_),
    .B(net3607),
    .X(_03809_));
 sky130_fd_sc_hd__clkbuf_1 _20401_ (.A(net3608),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _20402_ (.A0(net2833),
    .A1(net3660),
    .S(_03801_),
    .X(_03810_));
 sky130_fd_sc_hd__and2_1 _20403_ (.A(_03791_),
    .B(net3661),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _20404_ (.A(net3662),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _20405_ (.A0(net1298),
    .A1(net3466),
    .S(_03801_),
    .X(_03812_));
 sky130_fd_sc_hd__and2_1 _20406_ (.A(_03791_),
    .B(net3467),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _20407_ (.A(net3468),
    .X(_01188_));
 sky130_fd_sc_hd__buf_2 _20408_ (.A(_08275_),
    .X(_03814_));
 sky130_fd_sc_hd__mux2_1 _20409_ (.A0(net3388),
    .A1(net1168),
    .S(_03801_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _20410_ (.A(_03814_),
    .B(net3389),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _20411_ (.A(net3390),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _20412_ (.A0(net3453),
    .A1(net1162),
    .S(_03801_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_1 _20413_ (.A(_03814_),
    .B(net3454),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _20414_ (.A(net3455),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _20415_ (.A0(net3347),
    .A1(net1105),
    .S(_03801_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _20416_ (.A(_03814_),
    .B(net3348),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _20417_ (.A(net3349),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _20418_ (.A0(net3323),
    .A1(net1276),
    .S(_03801_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_1 _20419_ (.A(_03814_),
    .B(net3324),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _20420_ (.A(net3325),
    .X(_01192_));
 sky130_fd_sc_hd__clkbuf_4 _20421_ (.A(net3250),
    .X(_03823_));
 sky130_fd_sc_hd__mux2_1 _20422_ (.A0(net3229),
    .A1(net1294),
    .S(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_1 _20423_ (.A(_03814_),
    .B(net3230),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_1 _20424_ (.A(net3231),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _20425_ (.A0(net3449),
    .A1(net1389),
    .S(_03823_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_1 _20426_ (.A(_03814_),
    .B(net3450),
    .X(_03827_));
 sky130_fd_sc_hd__clkbuf_1 _20427_ (.A(net3451),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _20428_ (.A0(net3352),
    .A1(net1280),
    .S(_03823_),
    .X(_03828_));
 sky130_fd_sc_hd__and2_1 _20429_ (.A(_03814_),
    .B(net3353),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _20430_ (.A(net3354),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _20431_ (.A0(net1440),
    .A1(net3291),
    .S(_03823_),
    .X(_03830_));
 sky130_fd_sc_hd__and2_1 _20432_ (.A(_03814_),
    .B(net3292),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _20433_ (.A(net3293),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _20434_ (.A0(net3756),
    .A1(net1288),
    .S(_03823_),
    .X(_03832_));
 sky130_fd_sc_hd__and2_1 _20435_ (.A(_03814_),
    .B(net3757),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _20436_ (.A(net3758),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _20437_ (.A0(net3296),
    .A1(net1263),
    .S(_03823_),
    .X(_03834_));
 sky130_fd_sc_hd__and2_1 _20438_ (.A(_03814_),
    .B(net3297),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_1 _20439_ (.A(net3298),
    .X(_01198_));
 sky130_fd_sc_hd__clkbuf_2 _20440_ (.A(_08275_),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_1 _20441_ (.A0(net3728),
    .A1(net1292),
    .S(_03823_),
    .X(_03837_));
 sky130_fd_sc_hd__and2_1 _20442_ (.A(_03836_),
    .B(net3729),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_1 _20443_ (.A(net3730),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _20444_ (.A0(net3743),
    .A1(net3843),
    .S(_03823_),
    .X(_03839_));
 sky130_fd_sc_hd__and2_1 _20445_ (.A(_03836_),
    .B(net3844),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_1 _20446_ (.A(net3845),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _20447_ (.A0(net3547),
    .A1(net1335),
    .S(_03823_),
    .X(_03841_));
 sky130_fd_sc_hd__and2_1 _20448_ (.A(_03836_),
    .B(net3548),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_1 _20449_ (.A(net3549),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _20450_ (.A0(net1098),
    .A1(net3557),
    .S(_03823_),
    .X(_03843_));
 sky130_fd_sc_hd__and2_1 _20451_ (.A(_03836_),
    .B(net3558),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_1 _20452_ (.A(net3559),
    .X(_01202_));
 sky130_fd_sc_hd__clkbuf_4 _20453_ (.A(net3250),
    .X(_03845_));
 sky130_fd_sc_hd__mux2_1 _20454_ (.A0(net888),
    .A1(net3651),
    .S(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__and2_1 _20455_ (.A(_03836_),
    .B(net3652),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_1 _20456_ (.A(net3653),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _20457_ (.A0(net3833),
    .A1(net1470),
    .S(_03845_),
    .X(_03848_));
 sky130_fd_sc_hd__and2_1 _20458_ (.A(_03836_),
    .B(net3834),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_1 _20459_ (.A(net3835),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _20460_ (.A0(net2887),
    .A1(net3782),
    .S(_03845_),
    .X(_03850_));
 sky130_fd_sc_hd__and2_1 _20461_ (.A(_03836_),
    .B(net3783),
    .X(_03851_));
 sky130_fd_sc_hd__clkbuf_1 _20462_ (.A(net3784),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _20463_ (.A0(net3764),
    .A1(net1278),
    .S(_03845_),
    .X(_03852_));
 sky130_fd_sc_hd__and2_1 _20464_ (.A(_03836_),
    .B(net3765),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_1 _20465_ (.A(net3766),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _20466_ (.A0(net3709),
    .A1(net1274),
    .S(_03845_),
    .X(_03854_));
 sky130_fd_sc_hd__and2_1 _20467_ (.A(_03836_),
    .B(net3710),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_1 _20468_ (.A(net3711),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _20469_ (.A0(net3695),
    .A1(net1433),
    .S(_03845_),
    .X(_03856_));
 sky130_fd_sc_hd__and2_1 _20470_ (.A(_03836_),
    .B(net3696),
    .X(_03857_));
 sky130_fd_sc_hd__clkbuf_1 _20471_ (.A(net3697),
    .X(_01208_));
 sky130_fd_sc_hd__buf_2 _20472_ (.A(_08275_),
    .X(_03858_));
 sky130_fd_sc_hd__mux2_1 _20473_ (.A0(net3422),
    .A1(net1510),
    .S(_03845_),
    .X(_03859_));
 sky130_fd_sc_hd__and2_1 _20474_ (.A(_03858_),
    .B(net3423),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_1 _20475_ (.A(net3424),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _20476_ (.A0(net951),
    .A1(net3412),
    .S(_03845_),
    .X(_03861_));
 sky130_fd_sc_hd__and2_1 _20477_ (.A(_03858_),
    .B(net3413),
    .X(_03862_));
 sky130_fd_sc_hd__clkbuf_1 _20478_ (.A(net3414),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _20479_ (.A0(net721),
    .A1(net3665),
    .S(_03845_),
    .X(_03863_));
 sky130_fd_sc_hd__and2_1 _20480_ (.A(_03858_),
    .B(net3666),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_1 _20481_ (.A(net3667),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _20482_ (.A0(net3519),
    .A1(net1341),
    .S(_03845_),
    .X(_03865_));
 sky130_fd_sc_hd__and2_1 _20483_ (.A(_03858_),
    .B(net3520),
    .X(_03866_));
 sky130_fd_sc_hd__clkbuf_1 _20484_ (.A(net3521),
    .X(_01212_));
 sky130_fd_sc_hd__clkbuf_4 _20485_ (.A(net3250),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _20486_ (.A0(net3775),
    .A1(net1475),
    .S(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__and2_1 _20487_ (.A(_03858_),
    .B(net3776),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_1 _20488_ (.A(net3777),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _20489_ (.A0(net3139),
    .A1(net3530),
    .S(_03867_),
    .X(_03870_));
 sky130_fd_sc_hd__and2_1 _20490_ (.A(_03858_),
    .B(net3531),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _20491_ (.A(net3532),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _20492_ (.A0(net3337),
    .A1(net1491),
    .S(_03867_),
    .X(_03872_));
 sky130_fd_sc_hd__and2_1 _20493_ (.A(_03858_),
    .B(net3338),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _20494_ (.A(net3339),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _20495_ (.A0(net3305),
    .A1(net1318),
    .S(_03867_),
    .X(_03874_));
 sky130_fd_sc_hd__and2_1 _20496_ (.A(_03858_),
    .B(net3306),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_1 _20497_ (.A(net3307),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _20498_ (.A0(net3301),
    .A1(net1284),
    .S(_03867_),
    .X(_03876_));
 sky130_fd_sc_hd__and2_1 _20499_ (.A(_03858_),
    .B(net3302),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_1 _20500_ (.A(net3303),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _20501_ (.A0(net3440),
    .A1(net1228),
    .S(_03867_),
    .X(_03878_));
 sky130_fd_sc_hd__and2_1 _20502_ (.A(_03858_),
    .B(net3441),
    .X(_03879_));
 sky130_fd_sc_hd__clkbuf_1 _20503_ (.A(net3442),
    .X(_01218_));
 sky130_fd_sc_hd__buf_2 _20504_ (.A(_08274_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_1 _20505_ (.A0(net3365),
    .A1(net1290),
    .S(_03867_),
    .X(_03881_));
 sky130_fd_sc_hd__and2_1 _20506_ (.A(_03880_),
    .B(net3366),
    .X(_03882_));
 sky130_fd_sc_hd__clkbuf_1 _20507_ (.A(net3367),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _20508_ (.A0(net3573),
    .A1(net1270),
    .S(_03867_),
    .X(_03883_));
 sky130_fd_sc_hd__and2_1 _20509_ (.A(_03880_),
    .B(net3574),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_1 _20510_ (.A(net3575),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _20511_ (.A0(net3713),
    .A1(net1375),
    .S(_03867_),
    .X(_03885_));
 sky130_fd_sc_hd__and2_1 _20512_ (.A(_03880_),
    .B(net3714),
    .X(_03886_));
 sky130_fd_sc_hd__clkbuf_1 _20513_ (.A(net3715),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _20514_ (.A0(net3611),
    .A1(net1324),
    .S(_03867_),
    .X(_03887_));
 sky130_fd_sc_hd__and2_1 _20515_ (.A(_03880_),
    .B(net3612),
    .X(_03888_));
 sky130_fd_sc_hd__clkbuf_1 _20516_ (.A(net3613),
    .X(_01222_));
 sky130_fd_sc_hd__clkbuf_4 _20517_ (.A(net3249),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _20518_ (.A0(net2990),
    .A1(net3275),
    .S(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__and2_1 _20519_ (.A(_03880_),
    .B(net3276),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_1 _20520_ (.A(net3277),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _20521_ (.A0(net3580),
    .A1(net1493),
    .S(_03889_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _20522_ (.A(_03880_),
    .B(net3581),
    .X(_03893_));
 sky130_fd_sc_hd__clkbuf_1 _20523_ (.A(net3582),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _20524_ (.A0(net2956),
    .A1(net3342),
    .S(_03889_),
    .X(_03894_));
 sky130_fd_sc_hd__and2_1 _20525_ (.A(_03880_),
    .B(net3343),
    .X(_03895_));
 sky130_fd_sc_hd__clkbuf_1 _20526_ (.A(net3344),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _20527_ (.A0(net2914),
    .A1(net3435),
    .S(_03889_),
    .X(_03896_));
 sky130_fd_sc_hd__and2_1 _20528_ (.A(_03880_),
    .B(net3436),
    .X(_03897_));
 sky130_fd_sc_hd__clkbuf_1 _20529_ (.A(net3437),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _20530_ (.A0(net1018),
    .A1(net3800),
    .S(_03889_),
    .X(_03898_));
 sky130_fd_sc_hd__and2_1 _20531_ (.A(_03880_),
    .B(net3801),
    .X(_03899_));
 sky130_fd_sc_hd__clkbuf_1 _20532_ (.A(net3802),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _20533_ (.A0(net3360),
    .A1(net1337),
    .S(_03889_),
    .X(_03900_));
 sky130_fd_sc_hd__and2_1 _20534_ (.A(_03880_),
    .B(net3361),
    .X(_03901_));
 sky130_fd_sc_hd__clkbuf_1 _20535_ (.A(net3362),
    .X(_01228_));
 sky130_fd_sc_hd__clkbuf_2 _20536_ (.A(_08274_),
    .X(_03902_));
 sky130_fd_sc_hd__mux2_1 _20537_ (.A0(net3286),
    .A1(net1400),
    .S(_03889_),
    .X(_03903_));
 sky130_fd_sc_hd__and2_1 _20538_ (.A(_03902_),
    .B(net3287),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_1 _20539_ (.A(net3288),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _20540_ (.A0(net668),
    .A1(net3598),
    .S(_03889_),
    .X(_03905_));
 sky130_fd_sc_hd__and2_1 _20541_ (.A(_03902_),
    .B(net3599),
    .X(_03906_));
 sky130_fd_sc_hd__clkbuf_1 _20542_ (.A(net3600),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _20543_ (.A0(net747),
    .A1(net3646),
    .S(_03889_),
    .X(_03907_));
 sky130_fd_sc_hd__and2_1 _20544_ (.A(_03902_),
    .B(net3647),
    .X(_03908_));
 sky130_fd_sc_hd__clkbuf_1 _20545_ (.A(net3648),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _20546_ (.A0(net3081),
    .A1(net3568),
    .S(_03889_),
    .X(_03909_));
 sky130_fd_sc_hd__and2_1 _20547_ (.A(_03902_),
    .B(net3569),
    .X(_03910_));
 sky130_fd_sc_hd__clkbuf_1 _20548_ (.A(net3570),
    .X(_01232_));
 sky130_fd_sc_hd__clkbuf_4 _20549_ (.A(net3249),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_1 _20550_ (.A0(net3483),
    .A1(net1265),
    .S(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__and2_1 _20551_ (.A(_03902_),
    .B(net3484),
    .X(_03913_));
 sky130_fd_sc_hd__clkbuf_1 _20552_ (.A(net3485),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _20553_ (.A0(net733),
    .A1(net3488),
    .S(_03911_),
    .X(_03914_));
 sky130_fd_sc_hd__and2_1 _20554_ (.A(_03902_),
    .B(net3489),
    .X(_03915_));
 sky130_fd_sc_hd__clkbuf_1 _20555_ (.A(net3490),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _20556_ (.A0(net1156),
    .A1(net3476),
    .S(_03911_),
    .X(_03916_));
 sky130_fd_sc_hd__and2_1 _20557_ (.A(_03902_),
    .B(net3477),
    .X(_03917_));
 sky130_fd_sc_hd__clkbuf_1 _20558_ (.A(net3478),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _20559_ (.A0(net3258),
    .A1(net1282),
    .S(_03911_),
    .X(_03918_));
 sky130_fd_sc_hd__and2_1 _20560_ (.A(_03902_),
    .B(net3259),
    .X(_03919_));
 sky130_fd_sc_hd__clkbuf_1 _20561_ (.A(net3260),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _20562_ (.A0(net3030),
    .A1(net3705),
    .S(_03911_),
    .X(_03920_));
 sky130_fd_sc_hd__and2_1 _20563_ (.A(_03902_),
    .B(net3706),
    .X(_03921_));
 sky130_fd_sc_hd__clkbuf_1 _20564_ (.A(net3707),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _20565_ (.A0(net3732),
    .A1(net1209),
    .S(_03911_),
    .X(_03922_));
 sky130_fd_sc_hd__and2_1 _20566_ (.A(_03902_),
    .B(net3733),
    .X(_03923_));
 sky130_fd_sc_hd__clkbuf_1 _20567_ (.A(net3734),
    .X(_01238_));
 sky130_fd_sc_hd__clkbuf_2 _20568_ (.A(_08274_),
    .X(_03924_));
 sky130_fd_sc_hd__mux2_1 _20569_ (.A0(net2944),
    .A1(net3812),
    .S(_03911_),
    .X(_03925_));
 sky130_fd_sc_hd__and2_1 _20570_ (.A(_03924_),
    .B(net3813),
    .X(_03926_));
 sky130_fd_sc_hd__clkbuf_1 _20571_ (.A(net3814),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _20572_ (.A0(net2927),
    .A1(net3752),
    .S(_03911_),
    .X(_03927_));
 sky130_fd_sc_hd__and2_1 _20573_ (.A(_03924_),
    .B(net3753),
    .X(_03928_));
 sky130_fd_sc_hd__clkbuf_1 _20574_ (.A(net3754),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _20575_ (.A0(net2999),
    .A1(net3670),
    .S(_03911_),
    .X(_03929_));
 sky130_fd_sc_hd__and2_1 _20576_ (.A(_03924_),
    .B(net3671),
    .X(_03930_));
 sky130_fd_sc_hd__clkbuf_1 _20577_ (.A(net3672),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _20578_ (.A0(net1013),
    .A1(net3679),
    .S(_03911_),
    .X(_03931_));
 sky130_fd_sc_hd__and2_1 _20579_ (.A(_03924_),
    .B(net3680),
    .X(_03932_));
 sky130_fd_sc_hd__clkbuf_1 _20580_ (.A(net3681),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _20581_ (.A0(net744),
    .A1(net3514),
    .S(net3250),
    .X(_03933_));
 sky130_fd_sc_hd__and2_1 _20582_ (.A(_03924_),
    .B(net3515),
    .X(_03934_));
 sky130_fd_sc_hd__clkbuf_1 _20583_ (.A(net3516),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _20584_ (.A0(net2812),
    .A1(net3496),
    .S(net3250),
    .X(_03935_));
 sky130_fd_sc_hd__and2_1 _20585_ (.A(_03924_),
    .B(net3497),
    .X(_03936_));
 sky130_fd_sc_hd__clkbuf_1 _20586_ (.A(net3498),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _20587_ (.A0(net675),
    .A1(net3383),
    .S(net3250),
    .X(_03937_));
 sky130_fd_sc_hd__and2_1 _20588_ (.A(_03924_),
    .B(net3384),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_1 _20589_ (.A(net3385),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _20590_ (.A0(net3524),
    .A1(net1302),
    .S(net3250),
    .X(_03939_));
 sky130_fd_sc_hd__and2_1 _20591_ (.A(_03924_),
    .B(net3525),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_1 _20592_ (.A(net3526),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _20593_ (.A0(net3310),
    .A1(net1508),
    .S(net3250),
    .X(_03941_));
 sky130_fd_sc_hd__and2_1 _20594_ (.A(_03924_),
    .B(net3311),
    .X(_03942_));
 sky130_fd_sc_hd__clkbuf_1 _20595_ (.A(net3312),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _20596_ (.A0(net3156),
    .A1(net1187),
    .S(net3250),
    .X(_03943_));
 sky130_fd_sc_hd__and2_1 _20597_ (.A(_03924_),
    .B(net3251),
    .X(_03944_));
 sky130_fd_sc_hd__clkbuf_1 _20598_ (.A(net3252),
    .X(_01248_));
 sky130_fd_sc_hd__nor3b_1 _20599_ (.A(net2938),
    .B(_03782_),
    .C_N(net3562),
    .Y(_01249_));
 sky130_fd_sc_hd__and2_1 _20600_ (.A(net56),
    .B(_03026_),
    .X(_03945_));
 sky130_fd_sc_hd__clkbuf_1 _20601_ (.A(_03945_),
    .X(_01250_));
 sky130_fd_sc_hd__and2_1 _20602_ (.A(net6365),
    .B(_03026_),
    .X(_03946_));
 sky130_fd_sc_hd__clkbuf_1 _20603_ (.A(net1108),
    .X(_01251_));
 sky130_fd_sc_hd__or3b_1 _20604_ (.A(_04881_),
    .B(_05816_),
    .C_N(_03033_),
    .X(_03947_));
 sky130_fd_sc_hd__nor2_1 _20605_ (.A(net4014),
    .B(net3965),
    .Y(_03948_));
 sky130_fd_sc_hd__and4bb_1 _20606_ (.A_N(_03947_),
    .B_N(net4021),
    .C(_05825_),
    .D(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__or4b_1 _20607_ (.A(net4014),
    .B(_05825_),
    .C(net3965),
    .D_N(net4021),
    .X(_03950_));
 sky130_fd_sc_hd__o221a_1 _20608_ (.A1(net4103),
    .A2(net6266),
    .B1(net4015),
    .B2(_03947_),
    .C1(_08276_),
    .X(_01252_));
 sky130_fd_sc_hd__or4b_1 _20609_ (.A(_04162_),
    .B(_04601_),
    .C(net2987),
    .D_N(_09924_),
    .X(_03951_));
 sky130_fd_sc_hd__nor2_1 _20610_ (.A(_04777_),
    .B(net2987),
    .Y(_03952_));
 sky130_fd_sc_hd__a41o_1 _20611_ (.A1(_04760_),
    .A2(_04166_),
    .A3(_04852_),
    .A4(_03952_),
    .B1(net4962),
    .X(_03953_));
 sky130_fd_sc_hd__o211a_1 _20612_ (.A1(_04777_),
    .A2(net2988),
    .B1(_03953_),
    .C1(_08276_),
    .X(_01253_));
 sky130_fd_sc_hd__or3b_1 _20613_ (.A(net3930),
    .B(_05196_),
    .C_N(net3937),
    .X(_03954_));
 sky130_fd_sc_hd__or4_1 _20614_ (.A(net4002),
    .B(_04802_),
    .C(net4015),
    .D(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__inv_2 _20615_ (.A(net4016),
    .Y(_03956_));
 sky130_fd_sc_hd__nor2_1 _20616_ (.A(_09929_),
    .B(net4017),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2_1 _20617_ (.A(net3965),
    .B(net3979),
    .Y(_03958_));
 sky130_fd_sc_hd__o211a_1 _20618_ (.A1(net3965),
    .A2(net4018),
    .B1(net3966),
    .C1(_08276_),
    .X(_01254_));
 sky130_fd_sc_hd__inv_2 _20619_ (.A(_05825_),
    .Y(_03959_));
 sky130_fd_sc_hd__a31o_1 _20620_ (.A1(_05825_),
    .A2(net3965),
    .A3(net3979),
    .B1(_04597_),
    .X(_03960_));
 sky130_fd_sc_hd__a21oi_1 _20621_ (.A1(_03959_),
    .A2(net3966),
    .B1(_03960_),
    .Y(_01255_));
 sky130_fd_sc_hd__inv_2 _20622_ (.A(net3898),
    .Y(_03961_));
 sky130_fd_sc_hd__a22o_1 _20623_ (.A1(net4021),
    .A2(_09929_),
    .B1(_03961_),
    .B2(net4018),
    .X(_03962_));
 sky130_fd_sc_hd__a21o_1 _20624_ (.A1(_05825_),
    .A2(net3965),
    .B1(net4021),
    .X(_03963_));
 sky130_fd_sc_hd__and3_1 _20625_ (.A(_02992_),
    .B(_03962_),
    .C(net4022),
    .X(_03964_));
 sky130_fd_sc_hd__clkbuf_1 _20626_ (.A(net4023),
    .X(_01256_));
 sky130_fd_sc_hd__a22o_1 _20627_ (.A1(_05299_),
    .A2(_09929_),
    .B1(_03031_),
    .B2(_03957_),
    .X(_03965_));
 sky130_fd_sc_hd__o211a_1 _20628_ (.A1(_05299_),
    .A2(net3898),
    .B1(_03965_),
    .C1(_08276_),
    .X(_01257_));
 sky130_fd_sc_hd__a21oi_1 _20629_ (.A1(_05816_),
    .A2(_03032_),
    .B1(_03083_),
    .Y(_03966_));
 sky130_fd_sc_hd__o21a_1 _20630_ (.A1(_05816_),
    .A2(_03032_),
    .B1(_03966_),
    .X(_01258_));
 sky130_fd_sc_hd__and3_1 _20631_ (.A(net4060),
    .B(_05816_),
    .C(_03032_),
    .X(_03967_));
 sky130_fd_sc_hd__a21o_1 _20632_ (.A1(_05816_),
    .A2(_03032_),
    .B1(net4060),
    .X(_03968_));
 sky130_fd_sc_hd__and3b_1 _20633_ (.A_N(net4061),
    .B(_08275_),
    .C(net4100),
    .X(_03969_));
 sky130_fd_sc_hd__clkbuf_1 _20634_ (.A(net4101),
    .X(_01259_));
 sky130_fd_sc_hd__and2_1 _20635_ (.A(_04802_),
    .B(net4061),
    .X(_03970_));
 sky130_fd_sc_hd__nor2_1 _20636_ (.A(_03083_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__o21a_1 _20637_ (.A1(_04802_),
    .A2(net4061),
    .B1(_03971_),
    .X(_01260_));
 sky130_fd_sc_hd__and3_1 _20638_ (.A(net4002),
    .B(_04802_),
    .C(net4061),
    .X(_03972_));
 sky130_fd_sc_hd__nor2_1 _20639_ (.A(_03083_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__o21a_1 _20640_ (.A1(net4002),
    .A2(_03970_),
    .B1(_03973_),
    .X(_01261_));
 sky130_fd_sc_hd__and2_1 _20641_ (.A(net3930),
    .B(_03972_),
    .X(_03974_));
 sky130_fd_sc_hd__nor2_1 _20642_ (.A(_03083_),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__o21a_1 _20643_ (.A1(net3930),
    .A2(_03972_),
    .B1(_03975_),
    .X(_01262_));
 sky130_fd_sc_hd__a221o_1 _20644_ (.A1(net3979),
    .A2(net4017),
    .B1(_03974_),
    .B2(net3937),
    .C1(_04597_),
    .X(_03976_));
 sky130_fd_sc_hd__o21ba_1 _20645_ (.A1(net3937),
    .A2(_03974_),
    .B1_N(_03976_),
    .X(_01263_));
 sky130_fd_sc_hd__and2_2 _20646_ (.A(net46),
    .B(_03026_),
    .X(_03977_));
 sky130_fd_sc_hd__clkbuf_1 _20647_ (.A(_03977_),
    .X(_01264_));
 sky130_fd_sc_hd__and2_1 _20648_ (.A(net6363),
    .B(_03026_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _20649_ (.A(net1173),
    .X(_01265_));
 sky130_fd_sc_hd__and2_1 _20650_ (.A(net6557),
    .B(_03026_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_1 _20651_ (.A(net1578),
    .X(_01266_));
 sky130_fd_sc_hd__inv_2 _20652__91 (.A(clknet_1_1__leaf__03781_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _20653__92 (.A(clknet_1_1__leaf__03781_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _20654__93 (.A(clknet_1_1__leaf__03781_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _20655__94 (.A(clknet_1_1__leaf__03781_),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _20656__95 (.A(clknet_1_1__leaf__03781_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _20657__96 (.A(clknet_1_1__leaf__03781_),
    .Y(net235));
 sky130_fd_sc_hd__buf_1 _20658_ (.A(clknet_1_1__leaf__03780_),
    .X(_03980_));
 sky130_fd_sc_hd__inv_2 _20659__97 (.A(clknet_1_0__leaf__03980_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20660__98 (.A(clknet_1_0__leaf__03980_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20661__99 (.A(clknet_1_0__leaf__03980_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _20662__100 (.A(clknet_1_0__leaf__03980_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20663__101 (.A(clknet_1_1__leaf__03980_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _20664__102 (.A(clknet_1_1__leaf__03980_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _20665__103 (.A(clknet_1_1__leaf__03980_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20666__104 (.A(clknet_1_1__leaf__03980_),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _20667__105 (.A(clknet_1_1__leaf__03980_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _20668__106 (.A(clknet_1_1__leaf__03980_),
    .Y(net245));
 sky130_fd_sc_hd__buf_1 _20669_ (.A(clknet_1_1__leaf__03780_),
    .X(_03981_));
 sky130_fd_sc_hd__inv_2 _20670__107 (.A(clknet_1_1__leaf__03981_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20671__108 (.A(clknet_1_1__leaf__03981_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20672__109 (.A(clknet_1_1__leaf__03981_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _20673__110 (.A(clknet_1_1__leaf__03981_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20674__111 (.A(clknet_1_1__leaf__03981_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _20675__112 (.A(clknet_1_1__leaf__03981_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _20676__113 (.A(clknet_1_0__leaf__03981_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20677__114 (.A(clknet_1_0__leaf__03981_),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _20678__115 (.A(clknet_1_0__leaf__03981_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _20679__116 (.A(clknet_1_0__leaf__03981_),
    .Y(net255));
 sky130_fd_sc_hd__buf_1 _20680_ (.A(clknet_1_1__leaf__03780_),
    .X(_03982_));
 sky130_fd_sc_hd__inv_2 _20681__117 (.A(clknet_1_0__leaf__03982_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20682__118 (.A(clknet_1_0__leaf__03982_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20683__119 (.A(clknet_1_0__leaf__03982_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _20684__120 (.A(clknet_1_0__leaf__03982_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20685__121 (.A(clknet_1_0__leaf__03982_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _20686__122 (.A(clknet_1_0__leaf__03982_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _20687__123 (.A(clknet_1_1__leaf__03982_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20688__124 (.A(clknet_1_1__leaf__03982_),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _20689__125 (.A(clknet_1_1__leaf__03982_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _20690__126 (.A(clknet_1_1__leaf__03982_),
    .Y(net265));
 sky130_fd_sc_hd__buf_1 _20691_ (.A(clknet_1_1__leaf__03780_),
    .X(_03983_));
 sky130_fd_sc_hd__inv_2 _20692__127 (.A(clknet_1_0__leaf__03983_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20693__128 (.A(clknet_1_0__leaf__03983_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20694__129 (.A(clknet_1_0__leaf__03983_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _20695__130 (.A(clknet_1_1__leaf__03983_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20696__131 (.A(clknet_1_1__leaf__03983_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _20697__132 (.A(clknet_1_1__leaf__03983_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _20698__133 (.A(clknet_1_1__leaf__03983_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20699__134 (.A(clknet_1_1__leaf__03983_),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _20700__135 (.A(clknet_1_1__leaf__03983_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _20701__136 (.A(clknet_1_0__leaf__03983_),
    .Y(net275));
 sky130_fd_sc_hd__buf_1 _20702_ (.A(clknet_1_1__leaf__03780_),
    .X(_03984_));
 sky130_fd_sc_hd__inv_2 _20703__137 (.A(clknet_1_1__leaf__03984_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20704__138 (.A(clknet_1_1__leaf__03984_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20705__139 (.A(clknet_1_1__leaf__03984_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _20706__140 (.A(clknet_1_0__leaf__03984_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20707__141 (.A(clknet_1_0__leaf__03984_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _20708__142 (.A(clknet_1_0__leaf__03984_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _20709__143 (.A(clknet_1_0__leaf__03984_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20710__144 (.A(clknet_1_0__leaf__03984_),
    .Y(net283));
 sky130_fd_sc_hd__inv_2 _20711__145 (.A(clknet_1_0__leaf__03984_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _20712__146 (.A(clknet_1_1__leaf__03984_),
    .Y(net285));
 sky130_fd_sc_hd__buf_1 _20713_ (.A(clknet_1_0__leaf__03780_),
    .X(_03985_));
 sky130_fd_sc_hd__inv_2 _20714__147 (.A(clknet_1_1__leaf__03985_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20715__148 (.A(clknet_1_1__leaf__03985_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20716__149 (.A(clknet_1_1__leaf__03985_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _20717__150 (.A(clknet_1_1__leaf__03985_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20718__151 (.A(clknet_1_1__leaf__03985_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _20719__152 (.A(clknet_1_1__leaf__03985_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _20720__153 (.A(clknet_1_0__leaf__03985_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20721__154 (.A(clknet_1_0__leaf__03985_),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _20722__155 (.A(clknet_1_0__leaf__03985_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _20723__156 (.A(clknet_1_0__leaf__03985_),
    .Y(net295));
 sky130_fd_sc_hd__buf_1 _20724_ (.A(clknet_1_0__leaf__03780_),
    .X(_03986_));
 sky130_fd_sc_hd__inv_2 _20725__157 (.A(clknet_1_1__leaf__03986_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20726__158 (.A(clknet_1_1__leaf__03986_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20727__159 (.A(clknet_1_1__leaf__03986_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _20728__160 (.A(clknet_1_1__leaf__03986_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20729__161 (.A(clknet_1_1__leaf__03986_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _20730__162 (.A(clknet_1_0__leaf__03986_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _20731__163 (.A(clknet_1_0__leaf__03986_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20732__164 (.A(clknet_1_0__leaf__03986_),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _20733__165 (.A(clknet_1_0__leaf__03986_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _20734__166 (.A(clknet_1_0__leaf__03986_),
    .Y(net305));
 sky130_fd_sc_hd__buf_1 _20735_ (.A(clknet_1_0__leaf__03780_),
    .X(_03987_));
 sky130_fd_sc_hd__inv_2 _20736__167 (.A(clknet_1_1__leaf__03987_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20737__168 (.A(clknet_1_1__leaf__03987_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20738__169 (.A(clknet_1_1__leaf__03987_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _20739__170 (.A(clknet_1_1__leaf__03987_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20740__171 (.A(clknet_1_0__leaf__03987_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _20741__172 (.A(clknet_1_0__leaf__03987_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _20742__173 (.A(clknet_1_0__leaf__03987_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20743__174 (.A(clknet_1_0__leaf__03987_),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 _20744__175 (.A(clknet_1_0__leaf__03987_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _20745__176 (.A(clknet_1_0__leaf__03987_),
    .Y(net315));
 sky130_fd_sc_hd__buf_1 _20746_ (.A(clknet_1_0__leaf__03780_),
    .X(_03988_));
 sky130_fd_sc_hd__inv_2 _20747__177 (.A(clknet_1_0__leaf__03988_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20748__178 (.A(clknet_1_0__leaf__03988_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20749__179 (.A(clknet_1_0__leaf__03988_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _20750__180 (.A(clknet_1_0__leaf__03988_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20751__181 (.A(clknet_1_0__leaf__03988_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _20752__182 (.A(clknet_1_0__leaf__03988_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _20753__183 (.A(clknet_1_1__leaf__03988_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20754__184 (.A(clknet_1_1__leaf__03988_),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _20755__185 (.A(clknet_1_1__leaf__03988_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _20756__186 (.A(clknet_1_1__leaf__03988_),
    .Y(net325));
 sky130_fd_sc_hd__buf_1 _20757_ (.A(clknet_1_0__leaf__04800_),
    .X(_03989_));
 sky130_fd_sc_hd__buf_1 _20758_ (.A(clknet_1_0__leaf__03989_),
    .X(_03990_));
 sky130_fd_sc_hd__inv_2 _20759__187 (.A(clknet_1_0__leaf__03990_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20760__188 (.A(clknet_1_0__leaf__03990_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20761__189 (.A(clknet_1_0__leaf__03990_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _20762__190 (.A(clknet_1_0__leaf__03990_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20763__191 (.A(clknet_1_0__leaf__03990_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _20764__192 (.A(clknet_1_1__leaf__03990_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _20765__193 (.A(clknet_1_1__leaf__03990_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20766__194 (.A(clknet_1_1__leaf__03990_),
    .Y(net333));
 sky130_fd_sc_hd__inv_2 _20767__195 (.A(clknet_1_1__leaf__03990_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _20768__196 (.A(clknet_1_1__leaf__03990_),
    .Y(net335));
 sky130_fd_sc_hd__buf_1 _20769_ (.A(clknet_1_0__leaf__03989_),
    .X(_03991_));
 sky130_fd_sc_hd__inv_2 _20770__197 (.A(clknet_1_1__leaf__03991_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20771__198 (.A(clknet_1_1__leaf__03991_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20772__199 (.A(clknet_1_1__leaf__03991_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _20773__200 (.A(clknet_1_1__leaf__03991_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20774__201 (.A(clknet_1_1__leaf__03991_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _20775__202 (.A(clknet_1_0__leaf__03991_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _20776__203 (.A(clknet_1_0__leaf__03991_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20777__204 (.A(clknet_1_0__leaf__03991_),
    .Y(net343));
 sky130_fd_sc_hd__inv_2 _20778__205 (.A(clknet_1_0__leaf__03991_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _20779__206 (.A(clknet_1_0__leaf__03991_),
    .Y(net345));
 sky130_fd_sc_hd__buf_1 _20780_ (.A(clknet_1_0__leaf__03989_),
    .X(_03992_));
 sky130_fd_sc_hd__inv_2 _20781__207 (.A(clknet_1_0__leaf__03992_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20782__208 (.A(clknet_1_0__leaf__03992_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20783__209 (.A(clknet_1_0__leaf__03992_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _20784__210 (.A(clknet_1_0__leaf__03992_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20785__211 (.A(clknet_1_0__leaf__03992_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _20786__212 (.A(clknet_1_1__leaf__03992_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _20787__213 (.A(clknet_1_1__leaf__03992_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20788__214 (.A(clknet_1_1__leaf__03992_),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _20789__215 (.A(clknet_1_1__leaf__03992_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _20790__216 (.A(clknet_1_1__leaf__03992_),
    .Y(net355));
 sky130_fd_sc_hd__buf_1 _20791_ (.A(clknet_1_0__leaf__03989_),
    .X(_03993_));
 sky130_fd_sc_hd__inv_2 _20792__217 (.A(clknet_1_0__leaf__03993_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20793__218 (.A(clknet_1_0__leaf__03993_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20794__219 (.A(clknet_1_1__leaf__03993_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _20795__220 (.A(clknet_1_1__leaf__03993_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20796__221 (.A(clknet_1_1__leaf__03993_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _20797__222 (.A(clknet_1_1__leaf__03993_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _20798__223 (.A(clknet_1_0__leaf__03993_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20799__224 (.A(clknet_1_0__leaf__03993_),
    .Y(net363));
 sky130_fd_sc_hd__inv_2 _20800__225 (.A(clknet_1_0__leaf__03993_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _20801__226 (.A(clknet_1_0__leaf__03993_),
    .Y(net365));
 sky130_fd_sc_hd__buf_1 _20802_ (.A(clknet_1_1__leaf__03989_),
    .X(_03994_));
 sky130_fd_sc_hd__inv_2 _20803__227 (.A(clknet_1_0__leaf__03994_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20804__228 (.A(clknet_1_1__leaf__03994_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20805__229 (.A(clknet_1_1__leaf__03994_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _20806__230 (.A(clknet_1_1__leaf__03994_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20807__231 (.A(clknet_1_0__leaf__03994_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _20808__232 (.A(clknet_1_0__leaf__03994_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _20809__233 (.A(clknet_1_0__leaf__03994_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20810__234 (.A(clknet_1_1__leaf__03994_),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _20811__235 (.A(clknet_1_1__leaf__03994_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _20812__236 (.A(clknet_1_1__leaf__03994_),
    .Y(net375));
 sky130_fd_sc_hd__buf_1 _20813_ (.A(clknet_1_1__leaf__03989_),
    .X(_03995_));
 sky130_fd_sc_hd__inv_2 _20814__237 (.A(clknet_1_1__leaf__03995_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20815__238 (.A(clknet_1_1__leaf__03995_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20816__239 (.A(clknet_1_1__leaf__03995_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _20817__240 (.A(clknet_1_1__leaf__03995_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20818__241 (.A(clknet_1_1__leaf__03995_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _20819__242 (.A(clknet_1_1__leaf__03995_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _20820__243 (.A(clknet_1_0__leaf__03995_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20821__244 (.A(clknet_1_0__leaf__03995_),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _20822__245 (.A(clknet_1_0__leaf__03995_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _20823__246 (.A(clknet_1_0__leaf__03995_),
    .Y(net385));
 sky130_fd_sc_hd__buf_1 _20824_ (.A(clknet_1_1__leaf__03989_),
    .X(_03996_));
 sky130_fd_sc_hd__inv_2 _20825__247 (.A(clknet_1_1__leaf__03996_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20826__248 (.A(clknet_1_1__leaf__03996_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20827__249 (.A(clknet_1_0__leaf__03996_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _20828__250 (.A(clknet_1_0__leaf__03996_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20829__251 (.A(clknet_1_0__leaf__03996_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _20830__252 (.A(clknet_1_0__leaf__03996_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _20831__253 (.A(clknet_1_0__leaf__03996_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20832__254 (.A(clknet_1_1__leaf__03996_),
    .Y(net393));
 sky130_fd_sc_hd__inv_2 _20833__255 (.A(clknet_1_1__leaf__03996_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _20834__256 (.A(clknet_1_1__leaf__03996_),
    .Y(net395));
 sky130_fd_sc_hd__buf_1 _20835_ (.A(clknet_1_1__leaf__03989_),
    .X(_03997_));
 sky130_fd_sc_hd__inv_2 _20836__257 (.A(clknet_1_1__leaf__03997_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20837__258 (.A(clknet_1_1__leaf__03997_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20838__259 (.A(clknet_1_1__leaf__03997_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _20839__260 (.A(clknet_1_1__leaf__03997_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20840__261 (.A(clknet_1_0__leaf__03997_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _20841__262 (.A(clknet_1_0__leaf__03997_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _20842__263 (.A(clknet_1_0__leaf__03997_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20843__264 (.A(clknet_1_0__leaf__03997_),
    .Y(net403));
 sky130_fd_sc_hd__inv_2 _20844__265 (.A(clknet_1_0__leaf__03997_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _20845__266 (.A(clknet_1_0__leaf__03997_),
    .Y(net405));
 sky130_fd_sc_hd__buf_1 _20846_ (.A(clknet_1_1__leaf__03989_),
    .X(_03998_));
 sky130_fd_sc_hd__inv_2 _20847__267 (.A(clknet_1_1__leaf__03998_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20848__268 (.A(clknet_1_1__leaf__03998_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20849__269 (.A(clknet_1_1__leaf__03998_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _20850__270 (.A(clknet_1_1__leaf__03998_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20851__271 (.A(clknet_1_1__leaf__03998_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _20852__272 (.A(clknet_1_0__leaf__03998_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _20853__273 (.A(clknet_1_0__leaf__03998_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20854__274 (.A(clknet_1_0__leaf__03998_),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _20855__275 (.A(clknet_1_0__leaf__03998_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _20856__276 (.A(clknet_1_0__leaf__03998_),
    .Y(net415));
 sky130_fd_sc_hd__buf_1 _20857_ (.A(clknet_1_0__leaf__03989_),
    .X(_03999_));
 sky130_fd_sc_hd__inv_2 _20858__277 (.A(clknet_1_0__leaf__03999_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20859__278 (.A(clknet_1_0__leaf__03999_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20860__279 (.A(clknet_1_0__leaf__03999_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _20861__280 (.A(clknet_1_0__leaf__03999_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20862__281 (.A(clknet_1_0__leaf__03999_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _20863__282 (.A(clknet_1_0__leaf__03999_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _20864__283 (.A(clknet_1_1__leaf__03999_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20865__284 (.A(clknet_1_1__leaf__03999_),
    .Y(net423));
 sky130_fd_sc_hd__inv_2 _20866__285 (.A(clknet_1_1__leaf__03999_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _20867__286 (.A(clknet_1_1__leaf__03999_),
    .Y(net425));
 sky130_fd_sc_hd__buf_1 _20868_ (.A(clknet_1_0__leaf__04800_),
    .X(_04000_));
 sky130_fd_sc_hd__buf_1 _20869_ (.A(clknet_1_1__leaf__04000_),
    .X(_04001_));
 sky130_fd_sc_hd__inv_2 _20870__287 (.A(clknet_1_1__leaf__04001_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20871__288 (.A(clknet_1_1__leaf__04001_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20872__289 (.A(clknet_1_1__leaf__04001_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _20873__290 (.A(clknet_1_1__leaf__04001_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20874__291 (.A(clknet_1_1__leaf__04001_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _20875__292 (.A(clknet_1_1__leaf__04001_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _20876__293 (.A(clknet_1_0__leaf__04001_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20877__294 (.A(clknet_1_0__leaf__04001_),
    .Y(net433));
 sky130_fd_sc_hd__inv_2 _20878__295 (.A(clknet_1_0__leaf__04001_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _20879__296 (.A(clknet_1_0__leaf__04001_),
    .Y(net435));
 sky130_fd_sc_hd__buf_1 _20880_ (.A(clknet_1_1__leaf__04000_),
    .X(_04002_));
 sky130_fd_sc_hd__inv_2 _20881__297 (.A(clknet_1_1__leaf__04002_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20882__298 (.A(clknet_1_1__leaf__04002_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20883__299 (.A(clknet_1_1__leaf__04002_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _20884__300 (.A(clknet_1_1__leaf__04002_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20885__301 (.A(clknet_1_1__leaf__04002_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _20886__302 (.A(clknet_1_0__leaf__04002_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _20887__303 (.A(clknet_1_0__leaf__04002_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20888__304 (.A(clknet_1_0__leaf__04002_),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 _20889__305 (.A(clknet_1_0__leaf__04002_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _20890__306 (.A(clknet_1_0__leaf__04002_),
    .Y(net445));
 sky130_fd_sc_hd__buf_1 _20891_ (.A(clknet_1_1__leaf__04000_),
    .X(_04003_));
 sky130_fd_sc_hd__inv_2 _20892__307 (.A(clknet_1_0__leaf__04003_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20893__308 (.A(clknet_1_0__leaf__04003_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20894__309 (.A(clknet_1_0__leaf__04003_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _20895__310 (.A(clknet_1_0__leaf__04003_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20896__311 (.A(clknet_1_1__leaf__04003_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _20897__312 (.A(clknet_1_1__leaf__04003_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _20898__313 (.A(clknet_1_1__leaf__04003_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20899__314 (.A(clknet_1_1__leaf__04003_),
    .Y(net453));
 sky130_fd_sc_hd__inv_2 _20900__315 (.A(clknet_1_1__leaf__04003_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _20901__316 (.A(clknet_1_1__leaf__04003_),
    .Y(net455));
 sky130_fd_sc_hd__buf_1 _20902_ (.A(clknet_1_1__leaf__04000_),
    .X(_04004_));
 sky130_fd_sc_hd__inv_2 _20903__317 (.A(clknet_1_0__leaf__04004_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20904__318 (.A(clknet_1_0__leaf__04004_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20905__319 (.A(clknet_1_0__leaf__04004_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _20906__320 (.A(clknet_1_0__leaf__04004_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20907__321 (.A(clknet_1_0__leaf__04004_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _20908__322 (.A(clknet_1_1__leaf__04004_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _20909__323 (.A(clknet_1_1__leaf__04004_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20910__324 (.A(clknet_1_1__leaf__04004_),
    .Y(net463));
 sky130_fd_sc_hd__inv_2 _20911__325 (.A(clknet_1_1__leaf__04004_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _20912__326 (.A(clknet_1_1__leaf__04004_),
    .Y(net465));
 sky130_fd_sc_hd__buf_1 _20913_ (.A(clknet_1_1__leaf__04000_),
    .X(_04005_));
 sky130_fd_sc_hd__inv_2 _20914__327 (.A(clknet_1_1__leaf__04005_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20915__328 (.A(clknet_1_1__leaf__04005_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20916__329 (.A(clknet_1_1__leaf__04005_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _20917__330 (.A(clknet_1_1__leaf__04005_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20918__331 (.A(clknet_1_1__leaf__04005_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _20919__332 (.A(clknet_1_0__leaf__04005_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _20920__333 (.A(clknet_1_0__leaf__04005_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20921__334 (.A(clknet_1_0__leaf__04005_),
    .Y(net473));
 sky130_fd_sc_hd__inv_2 _20922__335 (.A(clknet_1_0__leaf__04005_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _20923__336 (.A(clknet_1_0__leaf__04005_),
    .Y(net475));
 sky130_fd_sc_hd__buf_1 _20924_ (.A(clknet_1_1__leaf__04000_),
    .X(_04006_));
 sky130_fd_sc_hd__inv_2 _20925__337 (.A(clknet_1_0__leaf__04006_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20926__338 (.A(clknet_1_0__leaf__04006_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20927__339 (.A(clknet_1_0__leaf__04006_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _20928__340 (.A(clknet_1_0__leaf__04006_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20929__341 (.A(clknet_1_0__leaf__04006_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _20930__342 (.A(clknet_1_1__leaf__04006_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _20931__343 (.A(clknet_1_1__leaf__04006_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20932__344 (.A(clknet_1_1__leaf__04006_),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _20933__345 (.A(clknet_1_1__leaf__04006_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _20934__346 (.A(clknet_1_1__leaf__04006_),
    .Y(net485));
 sky130_fd_sc_hd__buf_1 _20935_ (.A(clknet_1_0__leaf__04000_),
    .X(_04007_));
 sky130_fd_sc_hd__inv_2 _20936__347 (.A(clknet_1_1__leaf__04007_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20937__348 (.A(clknet_1_1__leaf__04007_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20938__349 (.A(clknet_1_1__leaf__04007_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _20939__350 (.A(clknet_1_1__leaf__04007_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20940__351 (.A(clknet_1_1__leaf__04007_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _20941__352 (.A(clknet_1_0__leaf__04007_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _20942__353 (.A(clknet_1_0__leaf__04007_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20943__354 (.A(clknet_1_0__leaf__04007_),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _20944__355 (.A(clknet_1_0__leaf__04007_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _20945__356 (.A(clknet_1_0__leaf__04007_),
    .Y(net495));
 sky130_fd_sc_hd__buf_1 _20946_ (.A(clknet_1_0__leaf__04000_),
    .X(_04008_));
 sky130_fd_sc_hd__inv_2 _20947__357 (.A(clknet_1_1__leaf__04008_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20948__358 (.A(clknet_1_1__leaf__04008_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20949__359 (.A(clknet_1_1__leaf__04008_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _20950__360 (.A(clknet_1_1__leaf__04008_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20951__361 (.A(clknet_1_1__leaf__04008_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _20952__362 (.A(clknet_1_1__leaf__04008_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _20953__363 (.A(clknet_1_0__leaf__04008_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20954__364 (.A(clknet_1_0__leaf__04008_),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _20955__365 (.A(clknet_1_0__leaf__04008_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _20956__366 (.A(clknet_1_0__leaf__04008_),
    .Y(net505));
 sky130_fd_sc_hd__buf_1 _20957_ (.A(clknet_1_0__leaf__04000_),
    .X(_04009_));
 sky130_fd_sc_hd__inv_2 _20958__367 (.A(clknet_1_1__leaf__04009_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20959__368 (.A(clknet_1_1__leaf__04009_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20960__369 (.A(clknet_1_1__leaf__04009_),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _20961__370 (.A(clknet_1_1__leaf__04009_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _20962__371 (.A(clknet_1_0__leaf__04009_),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _20963__372 (.A(clknet_1_0__leaf__04009_),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _20964__373 (.A(clknet_1_0__leaf__04009_),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _20965__374 (.A(clknet_1_0__leaf__04009_),
    .Y(net513));
 sky130_fd_sc_hd__inv_2 _20966__375 (.A(clknet_1_0__leaf__04009_),
    .Y(net514));
 sky130_fd_sc_hd__inv_2 _20967__376 (.A(clknet_1_0__leaf__04009_),
    .Y(net515));
 sky130_fd_sc_hd__buf_1 _20968_ (.A(clknet_1_0__leaf__04000_),
    .X(_04010_));
 sky130_fd_sc_hd__inv_2 _20969__377 (.A(clknet_1_1__leaf__04010_),
    .Y(net516));
 sky130_fd_sc_hd__inv_2 _20970__378 (.A(clknet_1_1__leaf__04010_),
    .Y(net517));
 sky130_fd_sc_hd__inv_2 _20971__379 (.A(clknet_1_1__leaf__04010_),
    .Y(net518));
 sky130_fd_sc_hd__inv_2 _20972__380 (.A(clknet_1_1__leaf__04010_),
    .Y(net519));
 sky130_fd_sc_hd__inv_2 _20973__381 (.A(clknet_1_1__leaf__04010_),
    .Y(net520));
 sky130_fd_sc_hd__inv_2 _20974__382 (.A(clknet_1_0__leaf__04010_),
    .Y(net521));
 sky130_fd_sc_hd__inv_2 _20975__383 (.A(clknet_1_0__leaf__04010_),
    .Y(net522));
 sky130_fd_sc_hd__inv_2 _20976__384 (.A(clknet_1_0__leaf__04010_),
    .Y(net523));
 sky130_fd_sc_hd__inv_2 _20977__385 (.A(clknet_1_0__leaf__04010_),
    .Y(net524));
 sky130_fd_sc_hd__inv_2 _20978__386 (.A(clknet_1_0__leaf__04010_),
    .Y(net525));
 sky130_fd_sc_hd__buf_1 _20979_ (.A(clknet_1_0__leaf__04800_),
    .X(_04011_));
 sky130_fd_sc_hd__inv_2 _20980__7 (.A(clknet_1_0__leaf__04011_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20981__8 (.A(clknet_1_0__leaf__04011_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20982__9 (.A(clknet_1_0__leaf__04011_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _20983__10 (.A(clknet_1_0__leaf__04011_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _20984__11 (.A(clknet_1_0__leaf__04011_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _20985__12 (.A(clknet_1_1__leaf__04011_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _20986__13 (.A(clknet_1_1__leaf__04011_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _20987__14 (.A(clknet_1_1__leaf__04011_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _20988__15 (.A(clknet_1_1__leaf__04011_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _20989__16 (.A(clknet_1_1__leaf__04011_),
    .Y(net155));
 sky130_fd_sc_hd__buf_1 _20990_ (.A(clknet_1_0__leaf__04800_),
    .X(_04012_));
 sky130_fd_sc_hd__inv_2 _20991__17 (.A(clknet_1_0__leaf__04012_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _20992__18 (.A(clknet_1_0__leaf__04012_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _20993__19 (.A(clknet_1_0__leaf__04012_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _20994__20 (.A(clknet_1_0__leaf__04012_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _20995__21 (.A(clknet_1_1__leaf__04012_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _20996__22 (.A(clknet_1_1__leaf__04012_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _20997__23 (.A(clknet_1_1__leaf__04012_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _20998__24 (.A(clknet_1_1__leaf__04012_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _20999__25 (.A(clknet_1_1__leaf__04012_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _21000__26 (.A(clknet_1_1__leaf__04012_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _21001__3 (.A(clknet_1_0__leaf__03773_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _21002__4 (.A(clknet_1_0__leaf__03773_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _21003__5 (.A(clknet_1_0__leaf__03773_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _21004__6 (.A(clknet_1_0__leaf__03773_),
    .Y(net145));
 sky130_fd_sc_hd__nor2_1 _21005_ (.A(net4945),
    .B(net65),
    .Y(_01587_));
 sky130_fd_sc_hd__xnor2_1 _21006_ (.A(net6347),
    .B(net4945),
    .Y(_04013_));
 sky130_fd_sc_hd__nor2_1 _21007_ (.A(_03502_),
    .B(net1081),
    .Y(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _21008_ (.A(_09920_),
    .X(_04014_));
 sky130_fd_sc_hd__or2_1 _21009_ (.A(net773),
    .B(net4987),
    .X(_04015_));
 sky130_fd_sc_hd__nand2_1 _21010_ (.A(net773),
    .B(net4987),
    .Y(_04016_));
 sky130_fd_sc_hd__clkbuf_4 _21011_ (.A(_04597_),
    .X(_04017_));
 sky130_fd_sc_hd__a32o_1 _21012_ (.A1(_04014_),
    .A2(_04015_),
    .A3(_04016_),
    .B1(_04017_),
    .B2(net4987),
    .X(_01589_));
 sky130_fd_sc_hd__clkbuf_4 _21013_ (.A(_09920_),
    .X(_04018_));
 sky130_fd_sc_hd__or2_1 _21014_ (.A(net839),
    .B(net4975),
    .X(_04019_));
 sky130_fd_sc_hd__nand2_1 _21015_ (.A(net839),
    .B(net4975),
    .Y(_04020_));
 sky130_fd_sc_hd__nand3b_1 _21016_ (.A_N(_04016_),
    .B(_04019_),
    .C(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21bo_1 _21017_ (.A1(_04019_),
    .A2(_04020_),
    .B1_N(_04016_),
    .X(_04022_));
 sky130_fd_sc_hd__a32o_1 _21018_ (.A1(_04018_),
    .A2(_04021_),
    .A3(_04022_),
    .B1(_04017_),
    .B2(net4975),
    .X(_01590_));
 sky130_fd_sc_hd__and2_1 _21019_ (.A(_04020_),
    .B(_04021_),
    .X(_04023_));
 sky130_fd_sc_hd__nor2_1 _21020_ (.A(net1011),
    .B(net5271),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _21021_ (.A(net1011),
    .B(net5271),
    .Y(_04025_));
 sky130_fd_sc_hd__or2b_1 _21022_ (.A(_04024_),
    .B_N(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__xor2_1 _21023_ (.A(_04023_),
    .B(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__a22o_1 _21024_ (.A1(net5271),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04027_),
    .X(_01591_));
 sky130_fd_sc_hd__o21a_1 _21025_ (.A1(_04023_),
    .A2(_04024_),
    .B1(_04025_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_1 _21026_ (.A(net890),
    .B(net5334),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _21027_ (.A(net890),
    .B(net5334),
    .Y(_04030_));
 sky130_fd_sc_hd__and2b_1 _21028_ (.A_N(_04029_),
    .B(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__xnor2_1 _21029_ (.A(_04028_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__a22o_1 _21030_ (.A1(net5334),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04032_),
    .X(_01592_));
 sky130_fd_sc_hd__o21a_1 _21031_ (.A1(_04028_),
    .A2(_04029_),
    .B1(_04030_),
    .X(_04033_));
 sky130_fd_sc_hd__nor2_1 _21032_ (.A(net5379),
    .B(net5168),
    .Y(_04034_));
 sky130_fd_sc_hd__nand2_1 _21033_ (.A(net5379),
    .B(net5168),
    .Y(_04035_));
 sky130_fd_sc_hd__and2b_1 _21034_ (.A_N(_04034_),
    .B(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__xnor2_1 _21035_ (.A(_04033_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__a22o_1 _21036_ (.A1(net5168),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04037_),
    .X(_01593_));
 sky130_fd_sc_hd__o21a_1 _21037_ (.A1(_04033_),
    .A2(_04034_),
    .B1(_04035_),
    .X(_04038_));
 sky130_fd_sc_hd__nor2_1 _21038_ (.A(net985),
    .B(net5424),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _21039_ (.A(net985),
    .B(net5424),
    .Y(_04040_));
 sky130_fd_sc_hd__and2b_1 _21040_ (.A_N(_04039_),
    .B(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__xnor2_1 _21041_ (.A(_04038_),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__a22o_1 _21042_ (.A1(net5424),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04042_),
    .X(_01594_));
 sky130_fd_sc_hd__o21a_1 _21043_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_04040_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_1 _21044_ (.A(net5310),
    .B(net5455),
    .Y(_04044_));
 sky130_fd_sc_hd__nand2_1 _21045_ (.A(net5310),
    .B(net5455),
    .Y(_04045_));
 sky130_fd_sc_hd__and2b_1 _21046_ (.A_N(_04044_),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__xnor2_1 _21047_ (.A(_04043_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__a22o_1 _21048_ (.A1(net5455),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04047_),
    .X(_01595_));
 sky130_fd_sc_hd__o21a_1 _21049_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_04045_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_1 _21050_ (.A(net4152),
    .B(net4763),
    .Y(_04049_));
 sky130_fd_sc_hd__nand2_1 _21051_ (.A(net4152),
    .B(net4763),
    .Y(_04050_));
 sky130_fd_sc_hd__and2b_1 _21052_ (.A_N(_04049_),
    .B(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__xnor2_1 _21053_ (.A(_04048_),
    .B(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__a22o_1 _21054_ (.A1(net4763),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04052_),
    .X(_01596_));
 sky130_fd_sc_hd__o21a_1 _21055_ (.A1(_04048_),
    .A2(_04049_),
    .B1(_04050_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_1 _21056_ (.A(net4146),
    .B(net4736),
    .Y(_04054_));
 sky130_fd_sc_hd__nand2_1 _21057_ (.A(net4146),
    .B(net4736),
    .Y(_04055_));
 sky130_fd_sc_hd__and2b_1 _21058_ (.A_N(_04054_),
    .B(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__xnor2_1 _21059_ (.A(_04053_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__a22o_1 _21060_ (.A1(net4736),
    .A2(_03519_),
    .B1(_04014_),
    .B2(_04057_),
    .X(_01597_));
 sky130_fd_sc_hd__o21ai_2 _21061_ (.A1(_04053_),
    .A2(_04054_),
    .B1(_04055_),
    .Y(_04058_));
 sky130_fd_sc_hd__or2_1 _21062_ (.A(net4130),
    .B(net4395),
    .X(_04059_));
 sky130_fd_sc_hd__nand2_1 _21063_ (.A(net4130),
    .B(net4395),
    .Y(_04060_));
 sky130_fd_sc_hd__nand3_1 _21064_ (.A(_04058_),
    .B(_04059_),
    .C(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__a21o_1 _21065_ (.A1(_04059_),
    .A2(_04060_),
    .B1(_04058_),
    .X(_04062_));
 sky130_fd_sc_hd__a32o_1 _21066_ (.A1(_04018_),
    .A2(_04061_),
    .A3(_04062_),
    .B1(_04017_),
    .B2(net4395),
    .X(_01598_));
 sky130_fd_sc_hd__or2_1 _21067_ (.A(net4173),
    .B(net4546),
    .X(_04063_));
 sky130_fd_sc_hd__nand2_1 _21068_ (.A(net4173),
    .B(net4546),
    .Y(_04064_));
 sky130_fd_sc_hd__a21bo_1 _21069_ (.A1(_04058_),
    .A2(_04059_),
    .B1_N(_04060_),
    .X(_04065_));
 sky130_fd_sc_hd__and3_1 _21070_ (.A(_04063_),
    .B(_04064_),
    .C(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__inv_2 _21071_ (.A(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a21o_1 _21072_ (.A1(_04063_),
    .A2(_04064_),
    .B1(_04065_),
    .X(_04068_));
 sky130_fd_sc_hd__a32o_1 _21073_ (.A1(_04018_),
    .A2(_04067_),
    .A3(_04068_),
    .B1(_04017_),
    .B2(net4546),
    .X(_01599_));
 sky130_fd_sc_hd__or2_1 _21074_ (.A(net4167),
    .B(net4503),
    .X(_04069_));
 sky130_fd_sc_hd__nand2_1 _21075_ (.A(net4167),
    .B(net4503),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_1 _21076_ (.A(_04064_),
    .B(_04067_),
    .Y(_04071_));
 sky130_fd_sc_hd__a21o_1 _21077_ (.A1(_04069_),
    .A2(_04070_),
    .B1(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__and3_1 _21078_ (.A(_04069_),
    .B(_04070_),
    .C(_04071_),
    .X(_04073_));
 sky130_fd_sc_hd__inv_2 _21079_ (.A(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__a32o_1 _21080_ (.A1(_04018_),
    .A2(_04072_),
    .A3(_04074_),
    .B1(_04017_),
    .B2(net4503),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _21081_ (.A(net4179),
    .B(net4542),
    .X(_04075_));
 sky130_fd_sc_hd__nand2_1 _21082_ (.A(net4179),
    .B(net4542),
    .Y(_04076_));
 sky130_fd_sc_hd__nand2_1 _21083_ (.A(_04070_),
    .B(_04074_),
    .Y(_04077_));
 sky130_fd_sc_hd__and3_1 _21084_ (.A(_04075_),
    .B(_04076_),
    .C(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__inv_2 _21085_ (.A(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__a21o_1 _21086_ (.A1(_04075_),
    .A2(_04076_),
    .B1(_04077_),
    .X(_04080_));
 sky130_fd_sc_hd__a32o_1 _21087_ (.A1(_04018_),
    .A2(_04079_),
    .A3(_04080_),
    .B1(_04017_),
    .B2(net4542),
    .X(_01601_));
 sky130_fd_sc_hd__or2_1 _21088_ (.A(net1100),
    .B(net4701),
    .X(_04081_));
 sky130_fd_sc_hd__nand2_1 _21089_ (.A(net1100),
    .B(net4701),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _21090_ (.A(_04076_),
    .B(_04079_),
    .Y(_04083_));
 sky130_fd_sc_hd__a21o_1 _21091_ (.A1(_04081_),
    .A2(_04082_),
    .B1(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__and3_1 _21092_ (.A(_04081_),
    .B(_04082_),
    .C(_04083_),
    .X(_04085_));
 sky130_fd_sc_hd__inv_2 _21093_ (.A(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__a32o_1 _21094_ (.A1(_04018_),
    .A2(_04084_),
    .A3(_04086_),
    .B1(_04017_),
    .B2(net4701),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _21095_ (.A(net4936),
    .B(net1886),
    .X(_04087_));
 sky130_fd_sc_hd__nand2_1 _21096_ (.A(net4936),
    .B(net1886),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _21097_ (.A(_04082_),
    .B(_04086_),
    .Y(_04089_));
 sky130_fd_sc_hd__and3_1 _21098_ (.A(_04087_),
    .B(net4937),
    .C(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__inv_2 _21099_ (.A(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21o_1 _21100_ (.A1(_04087_),
    .A2(net4937),
    .B1(_04089_),
    .X(_04092_));
 sky130_fd_sc_hd__a32o_1 _21101_ (.A1(_04018_),
    .A2(_04091_),
    .A3(net4938),
    .B1(_04017_),
    .B2(net1886),
    .X(_01603_));
 sky130_fd_sc_hd__or2_1 _21102_ (.A(net4186),
    .B(net4469),
    .X(_04093_));
 sky130_fd_sc_hd__nand2_1 _21103_ (.A(net4186),
    .B(net4469),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_1 _21104_ (.A(_04088_),
    .B(_04091_),
    .Y(_04095_));
 sky130_fd_sc_hd__a21o_1 _21105_ (.A1(_04093_),
    .A2(_04094_),
    .B1(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__nand3_1 _21106_ (.A(_04093_),
    .B(_04094_),
    .C(_04095_),
    .Y(_04097_));
 sky130_fd_sc_hd__a32o_1 _21107_ (.A1(_04018_),
    .A2(_04096_),
    .A3(_04097_),
    .B1(_03083_),
    .B2(net4469),
    .X(_01604_));
 sky130_fd_sc_hd__a21boi_1 _21108_ (.A1(_04093_),
    .A2(_04095_),
    .B1_N(_04094_),
    .Y(_04098_));
 sky130_fd_sc_hd__nor2_1 _21109_ (.A(net4143),
    .B(net4649),
    .Y(_04099_));
 sky130_fd_sc_hd__and2_1 _21110_ (.A(net4143),
    .B(net4649),
    .X(_04100_));
 sky130_fd_sc_hd__or3_1 _21111_ (.A(_04098_),
    .B(_04099_),
    .C(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__o21ai_1 _21112_ (.A1(_04099_),
    .A2(_04100_),
    .B1(_04098_),
    .Y(_04102_));
 sky130_fd_sc_hd__a32o_1 _21113_ (.A1(_04018_),
    .A2(_04101_),
    .A3(_04102_),
    .B1(_03083_),
    .B2(net4649),
    .X(_01605_));
 sky130_fd_sc_hd__o21ba_1 _21114_ (.A1(_04098_),
    .A2(_04099_),
    .B1_N(_04100_),
    .X(_04103_));
 sky130_fd_sc_hd__nor2_1 _21115_ (.A(net4160),
    .B(net4653),
    .Y(_04104_));
 sky130_fd_sc_hd__and2_1 _21116_ (.A(net4160),
    .B(net4653),
    .X(_04105_));
 sky130_fd_sc_hd__or3_1 _21117_ (.A(_04103_),
    .B(_04104_),
    .C(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__o21ai_1 _21118_ (.A1(_04104_),
    .A2(_04105_),
    .B1(_04103_),
    .Y(_04107_));
 sky130_fd_sc_hd__a32o_1 _21119_ (.A1(_04018_),
    .A2(_04106_),
    .A3(_04107_),
    .B1(_03083_),
    .B2(net4653),
    .X(_01606_));
 sky130_fd_sc_hd__o21ba_1 _21120_ (.A1(_04103_),
    .A2(_04104_),
    .B1_N(_04105_),
    .X(_04108_));
 sky130_fd_sc_hd__nor2_1 _21121_ (.A(net4176),
    .B(net4744),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_1 _21122_ (.A(net4176),
    .B(net4744),
    .Y(_04110_));
 sky130_fd_sc_hd__and2b_1 _21123_ (.A_N(_04109_),
    .B(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__xnor2_1 _21124_ (.A(_04108_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__a22o_1 _21125_ (.A1(net4744),
    .A2(_04017_),
    .B1(_04014_),
    .B2(_04112_),
    .X(_01607_));
 sky130_fd_sc_hd__o21a_1 _21126_ (.A1(_04108_),
    .A2(_04109_),
    .B1(_04110_),
    .X(_04113_));
 sky130_fd_sc_hd__nor2_1 _21127_ (.A(net4133),
    .B(net4740),
    .Y(_04114_));
 sky130_fd_sc_hd__and2_1 _21128_ (.A(net4133),
    .B(net4740),
    .X(_04115_));
 sky130_fd_sc_hd__nor2_1 _21129_ (.A(_04114_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__xnor2_1 _21130_ (.A(_04113_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__a22o_1 _21131_ (.A1(net4740),
    .A2(_04017_),
    .B1(_04014_),
    .B2(_04117_),
    .X(_01608_));
 sky130_fd_sc_hd__nor2_1 _21132_ (.A(_04113_),
    .B(_04114_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand2_2 _21133_ (.A(net4136),
    .B(net4679),
    .Y(_04119_));
 sky130_fd_sc_hd__or2_1 _21134_ (.A(net4136),
    .B(net4679),
    .X(_04120_));
 sky130_fd_sc_hd__o211ai_2 _21135_ (.A1(_04115_),
    .A2(_04118_),
    .B1(_04119_),
    .C1(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a211o_1 _21136_ (.A1(_04120_),
    .A2(_04119_),
    .B1(_04118_),
    .C1(_04115_),
    .X(_04122_));
 sky130_fd_sc_hd__a32o_1 _21137_ (.A1(_09920_),
    .A2(_04121_),
    .A3(_04122_),
    .B1(_03083_),
    .B2(net4679),
    .X(_01609_));
 sky130_fd_sc_hd__xnor2_1 _21138_ (.A(net4155),
    .B(net4705),
    .Y(_04123_));
 sky130_fd_sc_hd__a21oi_1 _21139_ (.A1(_04119_),
    .A2(_04121_),
    .B1(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__a31o_1 _21140_ (.A1(_04119_),
    .A2(_04121_),
    .A3(_04123_),
    .B1(_09919_),
    .X(_04125_));
 sky130_fd_sc_hd__a2bb2o_1 _21141_ (.A1_N(_04124_),
    .A2_N(_04125_),
    .B1(net4705),
    .B2(net65),
    .X(_01610_));
 sky130_fd_sc_hd__o21ai_1 _21142_ (.A1(_04626_),
    .A2(_04818_),
    .B1(net4027),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _21143_ (.A(_04627_),
    .B(net3979),
    .Y(_04127_));
 sky130_fd_sc_hd__a41o_1 _21144_ (.A1(net3402),
    .A2(net2982),
    .A3(_04626_),
    .A4(net3980),
    .B1(_08200_),
    .X(_04128_));
 sky130_fd_sc_hd__mux2_1 _21145_ (.A0(net4028),
    .A1(net4027),
    .S(net3981),
    .X(_04129_));
 sky130_fd_sc_hd__and2_1 _21146_ (.A(_08195_),
    .B(net4029),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _21147_ (.A(net4030),
    .X(_01611_));
 sky130_fd_sc_hd__o211a_1 _21148_ (.A1(net3535),
    .A2(net3981),
    .B1(_08195_),
    .C1(net3507),
    .X(_01612_));
 sky130_fd_sc_hd__o21ai_1 _21149_ (.A1(net3535),
    .A2(net3981),
    .B1(net2982),
    .Y(_04131_));
 sky130_fd_sc_hd__or3_1 _21150_ (.A(net6168),
    .B(net3535),
    .C(_08200_),
    .X(_04132_));
 sky130_fd_sc_hd__a21oi_1 _21151_ (.A1(net2983),
    .A2(_04132_),
    .B1(_04633_),
    .Y(_01613_));
 sky130_fd_sc_hd__o21ai_1 _21152_ (.A1(_04626_),
    .A2(_04818_),
    .B1(net4910),
    .Y(_04133_));
 sky130_fd_sc_hd__o31a_1 _21153_ (.A1(_09486_),
    .A2(net3981),
    .A3(_04133_),
    .B1(_01622_),
    .X(_01614_));
 sky130_fd_sc_hd__and2_2 _21154_ (.A(_02488_),
    .B(clknet_1_1__leaf__05840_),
    .X(_04134_));
 sky130_fd_sc_hd__buf_1 _21155_ (.A(_04134_),
    .X(_01615_));
 sky130_fd_sc_hd__and2_2 _21156_ (.A(_02488_),
    .B(clknet_1_0__leaf__05891_),
    .X(_04135_));
 sky130_fd_sc_hd__buf_1 _21157_ (.A(_04135_),
    .X(_01616_));
 sky130_fd_sc_hd__and2_2 _21158_ (.A(_02488_),
    .B(clknet_1_0__leaf__05942_),
    .X(_04136_));
 sky130_fd_sc_hd__buf_1 _21159_ (.A(_04136_),
    .X(_01617_));
 sky130_fd_sc_hd__and2_2 _21160_ (.A(_02488_),
    .B(clknet_1_0__leaf__05994_),
    .X(_04137_));
 sky130_fd_sc_hd__buf_1 _21161_ (.A(_04137_),
    .X(_01618_));
 sky130_fd_sc_hd__and2_2 _21162_ (.A(_02488_),
    .B(clknet_1_0__leaf__06044_),
    .X(_04138_));
 sky130_fd_sc_hd__buf_1 _21163_ (.A(_04138_),
    .X(_01619_));
 sky130_fd_sc_hd__and2_2 _21164_ (.A(_02488_),
    .B(clknet_1_0__leaf__06092_),
    .X(_04139_));
 sky130_fd_sc_hd__buf_1 _21165_ (.A(_04139_),
    .X(_01620_));
 sky130_fd_sc_hd__nor2_1 _21166_ (.A(net4962),
    .B(net65),
    .Y(_01621_));
 sky130_fd_sc_hd__a22o_1 _21167_ (.A1(net4111),
    .A2(_09941_),
    .B1(_09942_),
    .B2(_09284_),
    .X(_01623_));
 sky130_fd_sc_hd__clkbuf_4 _21168_ (.A(_09933_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_4 _21169_ (.A(_09935_),
    .X(_04141_));
 sky130_fd_sc_hd__a22o_1 _21170_ (.A1(net4190),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09281_),
    .X(_01624_));
 sky130_fd_sc_hd__a22o_1 _21171_ (.A1(net4159),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09276_),
    .X(_01625_));
 sky130_fd_sc_hd__a22o_1 _21172_ (.A1(net4183),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09403_),
    .X(_01626_));
 sky130_fd_sc_hd__a22o_1 _21173_ (.A1(net4164),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09521_),
    .X(_01627_));
 sky130_fd_sc_hd__a22o_1 _21174_ (.A1(net4166),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09642_),
    .X(_01628_));
 sky130_fd_sc_hd__a22o_1 _21175_ (.A1(net4140),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09769_),
    .X(_01629_));
 sky130_fd_sc_hd__a22o_1 _21176_ (.A1(net4142),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_09908_),
    .X(_01630_));
 sky130_fd_sc_hd__a22o_1 _21177_ (.A1(net4185),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_10205_),
    .X(_01631_));
 sky130_fd_sc_hd__a22o_1 _21178_ (.A1(net4201),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_10329_),
    .X(_01632_));
 sky130_fd_sc_hd__a22o_1 _21179_ (.A1(net4231),
    .A2(_04140_),
    .B1(_04141_),
    .B2(_10454_),
    .X(_01633_));
 sky130_fd_sc_hd__nor2_1 _21180_ (.A(net4951),
    .B(net65),
    .Y(_01634_));
 sky130_fd_sc_hd__xnor2_1 _21181_ (.A(net6349),
    .B(net4951),
    .Y(_04142_));
 sky130_fd_sc_hd__nor2_1 _21182_ (.A(_03502_),
    .B(net1128),
    .Y(_01635_));
 sky130_fd_sc_hd__or2_1 _21183_ (.A(net4424),
    .B(net701),
    .X(_04143_));
 sky130_fd_sc_hd__a32o_1 _21184_ (.A1(_02529_),
    .A2(net4425),
    .A3(_04143_),
    .B1(_02528_),
    .B2(net701),
    .X(_01636_));
 sky130_fd_sc_hd__a21bo_1 _21185_ (.A1(_02532_),
    .A2(net4657),
    .B1_N(net4425),
    .X(_04144_));
 sky130_fd_sc_hd__a32o_1 _21186_ (.A1(_02529_),
    .A2(_02535_),
    .A3(net4658),
    .B1(_02528_),
    .B2(net715),
    .X(_01637_));
 sky130_fd_sc_hd__or2b_1 _21187_ (.A(_02531_),
    .B_N(_02537_),
    .X(_04145_));
 sky130_fd_sc_hd__xor2_1 _21188_ (.A(_02536_),
    .B(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__a22o_1 _21189_ (.A1(net4806),
    .A2(_02528_),
    .B1(_02579_),
    .B2(_04146_),
    .X(_01638_));
 sky130_fd_sc_hd__and2b_1 _21190_ (.A_N(_02530_),
    .B(net4477),
    .X(_04147_));
 sky130_fd_sc_hd__xnor2_1 _21191_ (.A(_02538_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__a22o_1 _21192_ (.A1(net4791),
    .A2(_02528_),
    .B1(_02579_),
    .B2(_04148_),
    .X(_01639_));
 sky130_fd_sc_hd__or2_1 _21193_ (.A(net4438),
    .B(net723),
    .X(_04149_));
 sky130_fd_sc_hd__a32o_1 _21194_ (.A1(_02529_),
    .A2(net4439),
    .A3(_04149_),
    .B1(_02528_),
    .B2(net723),
    .X(_01640_));
 sky130_fd_sc_hd__a21bo_1 _21195_ (.A1(_02752_),
    .A2(net4621),
    .B1_N(net4439),
    .X(_04150_));
 sky130_fd_sc_hd__a32o_1 _21196_ (.A1(_02529_),
    .A2(_02755_),
    .A3(net4622),
    .B1(_02528_),
    .B2(net738),
    .X(_01641_));
 sky130_fd_sc_hd__or2b_1 _21197_ (.A(_02751_),
    .B_N(_02757_),
    .X(_04151_));
 sky130_fd_sc_hd__xor2_1 _21198_ (.A(_02756_),
    .B(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__a22o_1 _21199_ (.A1(net4905),
    .A2(_02528_),
    .B1(_02579_),
    .B2(_04152_),
    .X(_01642_));
 sky130_fd_sc_hd__and2b_1 _21200_ (.A_N(_02750_),
    .B(net4800),
    .X(_04153_));
 sky130_fd_sc_hd__xnor2_1 _21201_ (.A(_02758_),
    .B(net4801),
    .Y(_04154_));
 sky130_fd_sc_hd__a22o_1 _21202_ (.A1(net941),
    .A2(_02528_),
    .B1(_02579_),
    .B2(net4802),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_1 _21203_ (.A(net4956),
    .B(net65),
    .Y(_01644_));
 sky130_fd_sc_hd__xnor2_1 _21204_ (.A(net660),
    .B(net6555),
    .Y(_04155_));
 sky130_fd_sc_hd__nor2_1 _21205_ (.A(_03502_),
    .B(net1921),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _21206_ (.A(net4942),
    .B(net65),
    .Y(_01646_));
 sky130_fd_sc_hd__xnor2_1 _21207_ (.A(net4942),
    .B(net6355),
    .Y(_04156_));
 sky130_fd_sc_hd__nor2_1 _21208_ (.A(_03502_),
    .B(net1183),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(net4965),
    .B(net65),
    .Y(_01648_));
 sky130_fd_sc_hd__xnor2_1 _21210_ (.A(net4965),
    .B(net6357),
    .Y(_04157_));
 sky130_fd_sc_hd__nor2_1 _21211_ (.A(_03502_),
    .B(net1136),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _21212_ (.A(net4959),
    .B(net65),
    .Y(_01650_));
 sky130_fd_sc_hd__xnor2_1 _21213_ (.A(net6341),
    .B(net4959),
    .Y(_04158_));
 sky130_fd_sc_hd__nor2_1 _21214_ (.A(_03502_),
    .B(net1048),
    .Y(_01651_));
 sky130_fd_sc_hd__dfxtp_2 _21215_ (.CLK(clknet_leaf_74_i_clk),
    .D(net4949),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21216_ (.CLK(clknet_leaf_75_i_clk),
    .D(net4734),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_43_i_clk),
    .D(net4826),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_43_i_clk),
    .D(net5708),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_43_i_clk),
    .D(net4889),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21220_ (.CLK(clknet_leaf_43_i_clk),
    .D(net5493),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_43_i_clk),
    .D(net1065),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00391_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00392_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00393_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00394_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00395_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00396_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00397_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00398_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00399_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00400_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21244_ (.CLK(clknet_leaf_53_i_clk),
    .D(net3724),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _21245_ (.CLK(clknet_leaf_53_i_clk),
    .D(net3541),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _21246_ (.CLK(clknet_leaf_55_i_clk),
    .D(net3792),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21247_ (.CLK(clknet_leaf_53_i_clk),
    .D(net3335),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21248_ (.CLK(clknet_leaf_54_i_clk),
    .D(net3208),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_50_i_clk),
    .D(net3358),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_50_i_clk),
    .D(net3264),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_51_i_clk),
    .D(net3464),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_52_i_clk),
    .D(net3202),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_52_i_clk),
    .D(net3068),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_52_i_clk),
    .D(net3049),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_52_i_clk),
    .D(net3188),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_52_i_clk),
    .D(net4786),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_71_i_clk),
    .D(net4584),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(clknet_leaf_71_i_clk),
    .D(net3632),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(clknet_leaf_52_i_clk),
    .D(net3224),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(clknet_leaf_71_i_clk),
    .D(net3629),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21261_ (.CLK(clknet_leaf_71_i_clk),
    .D(net3720),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(clknet_leaf_71_i_clk),
    .D(net3774),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_71_i_clk),
    .D(net3635),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(clknet_leaf_71_i_clk),
    .D(net4782),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_71_i_clk),
    .D(net4831),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21276_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_88_i_clk),
    .D(net4097),
    .Q(\reg_rgb[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_75_i_clk),
    .D(net4008),
    .Q(\reg_rgb[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_89_i_clk),
    .D(net4047),
    .Q(\reg_rgb[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_75_i_clk),
    .D(net4068),
    .Q(\reg_rgb[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_75_i_clk),
    .D(net4085),
    .Q(\reg_rgb[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(clknet_leaf_75_i_clk),
    .D(net4080),
    .Q(\reg_rgb[23] ));
 sky130_fd_sc_hd__dfxtp_2 _21294_ (.CLK(clknet_leaf_27_i_clk),
    .D(net3626),
    .Q(\rbzero.wall_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21295_ (.CLK(clknet_leaf_27_i_clk),
    .D(net3512),
    .Q(\rbzero.wall_hot[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_74_i_clk),
    .D(net4089),
    .Q(\rbzero.side_hot ));
 sky130_fd_sc_hd__dfxtp_2 _21297_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00466_),
    .Q(\rbzero.texu_hot[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00467_),
    .Q(\rbzero.texu_hot[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00468_),
    .Q(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00469_),
    .Q(\rbzero.texu_hot[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21301_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00470_),
    .Q(\rbzero.texu_hot[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21302_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00471_),
    .Q(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00472_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_12_i_clk),
    .D(net3871),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_74_i_clk),
    .D(net3990),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_74_i_clk),
    .D(net3911),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_74_i_clk),
    .D(net3763),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_48_i_clk),
    .D(net4012),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(clknet_leaf_74_i_clk),
    .D(net4040),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00479_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_49_i_clk),
    .D(net4057),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(clknet_leaf_49_i_clk),
    .D(net3994),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_72_i_clk),
    .D(net4534),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_73_i_clk),
    .D(net4276),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00484_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_73_i_clk),
    .D(net4279),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(clknet_leaf_73_i_clk),
    .D(net4266),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(clknet_leaf_72_i_clk),
    .D(net2994),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00488_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00489_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00490_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4241),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4273),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4305),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4282),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4256),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_57_i_clk),
    .D(net4253),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_57_i_clk),
    .D(net4234),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_55_i_clk),
    .D(net4299),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_54_i_clk),
    .D(net4204),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_54_i_clk),
    .D(net5381),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(clknet_leaf_50_i_clk),
    .D(net5473),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_50_i_clk),
    .D(net5312),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_46_i_clk),
    .D(net4154),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_46_i_clk),
    .D(net4148),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4132),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4175),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4169),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4181),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(clknet_leaf_56_i_clk),
    .D(net4287),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(clknet_leaf_56_i_clk),
    .D(net4526),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_40_i_clk),
    .D(net4188),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4145),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4162),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4178),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4135),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4138),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4157),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(clknet_leaf_35_i_clk),
    .D(net3380),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(clknet_leaf_35_i_clk),
    .D(net3220),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4879),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_42_i_clk),
    .D(net5971),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(clknet_leaf_42_i_clk),
    .D(net4924),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(clknet_leaf_41_i_clk),
    .D(net5748),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(clknet_leaf_42_i_clk),
    .D(net5422),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00528_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00529_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00530_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00531_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00532_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00572_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1213),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_29_i_clk),
    .D(net3215),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00575_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(clknet_leaf_24_i_clk),
    .D(net629),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_79_i_clk),
    .D(net4481),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(clknet_leaf_79_i_clk),
    .D(net2921),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21410_ (.CLK(clknet_leaf_79_i_clk),
    .D(net3205),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21411_ (.CLK(clknet_leaf_79_i_clk),
    .D(net3239),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21412_ (.CLK(clknet_leaf_84_i_clk),
    .D(net4694),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21413_ (.CLK(clknet_leaf_84_i_clk),
    .D(net3596),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_84_i_clk),
    .D(net4670),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_78_i_clk),
    .D(net3798),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21416_ (.CLK(clknet_leaf_78_i_clk),
    .D(net4756),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_78_i_clk),
    .D(net3372),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_85_i_clk),
    .D(net4770),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21419_ (.CLK(clknet_leaf_85_i_clk),
    .D(net4699),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_85_i_clk),
    .D(net4814),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_85_i_clk),
    .D(net3196),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_85_i_clk),
    .D(net4789),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_85_i_clk),
    .D(net3199),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(clknet_leaf_45_i_clk),
    .D(net3920),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(clknet_leaf_43_i_clk),
    .D(net3884),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_44_i_clk),
    .D(net3806),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_44_i_clk),
    .D(net3896),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_44_i_clk),
    .D(net3282),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_43_i_clk),
    .D(net3036),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_81_i_clk),
    .D(net4554),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(clknet_leaf_82_i_clk),
    .D(net2886),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21432_ (.CLK(clknet_leaf_80_i_clk),
    .D(net3248),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21433_ (.CLK(clknet_leaf_82_i_clk),
    .D(net3459),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21434_ (.CLK(clknet_leaf_82_i_clk),
    .D(net4629),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(clknet_leaf_82_i_clk),
    .D(net3727),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21436_ (.CLK(clknet_leaf_83_i_clk),
    .D(net4712),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21437_ (.CLK(clknet_leaf_83_i_clk),
    .D(net3165),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21438_ (.CLK(clknet_leaf_83_i_clk),
    .D(net4725),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(clknet_leaf_87_i_clk),
    .D(net3410),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21440_ (.CLK(clknet_leaf_87_i_clk),
    .D(net4761),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21441_ (.CLK(clknet_leaf_88_i_clk),
    .D(net4665),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(clknet_leaf_86_i_clk),
    .D(net4820),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(clknet_leaf_88_i_clk),
    .D(net3137),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(clknet_leaf_86_i_clk),
    .D(net4873),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(clknet_leaf_86_i_clk),
    .D(net3020),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(clknet_leaf_45_i_clk),
    .D(net3824),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(clknet_leaf_47_i_clk),
    .D(net4000),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(clknet_leaf_45_i_clk),
    .D(net3986),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(clknet_leaf_45_i_clk),
    .D(net3924),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(clknet_leaf_46_i_clk),
    .D(net3856),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(clknet_leaf_46_i_clk),
    .D(net3267),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3750),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3892),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3916),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3907),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3888),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3377),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(clknet_leaf_30_i_clk),
    .D(net5621),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(clknet_leaf_25_i_clk),
    .D(net1469),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3951),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3959),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3935),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3947),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3943),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3113),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3051),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3094),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(clknet_leaf_24_i_clk),
    .D(net3053),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3098),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3023),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3039),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3089),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3071),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(clknet_leaf_0_i_clk),
    .D(net3101),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(clknet_leaf_102_i_clk),
    .D(net2844),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(clknet_leaf_102_i_clk),
    .D(net3073),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(clknet_leaf_102_i_clk),
    .D(net3110),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(clknet_leaf_102_i_clk),
    .D(net2972),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4320),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(clknet_leaf_21_i_clk),
    .D(net2963),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(clknet_leaf_21_i_clk),
    .D(net2981),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(clknet_leaf_21_i_clk),
    .D(net2950),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00652_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(clknet_leaf_93_i_clk),
    .D(net623),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(clknet_leaf_93_i_clk),
    .D(net2124),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21486_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2678),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2706),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2918),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2044),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2840),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21491_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2926),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2906),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2865),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2537),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2824),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(clknet_leaf_14_i_clk),
    .D(net4685),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(clknet_leaf_14_i_clk),
    .D(net2775),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(clknet_leaf_13_i_clk),
    .D(net2896),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(clknet_leaf_13_i_clk),
    .D(net2826),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(clknet_leaf_14_i_clk),
    .D(net4347),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(clknet_leaf_14_i_clk),
    .D(net638),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21502_ (.CLK(clknet_leaf_14_i_clk),
    .D(net1186),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(clknet_leaf_14_i_clk),
    .D(net2803),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(clknet_leaf_14_i_clk),
    .D(net2880),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_14_i_clk),
    .D(net2790),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(clknet_leaf_44_i_clk),
    .D(net2792),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_15_i_clk),
    .D(net2727),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1507),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1069),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1009),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(clknet_leaf_44_i_clk),
    .D(net1055),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(clknet_leaf_35_i_clk),
    .D(net1313),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(clknet_leaf_36_i_clk),
    .D(net5515),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(clknet_leaf_36_i_clk),
    .D(net4199),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(clknet_leaf_36_i_clk),
    .D(net5712),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(clknet_leaf_37_i_clk),
    .D(net5658),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(clknet_leaf_37_i_clk),
    .D(net5704),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(clknet_leaf_33_i_clk),
    .D(net1636),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_35_i_clk),
    .D(net3147),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_34_i_clk),
    .D(net5119),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(clknet_leaf_34_i_clk),
    .D(net2967),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(clknet_leaf_28_i_clk),
    .D(net5070),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(clknet_leaf_34_i_clk),
    .D(net2998),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5358),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5332),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_34_i_clk),
    .D(net2976),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_33_i_clk),
    .D(net5328),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(clknet_leaf_28_i_clk),
    .D(net2954),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(clknet_leaf_34_i_clk),
    .D(net5153),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_27_i_clk),
    .D(net3131),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1651),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1530),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1570),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(clknet_leaf_36_i_clk),
    .D(net2195),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(clknet_leaf_36_i_clk),
    .D(net2468),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(clknet_leaf_36_i_clk),
    .D(net1916),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(clknet_leaf_27_i_clk),
    .D(net1828),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(clknet_leaf_28_i_clk),
    .D(net1722),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(clknet_leaf_28_i_clk),
    .D(net1351),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(clknet_leaf_28_i_clk),
    .D(net1594),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(clknet_leaf_28_i_clk),
    .D(net1311),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(clknet_leaf_26_i_clk),
    .D(net1421),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5130),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(clknet_leaf_27_i_clk),
    .D(net877),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(clknet_leaf_27_i_clk),
    .D(net1005),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(clknet_leaf_27_i_clk),
    .D(net1321),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(clknet_leaf_17_i_clk),
    .D(net848),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4123),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4151),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4250),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4129),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1067),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1051),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(clknet_leaf_101_i_clk),
    .D(net918),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(clknet_leaf_101_i_clk),
    .D(net1087),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(clknet_leaf_101_i_clk),
    .D(net1380),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21557_ (.CLK(clknet_leaf_2_i_clk),
    .D(net806),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(clknet_leaf_20_i_clk),
    .D(net820),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21559_ (.CLK(clknet_leaf_19_i_clk),
    .D(net920),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(clknet_leaf_19_i_clk),
    .D(net1053),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(clknet_leaf_19_i_clk),
    .D(net5300),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(clknet_leaf_17_i_clk),
    .D(net5308),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(clknet_leaf_17_i_clk),
    .D(net5269),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5479),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(clknet_leaf_17_i_clk),
    .D(net5344),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(clknet_leaf_17_i_clk),
    .D(net5138),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5028),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5024),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(clknet_leaf_16_i_clk),
    .D(net4997),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(clknet_leaf_17_i_clk),
    .D(net4985),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(clknet_leaf_17_i_clk),
    .D(net4126),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5261),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5184),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5616),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5085),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5055),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(clknet_leaf_4_i_clk),
    .D(net4217),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5316),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5009),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5277),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(clknet_leaf_2_i_clk),
    .D(net893),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21582_ (.CLK(clknet_leaf_21_i_clk),
    .D(net5662),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(clknet_leaf_21_i_clk),
    .D(net5716),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(clknet_leaf_21_i_clk),
    .D(net5726),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(clknet_leaf_21_i_clk),
    .D(net4193),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(clknet_leaf_22_i_clk),
    .D(net5596),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(clknet_leaf_22_i_clk),
    .D(net5644),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(clknet_leaf_23_i_clk),
    .D(net5654),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(clknet_leaf_23_i_clk),
    .D(net5635),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(clknet_leaf_23_i_clk),
    .D(net5676),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(clknet_leaf_23_i_clk),
    .D(net4213),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(clknet_leaf_24_i_clk),
    .D(net5738),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21593_ (.CLK(clknet_leaf_24_i_clk),
    .D(net5760),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(clknet_leaf_23_i_clk),
    .D(net5752),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(clknet_leaf_21_i_clk),
    .D(net4270),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4246),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4229),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4263),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4293),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21600_ (.CLK(clknet_leaf_102_i_clk),
    .D(net4210),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(clknet_leaf_102_i_clk),
    .D(net4207),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(clknet_leaf_102_i_clk),
    .D(net5506),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21603_ (.CLK(clknet_leaf_102_i_clk),
    .D(net5529),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(clknet_leaf_2_i_clk),
    .D(net4172),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21605_ (.CLK(clknet_leaf_1_i_clk),
    .D(net5525),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5489),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5631),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(clknet_leaf_20_i_clk),
    .D(net4196),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5265),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(clknet_leaf_22_i_clk),
    .D(net5149),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(clknet_leaf_22_i_clk),
    .D(net5400),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5437),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_23_i_clk),
    .D(net5340),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21614_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5348),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5538),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5607),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5692),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_17_i_clk),
    .D(net5104),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_18_i_clk),
    .D(net5001),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4120),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4114),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5580),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_5_i_clk),
    .D(net5864),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5145),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5020),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_5_i_clk),
    .D(net5005),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_4_i_clk),
    .D(net5415),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5289),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_2_i_clk),
    .D(net5108),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_19_i_clk),
    .D(net4981),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21631_ (.CLK(clknet_leaf_19_i_clk),
    .D(net5293),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21632_ (.CLK(clknet_leaf_19_i_clk),
    .D(net5093),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_28_i_clk),
    .D(net3257),
    .Q(\rbzero.spi_registers.buf_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_34_i_clk),
    .D(net1597),
    .Q(\rbzero.spi_registers.buf_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21635_ (.CLK(clknet_leaf_32_i_clk),
    .D(net3183),
    .Q(\rbzero.spi_registers.buf_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21636_ (.CLK(clknet_leaf_28_i_clk),
    .D(net1533),
    .Q(\rbzero.spi_registers.buf_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_32_i_clk),
    .D(net3107),
    .Q(\rbzero.spi_registers.buf_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21638_ (.CLK(clknet_leaf_28_i_clk),
    .D(net6227),
    .Q(\rbzero.spi_registers.buf_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_34_i_clk),
    .D(net1536),
    .Q(\rbzero.spi_registers.buf_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_29_i_clk),
    .D(net3080),
    .Q(\rbzero.spi_registers.buf_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21641_ (.CLK(clknet_leaf_34_i_clk),
    .D(net1617),
    .Q(\rbzero.spi_registers.buf_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_29_i_clk),
    .D(net3126),
    .Q(\rbzero.spi_registers.buf_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(clknet_leaf_34_i_clk),
    .D(net1542),
    .Q(\rbzero.spi_registers.buf_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_27_i_clk),
    .D(net3119),
    .Q(\rbzero.spi_registers.buf_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21645_ (.CLK(clknet_leaf_34_i_clk),
    .D(net6273),
    .Q(\rbzero.spi_registers.buf_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21646_ (.CLK(clknet_leaf_33_i_clk),
    .D(net1609),
    .Q(\rbzero.spi_registers.buf_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(clknet_leaf_34_i_clk),
    .D(net2555),
    .Q(\rbzero.spi_registers.buf_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(clknet_leaf_33_i_clk),
    .D(net1737),
    .Q(\rbzero.spi_registers.buf_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21649_ (.CLK(clknet_leaf_33_i_clk),
    .D(net2592),
    .Q(\rbzero.spi_registers.buf_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(clknet_leaf_33_i_clk),
    .D(net5786),
    .Q(\rbzero.spi_registers.buf_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21651_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5257),
    .Q(\rbzero.spi_registers.buf_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5369),
    .Q(\rbzero.spi_registers.buf_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5564),
    .Q(\rbzero.spi_registers.buf_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5112),
    .Q(\rbzero.spi_registers.buf_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(clknet_leaf_15_i_clk),
    .D(net5404),
    .Q(\rbzero.spi_registers.buf_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_15_i_clk),
    .D(net5461),
    .Q(\rbzero.spi_registers.buf_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_15_i_clk),
    .D(net5408),
    .Q(\rbzero.spi_registers.buf_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_15_i_clk),
    .D(net5126),
    .Q(\rbzero.spi_registers.buf_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5047),
    .Q(\rbzero.spi_registers.buf_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_15_i_clk),
    .D(net5377),
    .Q(\rbzero.spi_registers.buf_othery[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5249),
    .Q(\rbzero.spi_registers.buf_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5430),
    .Q(\rbzero.spi_registers.buf_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5549),
    .Q(\rbzero.spi_registers.buf_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5180),
    .Q(\rbzero.spi_registers.buf_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5304),
    .Q(\rbzero.spi_registers.buf_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5362),
    .Q(\rbzero.spi_registers.buf_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(clknet_leaf_27_i_clk),
    .D(net3867),
    .Q(\rbzero.spi_registers.buf_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5134),
    .Q(\rbzero.spi_registers.buf_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(clknet_leaf_13_i_clk),
    .D(net899),
    .Q(\rbzero.spi_registers.buf_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(clknet_leaf_13_i_clk),
    .D(net854),
    .Q(\rbzero.spi_registers.buf_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(clknet_leaf_13_i_clk),
    .D(net825),
    .Q(\rbzero.spi_registers.buf_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21672_ (.CLK(clknet_leaf_13_i_clk),
    .D(net931),
    .Q(\rbzero.spi_registers.buf_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(clknet_leaf_14_i_clk),
    .D(net818),
    .Q(\rbzero.spi_registers.buf_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21674_ (.CLK(clknet_leaf_14_i_clk),
    .D(net808),
    .Q(\rbzero.spi_registers.buf_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(clknet_leaf_14_i_clk),
    .D(net5373),
    .Q(\rbzero.spi_registers.buf_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_14_i_clk),
    .D(net842),
    .Q(\rbzero.spi_registers.buf_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(clknet_leaf_16_i_clk),
    .D(net5016),
    .Q(\rbzero.spi_registers.buf_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_27_i_clk),
    .D(net5188),
    .Q(\rbzero.spi_registers.buf_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_44_i_clk),
    .D(net5081),
    .Q(\rbzero.spi_registers.buf_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5324),
    .Q(\rbzero.spi_registers.buf_mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5285),
    .Q(\rbzero.spi_registers.buf_mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5245),
    .Q(\rbzero.spi_registers.buf_mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_35_i_clk),
    .D(net5281),
    .Q(\rbzero.spi_registers.buf_mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_28_i_clk),
    .D(net5089),
    .Q(\rbzero.spi_registers.buf_texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(clknet_leaf_28_i_clk),
    .D(net5074),
    .Q(\rbzero.spi_registers.buf_texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(clknet_leaf_29_i_clk),
    .D(net5228),
    .Q(\rbzero.spi_registers.buf_texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21687_ (.CLK(clknet_leaf_28_i_clk),
    .D(net5238),
    .Q(\rbzero.spi_registers.buf_texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_29_i_clk),
    .D(net5059),
    .Q(\rbzero.spi_registers.buf_texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5320),
    .Q(\rbzero.spi_registers.buf_texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5199),
    .Q(\rbzero.spi_registers.buf_texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5203),
    .Q(\rbzero.spi_registers.buf_texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(clknet_leaf_26_i_clk),
    .D(net5224),
    .Q(\rbzero.spi_registers.buf_texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(clknet_leaf_25_i_clk),
    .D(net5393),
    .Q(\rbzero.spi_registers.buf_texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(clknet_leaf_3_i_clk),
    .D(net5032),
    .Q(\rbzero.spi_registers.buf_texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(clknet_leaf_2_i_clk),
    .D(net800),
    .Q(\rbzero.spi_registers.buf_texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(clknet_leaf_2_i_clk),
    .D(net970),
    .Q(\rbzero.spi_registers.buf_texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(clknet_leaf_3_i_clk),
    .D(net4117),
    .Q(\rbzero.spi_registers.buf_texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(clknet_leaf_2_i_clk),
    .D(net912),
    .Q(\rbzero.spi_registers.buf_texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21699_ (.CLK(clknet_leaf_5_i_clk),
    .D(net743),
    .Q(\rbzero.spi_registers.buf_texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(clknet_leaf_101_i_clk),
    .D(net5063),
    .Q(\rbzero.spi_registers.buf_texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(clknet_leaf_101_i_clk),
    .D(net4993),
    .Q(\rbzero.spi_registers.buf_texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21702_ (.CLK(clknet_leaf_101_i_clk),
    .D(net862),
    .Q(\rbzero.spi_registers.buf_texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(clknet_leaf_101_i_clk),
    .D(net5163),
    .Q(\rbzero.spi_registers.buf_texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21704_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4609),
    .Q(\rbzero.spi_registers.buf_texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21705_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5036),
    .Q(\rbzero.spi_registers.buf_texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5097),
    .Q(\rbzero.spi_registers.buf_texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(clknet_leaf_20_i_clk),
    .D(net5040),
    .Q(\rbzero.spi_registers.buf_texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21708_ (.CLK(clknet_leaf_19_i_clk),
    .D(net1705),
    .Q(\rbzero.spi_registers.buf_texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21709_ (.CLK(clknet_leaf_19_i_clk),
    .D(net1654),
    .Q(\rbzero.spi_registers.buf_texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21710_ (.CLK(clknet_leaf_19_i_clk),
    .D(net2078),
    .Q(\rbzero.spi_registers.buf_texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21711_ (.CLK(clknet_leaf_26_i_clk),
    .D(net1669),
    .Q(\rbzero.spi_registers.buf_texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21712_ (.CLK(clknet_leaf_25_i_clk),
    .D(net1831),
    .Q(\rbzero.spi_registers.buf_texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21713_ (.CLK(clknet_leaf_26_i_clk),
    .D(net1606),
    .Q(\rbzero.spi_registers.buf_texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21714_ (.CLK(clknet_leaf_25_i_clk),
    .D(net2276),
    .Q(\rbzero.spi_registers.buf_texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21715_ (.CLK(clknet_leaf_17_i_clk),
    .D(net2092),
    .Q(\rbzero.spi_registers.buf_texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21716_ (.CLK(clknet_leaf_26_i_clk),
    .D(net2258),
    .Q(\rbzero.spi_registers.buf_texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21717_ (.CLK(clknet_leaf_17_i_clk),
    .D(net1914),
    .Q(\rbzero.spi_registers.buf_texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21718_ (.CLK(clknet_leaf_8_i_clk),
    .D(net3013),
    .Q(\rbzero.spi_registers.buf_texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1649),
    .Q(\rbzero.spi_registers.buf_texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21720_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1627),
    .Q(\rbzero.spi_registers.buf_texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21721_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1694),
    .Q(\rbzero.spi_registers.buf_texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21722_ (.CLK(clknet_leaf_8_i_clk),
    .D(net2595),
    .Q(\rbzero.spi_registers.buf_texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(clknet_leaf_4_i_clk),
    .D(net2489),
    .Q(\rbzero.spi_registers.buf_texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21724_ (.CLK(clknet_leaf_4_i_clk),
    .D(net4226),
    .Q(\rbzero.spi_registers.buf_texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21725_ (.CLK(clknet_leaf_2_i_clk),
    .D(net6031),
    .Q(\rbzero.spi_registers.buf_texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21726_ (.CLK(clknet_leaf_2_i_clk),
    .D(net1731),
    .Q(\rbzero.spi_registers.buf_texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21727_ (.CLK(clknet_leaf_2_i_clk),
    .D(net6106),
    .Q(\rbzero.spi_registers.buf_texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_2_i_clk),
    .D(net1702),
    .Q(\rbzero.spi_registers.buf_texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1714),
    .Q(\rbzero.spi_registers.buf_texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1672),
    .Q(\rbzero.spi_registers.buf_texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1550),
    .Q(\rbzero.spi_registers.buf_texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(clknet_leaf_22_i_clk),
    .D(net5731),
    .Q(\rbzero.spi_registers.buf_texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21733_ (.CLK(clknet_leaf_22_i_clk),
    .D(net1911),
    .Q(\rbzero.spi_registers.buf_texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21734_ (.CLK(clknet_leaf_22_i_clk),
    .D(net1789),
    .Q(\rbzero.spi_registers.buf_texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1870),
    .Q(\rbzero.spi_registers.buf_texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(clknet_leaf_23_i_clk),
    .D(net2115),
    .Q(\rbzero.spi_registers.buf_texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21737_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1885),
    .Q(\rbzero.spi_registers.buf_texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21738_ (.CLK(clknet_leaf_24_i_clk),
    .D(net2089),
    .Q(\rbzero.spi_registers.buf_texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(clknet_leaf_24_i_clk),
    .D(net2457),
    .Q(\rbzero.spi_registers.buf_texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21740_ (.CLK(clknet_leaf_24_i_clk),
    .D(net2535),
    .Q(\rbzero.spi_registers.buf_texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21741_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1808),
    .Q(\rbzero.spi_registers.buf_texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(clknet_leaf_21_i_clk),
    .D(net4260),
    .Q(\rbzero.spi_registers.buf_texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4238),
    .Q(\rbzero.spi_registers.buf_texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(clknet_leaf_1_i_clk),
    .D(net617),
    .Q(\rbzero.spi_registers.buf_texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21745_ (.CLK(clknet_leaf_0_i_clk),
    .D(net2096),
    .Q(\rbzero.spi_registers.buf_texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21746_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1565),
    .Q(\rbzero.spi_registers.buf_texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21747_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1547),
    .Q(\rbzero.spi_registers.buf_texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1786),
    .Q(\rbzero.spi_registers.buf_texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(clknet_leaf_102_i_clk),
    .D(net1646),
    .Q(\rbzero.spi_registers.buf_texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(clknet_leaf_102_i_clk),
    .D(net2022),
    .Q(\rbzero.spi_registers.buf_texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(clknet_leaf_0_i_clk),
    .D(net1640),
    .Q(\rbzero.spi_registers.buf_texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4330),
    .Q(\rbzero.spi_registers.buf_texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21753_ (.CLK(clknet_leaf_21_i_clk),
    .D(net1576),
    .Q(\rbzero.spi_registers.buf_texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(clknet_leaf_21_i_clk),
    .D(net2356),
    .Q(\rbzero.spi_registers.buf_texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21755_ (.CLK(clknet_leaf_22_i_clk),
    .D(net5765),
    .Q(\rbzero.spi_registers.buf_texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(clknet_leaf_22_i_clk),
    .D(net1561),
    .Q(\rbzero.spi_registers.buf_texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(clknet_leaf_22_i_clk),
    .D(net1905),
    .Q(\rbzero.spi_registers.buf_texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1711),
    .Q(\rbzero.spi_registers.buf_texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1688),
    .Q(\rbzero.spi_registers.buf_texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1873),
    .Q(\rbzero.spi_registers.buf_texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_23_i_clk),
    .D(net1663),
    .Q(\rbzero.spi_registers.buf_texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(clknet_leaf_24_i_clk),
    .D(net1966),
    .Q(\rbzero.spi_registers.buf_texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(clknet_leaf_25_i_clk),
    .D(net6166),
    .Q(\rbzero.spi_registers.buf_texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(clknet_leaf_25_i_clk),
    .D(net6174),
    .Q(\rbzero.spi_registers.buf_texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(clknet_leaf_20_i_clk),
    .D(net1746),
    .Q(\rbzero.spi_registers.buf_texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21766_ (.CLK(clknet_leaf_18_i_clk),
    .D(net5840),
    .Q(\rbzero.spi_registers.buf_texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21767_ (.CLK(clknet_leaf_8_i_clk),
    .D(net2016),
    .Q(\rbzero.spi_registers.buf_texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1991),
    .Q(\rbzero.spi_registers.buf_texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21769_ (.CLK(clknet_leaf_4_i_clk),
    .D(net1720),
    .Q(\rbzero.spi_registers.buf_texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(clknet_leaf_4_i_clk),
    .D(net2157),
    .Q(\rbzero.spi_registers.buf_texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1545),
    .Q(\rbzero.spi_registers.buf_texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(clknet_leaf_5_i_clk),
    .D(net1568),
    .Q(\rbzero.spi_registers.buf_texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(clknet_leaf_102_i_clk),
    .D(net1846),
    .Q(\rbzero.spi_registers.buf_texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_102_i_clk),
    .D(net1849),
    .Q(\rbzero.spi_registers.buf_texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(clknet_leaf_2_i_clk),
    .D(net1633),
    .Q(\rbzero.spi_registers.buf_texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21776_ (.CLK(clknet_leaf_1_i_clk),
    .D(net4324),
    .Q(\rbzero.spi_registers.buf_texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21777_ (.CLK(clknet_leaf_20_i_clk),
    .D(net2232),
    .Q(\rbzero.spi_registers.buf_texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(clknet_leaf_20_i_clk),
    .D(net2284),
    .Q(\rbzero.spi_registers.buf_texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(clknet_leaf_20_i_clk),
    .D(net6035),
    .Q(\rbzero.spi_registers.buf_texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_30_i_clk),
    .D(net3154),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21781_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00950_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3963),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(clknet_leaf_31_i_clk),
    .D(net3928),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00953_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_93_i_clk),
    .D(net626),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(clknet_leaf_10_i_clk),
    .D(net4337),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21787_ (.CLK(clknet_leaf_11_i_clk),
    .D(net4308),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(clknet_leaf_11_i_clk),
    .D(net5465),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(clknet_leaf_11_i_clk),
    .D(net4340),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(clknet_leaf_11_i_clk),
    .D(net6012),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(clknet_leaf_11_i_clk),
    .D(net4302),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(clknet_leaf_11_i_clk),
    .D(net2930),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21793_ (.CLK(clknet_leaf_11_i_clk),
    .D(net3002),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21794_ (.CLK(clknet_leaf_11_i_clk),
    .D(net4221),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(clknet_leaf_12_i_clk),
    .D(net6157),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21796_ (.CLK(clknet_leaf_12_i_clk),
    .D(net2815),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(clknet_leaf_11_i_clk),
    .D(net6184),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(clknet_leaf_11_i_clk),
    .D(net727),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21799_ (.CLK(clknet_leaf_12_i_clk),
    .D(net1037),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21800_ (.CLK(clknet_leaf_12_i_clk),
    .D(net3160),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(clknet_leaf_89_i_clk),
    .D(net4357),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(clknet_leaf_89_i_clk),
    .D(net2838),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(clknet_leaf_89_i_clk),
    .D(net4895),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(clknet_leaf_89_i_clk),
    .D(net2924),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(clknet_leaf_89_i_clk),
    .D(net4296),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(clknet_leaf_90_i_clk),
    .D(net2891),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(clknet_leaf_10_i_clk),
    .D(net6193),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(clknet_leaf_90_i_clk),
    .D(net4360),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(clknet_leaf_10_i_clk),
    .D(net4290),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(clknet_leaf_10_i_clk),
    .D(net2894),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(clknet_leaf_10_i_clk),
    .D(net4677),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(clknet_leaf_10_i_clk),
    .D(net4389),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(clknet_leaf_10_i_clk),
    .D(net6215),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(clknet_leaf_9_i_clk),
    .D(net3084),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(clknet_leaf_9_i_clk),
    .D(net3955),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21816_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4633),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21817_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4366),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4445),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4523),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21820_ (.CLK(clknet_leaf_87_i_clk),
    .D(net3875),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(clknet_leaf_87_i_clk),
    .D(net3850),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(clknet_leaf_91_i_clk),
    .D(net3142),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21823_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4647),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(clknet_leaf_87_i_clk),
    .D(net3789),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4564),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4409),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(clknet_leaf_88_i_clk),
    .D(net3903),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21828_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4517),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(clknet_leaf_88_i_clk),
    .D(net3832),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(clknet_leaf_89_i_clk),
    .D(net3746),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(clknet_leaf_87_i_clk),
    .D(net3658),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(clknet_leaf_96_i_clk),
    .D(net4415),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21833_ (.CLK(clknet_leaf_91_i_clk),
    .D(net4421),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(clknet_leaf_88_i_clk),
    .D(net3771),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(clknet_leaf_83_i_clk),
    .D(net4603),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(clknet_leaf_83_i_clk),
    .D(net3860),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(clknet_leaf_83_i_clk),
    .D(net3879),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(clknet_leaf_81_i_clk),
    .D(net3546),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4778),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(clknet_leaf_81_i_clk),
    .D(net4449),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(clknet_leaf_81_i_clk),
    .D(net950),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(clknet_leaf_80_i_clk),
    .D(net3841),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(clknet_leaf_81_i_clk),
    .D(net3178),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(clknet_leaf_81_i_clk),
    .D(net1252),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(clknet_leaf_82_i_clk),
    .D(net3245),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(clknet_leaf_82_i_clk),
    .D(net1367),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(clknet_leaf_82_i_clk),
    .D(net1227),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21848_ (.CLK(clknet_leaf_83_i_clk),
    .D(net1441),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(clknet_leaf_81_i_clk),
    .D(net4617),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(clknet_leaf_81_i_clk),
    .D(net4731),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(clknet_leaf_98_i_clk),
    .D(net4643),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(clknet_leaf_81_i_clk),
    .D(net3677),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(clknet_leaf_81_i_clk),
    .D(net3618),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(clknet_leaf_82_i_clk),
    .D(net3810),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(clknet_leaf_97_i_clk),
    .D(net4462),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(clknet_leaf_82_i_clk),
    .D(net3703),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(clknet_leaf_82_i_clk),
    .D(net4750),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(clknet_leaf_97_i_clk),
    .D(net4637),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(clknet_leaf_83_i_clk),
    .D(net2901),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(clknet_leaf_94_i_clk),
    .D(net3228),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(clknet_leaf_94_i_clk),
    .D(net2631),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(clknet_leaf_94_i_clk),
    .D(net1602),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(clknet_leaf_94_i_clk),
    .D(net3331),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(clknet_leaf_94_i_clk),
    .D(net3828),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(clknet_leaf_94_i_clk),
    .D(net3564),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(clknet_leaf_6_i_clk),
    .D(net4970),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(clknet_leaf_100_i_clk),
    .D(net955),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(clknet_leaf_100_i_clk),
    .D(net1238),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(clknet_leaf_100_i_clk),
    .D(net1171),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(clknet_leaf_100_i_clk),
    .D(net1329),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(clknet_leaf_100_i_clk),
    .D(net1244),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(clknet_leaf_100_i_clk),
    .D(net1205),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(clknet_leaf_95_i_clk),
    .D(net5253),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1223),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1126),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1246),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1225),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1287),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(clknet_leaf_99_i_clk),
    .D(net1231),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(clknet_leaf_99_i_clk),
    .D(net1178),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(clknet_leaf_99_i_clk),
    .D(net1169),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(clknet_leaf_99_i_clk),
    .D(net1163),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(clknet_leaf_99_i_clk),
    .D(net5502),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1277),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(clknet_leaf_98_i_clk),
    .D(net5542),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(clknet_leaf_98_i_clk),
    .D(net1390),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1281),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(clknet_leaf_97_i_clk),
    .D(net1273),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(clknet_leaf_96_i_clk),
    .D(net1289),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(clknet_leaf_96_i_clk),
    .D(net1264),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(clknet_leaf_96_i_clk),
    .D(net1293),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(clknet_leaf_96_i_clk),
    .D(net1340),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1336),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1410),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1439),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1471),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1382),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1279),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(clknet_leaf_95_i_clk),
    .D(net5051),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(clknet_leaf_95_i_clk),
    .D(net1434),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(clknet_leaf_94_i_clk),
    .D(net1511),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1315),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1371),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1342),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1476),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1414),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(clknet_leaf_92_i_clk),
    .D(net1492),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(clknet_leaf_92_i_clk),
    .D(net5389),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(clknet_leaf_92_i_clk),
    .D(net5385),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(clknet_leaf_90_i_clk),
    .D(net5214),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21911_ (.CLK(clknet_leaf_90_i_clk),
    .D(net5195),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(clknet_leaf_90_i_clk),
    .D(net1271),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(clknet_leaf_90_i_clk),
    .D(net5207),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(clknet_leaf_90_i_clk),
    .D(net1325),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(clknet_leaf_92_i_clk),
    .D(net1240),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(clknet_leaf_92_i_clk),
    .D(net1494),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(clknet_leaf_92_i_clk),
    .D(net1344),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1396),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1307),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1338),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(clknet_leaf_93_i_clk),
    .D(net1401),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1363),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1323),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1317),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1266),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1248),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1176),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1283),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1254),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(clknet_leaf_8_i_clk),
    .D(net4835),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1484),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(clknet_leaf_8_i_clk),
    .D(net4842),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(clknet_leaf_8_i_clk),
    .D(net1242),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1200),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1361),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1412),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(clknet_leaf_7_i_clk),
    .D(net1221),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(clknet_leaf_9_i_clk),
    .D(net1303),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(clknet_leaf_9_i_clk),
    .D(net4870),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(clknet_leaf_9_i_clk),
    .D(net4863),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(net166),
    .D(net1523),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(net167),
    .D(net2652),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(net168),
    .D(net2372),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(net169),
    .D(net1805),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(net170),
    .D(net2795),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(net171),
    .D(net1359),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21947_ (.CLK(net172),
    .D(net2410),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(net173),
    .D(net2217),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(net174),
    .D(net1622),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(net175),
    .D(net730),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(net176),
    .D(net2694),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(net177),
    .D(net2811),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(net178),
    .D(net2736),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(net179),
    .D(net1949),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(net180),
    .D(net2610),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(net181),
    .D(net2818),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(net182),
    .D(net2270),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(net183),
    .D(net2513),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(net184),
    .D(net2658),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(net185),
    .D(net1033),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(net186),
    .D(net2205),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(net187),
    .D(net2713),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(net188),
    .D(net2032),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(net189),
    .D(net2483),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(net190),
    .D(net2806),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(net191),
    .D(net1444),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(net192),
    .D(net2279),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(net193),
    .D(net2432),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(net194),
    .D(net2297),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(net195),
    .D(net1419),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(net196),
    .D(net1896),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(net197),
    .D(net2621),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(net198),
    .D(net2029),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(net199),
    .D(net2333),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(net200),
    .D(net1499),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(net201),
    .D(net2053),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(net202),
    .D(net2075),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(net203),
    .D(net2583),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(net204),
    .D(net2401),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(net205),
    .D(net1198),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(net206),
    .D(net1826),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(net207),
    .D(net2392),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(net208),
    .D(net2532),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(net209),
    .D(net2318),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(net210),
    .D(net1755),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(net211),
    .D(net1388),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(net212),
    .D(net1963),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(net213),
    .D(net2504),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(net214),
    .D(net2348),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(net215),
    .D(net1104),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(net216),
    .D(net1817),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(net217),
    .D(net2801),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(net218),
    .D(net1740),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(net219),
    .D(net2148),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(net220),
    .D(net2615),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(net221),
    .D(net2162),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(net222),
    .D(net2291),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(net223),
    .D(net1969),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(net224),
    .D(net1972),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(net225),
    .D(net1463),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(net226),
    .D(net1908),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(net227),
    .D(net2417),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(net228),
    .D(net1931),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(net229),
    .D(net2036),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(clknet_leaf_10_i_clk),
    .D(net5469),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3271),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(clknet_leaf_100_i_clk),
    .D(net3644),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(clknet_leaf_100_i_clk),
    .D(net3593),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(clknet_leaf_100_i_clk),
    .D(net3820),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(clknet_leaf_100_i_clk),
    .D(net3740),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3192),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3431),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(clknet_leaf_97_i_clk),
    .D(net3639),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(clknet_leaf_97_i_clk),
    .D(net3588),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3320),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3687),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3609),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3663),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3469),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(clknet_leaf_81_i_clk),
    .D(net3391),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3456),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(clknet_leaf_99_i_clk),
    .D(net3350),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3326),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(clknet_leaf_98_i_clk),
    .D(net3232),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(clknet_leaf_97_i_clk),
    .D(net3452),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(clknet_leaf_97_i_clk),
    .D(net3355),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3294),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3759),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3299),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3731),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3846),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3550),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3560),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(clknet_leaf_96_i_clk),
    .D(net3654),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3836),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3785),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3767),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3712),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(clknet_leaf_95_i_clk),
    .D(net3698),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3425),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3415),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3668),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3522),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3778),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(clknet_leaf_92_i_clk),
    .D(net3533),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(clknet_leaf_91_i_clk),
    .D(net3340),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(clknet_leaf_91_i_clk),
    .D(net3308),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(clknet_leaf_91_i_clk),
    .D(net3304),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(clknet_leaf_91_i_clk),
    .D(net3443),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3368),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3576),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22052_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3716),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3614),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3278),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22055_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3583),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3345),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(clknet_leaf_90_i_clk),
    .D(net3438),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22058_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3803),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(clknet_leaf_10_i_clk),
    .D(net3363),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3289),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3601),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3649),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3571),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3486),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3491),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(clknet_leaf_7_i_clk),
    .D(net3479),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(clknet_leaf_8_i_clk),
    .D(net3261),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22068_ (.CLK(clknet_leaf_8_i_clk),
    .D(net3708),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(clknet_leaf_8_i_clk),
    .D(net3735),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(clknet_leaf_13_i_clk),
    .D(net3815),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(clknet_leaf_13_i_clk),
    .D(net3755),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(clknet_leaf_8_i_clk),
    .D(net3673),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(clknet_leaf_9_i_clk),
    .D(net3682),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _22074_ (.CLK(clknet_leaf_13_i_clk),
    .D(net3517),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _22075_ (.CLK(clknet_leaf_13_i_clk),
    .D(net3499),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _22076_ (.CLK(clknet_leaf_9_i_clk),
    .D(net3386),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _22077_ (.CLK(clknet_leaf_9_i_clk),
    .D(net3527),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _22078_ (.CLK(clknet_leaf_13_i_clk),
    .D(net3313),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _22079_ (.CLK(clknet_leaf_13_i_clk),
    .D(net3253),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _22080_ (.CLK(clknet_leaf_6_i_clk),
    .D(net6178),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _22081_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01250_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22082_ (.CLK(clknet_leaf_79_i_clk),
    .D(net1109),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _22083_ (.CLK(clknet_leaf_49_i_clk),
    .D(net1452),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _22084_ (.CLK(clknet_leaf_47_i_clk),
    .D(net6027),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_1 _22085_ (.CLK(clknet_leaf_74_i_clk),
    .D(net4019),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22086_ (.CLK(clknet_leaf_73_i_clk),
    .D(net3967),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22087_ (.CLK(clknet_leaf_74_i_clk),
    .D(net4024),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22088_ (.CLK(clknet_leaf_49_i_clk),
    .D(net3899),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22089_ (.CLK(clknet_leaf_48_i_clk),
    .D(net4035),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22090_ (.CLK(clknet_leaf_48_i_clk),
    .D(_01259_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22091_ (.CLK(clknet_leaf_47_i_clk),
    .D(net4062),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22092_ (.CLK(clknet_leaf_49_i_clk),
    .D(net4003),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22093_ (.CLK(clknet_leaf_49_i_clk),
    .D(net3931),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22094_ (.CLK(clknet_leaf_49_i_clk),
    .D(net3938),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22095_ (.CLK(clknet_leaf_6_i_clk),
    .D(_01264_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22096_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1174),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22097_ (.CLK(clknet_leaf_6_i_clk),
    .D(net1579),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22098_ (.CLK(net230),
    .D(net1482),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22099_ (.CLK(net231),
    .D(net2039),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22100_ (.CLK(net232),
    .D(net1876),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22101_ (.CLK(net233),
    .D(net2106),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22102_ (.CLK(net234),
    .D(net2438),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22103_ (.CLK(net235),
    .D(net762),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22104_ (.CLK(net236),
    .D(net2655),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22105_ (.CLK(net237),
    .D(net2607),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22106_ (.CLK(net238),
    .D(net2321),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22107_ (.CLK(net239),
    .D(net2860),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22108_ (.CLK(net240),
    .D(net2786),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22109_ (.CLK(net241),
    .D(net2883),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22110_ (.CLK(net242),
    .D(net2342),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22111_ (.CLK(net243),
    .D(net2586),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22112_ (.CLK(net244),
    .D(net2868),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22113_ (.CLK(net245),
    .D(net1090),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22114_ (.CLK(net246),
    .D(net1802),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22115_ (.CLK(net247),
    .D(net1882),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22116_ (.CLK(net248),
    .D(net1840),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22117_ (.CLK(net249),
    .D(net2168),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22118_ (.CLK(net250),
    .D(net2798),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22119_ (.CLK(net251),
    .D(net1437),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22120_ (.CLK(net252),
    .D(net2414),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22121_ (.CLK(net253),
    .D(net2181),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22122_ (.CLK(net254),
    .D(net2184),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22123_ (.CLK(net255),
    .D(net1385),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22124_ (.CLK(net256),
    .D(net2199),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22125_ (.CLK(net257),
    .D(net2121),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22126_ (.CLK(net258),
    .D(net2466),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22127_ (.CLK(net259),
    .D(net2187),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22128_ (.CLK(net260),
    .D(net2510),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22129_ (.CLK(net261),
    .D(net1399),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22130_ (.CLK(net262),
    .D(net1811),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22131_ (.CLK(net263),
    .D(net2208),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22132_ (.CLK(net264),
    .D(net2229),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22133_ (.CLK(net265),
    .D(net1236),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22134_ (.CLK(net266),
    .D(net2589),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22135_ (.CLK(net267),
    .D(net2598),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22136_ (.CLK(net268),
    .D(net1758),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22137_ (.CLK(net269),
    .D(net2175),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22138_ (.CLK(net270),
    .D(net1925),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22139_ (.CLK(net271),
    .D(net1858),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22140_ (.CLK(net272),
    .D(net2178),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22141_ (.CLK(net273),
    .D(net2190),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22142_ (.CLK(net274),
    .D(net1374),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22143_ (.CLK(net275),
    .D(net1140),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22144_ (.CLK(net276),
    .D(net2202),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22145_ (.CLK(net277),
    .D(net2546),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22146_ (.CLK(net278),
    .D(net2287),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22147_ (.CLK(net279),
    .D(net2324),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22148_ (.CLK(net280),
    .D(net2251),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22149_ (.CLK(net281),
    .D(net2435),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22150_ (.CLK(net282),
    .D(net2745),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22151_ (.CLK(net283),
    .D(net2151),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22152_ (.CLK(net284),
    .D(net1487),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22153_ (.CLK(net285),
    .D(net1269),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22154_ (.CLK(net286),
    .D(net2580),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22155_ (.CLK(net287),
    .D(net2567),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22156_ (.CLK(net288),
    .D(net2214),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22157_ (.CLK(net289),
    .D(net2142),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22158_ (.CLK(net290),
    .D(net1834),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22159_ (.CLK(net291),
    .D(net1520),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22160_ (.CLK(net292),
    .D(net2245),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22161_ (.CLK(net293),
    .D(net2451),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22162_ (.CLK(net294),
    .D(net2193),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22163_ (.CLK(net295),
    .D(net752),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22164_ (.CLK(net296),
    .D(net1612),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22165_ (.CLK(net297),
    .D(net2351),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22166_ (.CLK(net298),
    .D(net1928),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22167_ (.CLK(net299),
    .D(net2618),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22168_ (.CLK(net300),
    .D(net1796),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22169_ (.CLK(net301),
    .D(net2523),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22170_ (.CLK(net302),
    .D(net1717),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22171_ (.CLK(net303),
    .D(net2118),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22172_ (.CLK(net304),
    .D(net1752),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22173_ (.CLK(net305),
    .D(net1075),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22174_ (.CLK(net306),
    .D(net1890),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22175_ (.CLK(net307),
    .D(net1987),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22176_ (.CLK(net308),
    .D(net2273),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22177_ (.CLK(net309),
    .D(net1937),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22178_ (.CLK(net310),
    .D(net1852),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22179_ (.CLK(net311),
    .D(net2667),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22180_ (.CLK(net312),
    .D(net2719),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22181_ (.CLK(net313),
    .D(net1919),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22182_ (.CLK(net314),
    .D(net2742),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22183_ (.CLK(net315),
    .D(net1095),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22184_ (.CLK(net316),
    .D(net1676),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22185_ (.CLK(net317),
    .D(net2362),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22186_ (.CLK(net318),
    .D(net2130),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22187_ (.CLK(net319),
    .D(net1946),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22188_ (.CLK(net320),
    .D(net2529),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22189_ (.CLK(net321),
    .D(net1334),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22190_ (.CLK(net322),
    .D(net2050),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22191_ (.CLK(net323),
    .D(net2404),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22192_ (.CLK(net324),
    .D(net2315),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22193_ (.CLK(net325),
    .D(net635),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22194_ (.CLK(net326),
    .D(net2026),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22195_ (.CLK(net327),
    .D(net1958),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22196_ (.CLK(net328),
    .D(net1940),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22197_ (.CLK(net329),
    .D(net2239),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22198_ (.CLK(net330),
    .D(net1879),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22199_ (.CLK(net331),
    .D(net2872),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22200_ (.CLK(net332),
    .D(net1814),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22201_ (.CLK(net333),
    .D(net2426),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22202_ (.CLK(net334),
    .D(net1767),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22203_ (.CLK(net335),
    .D(net1193),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22204_ (.CLK(net336),
    .D(net2220),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22205_ (.CLK(net337),
    .D(net2267),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22206_ (.CLK(net338),
    .D(net2540),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22207_ (.CLK(net339),
    .D(net2552),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22208_ (.CLK(net340),
    .D(net1643),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22209_ (.CLK(net341),
    .D(net2664),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22210_ (.CLK(net342),
    .D(net1660),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22211_ (.CLK(net343),
    .D(net1997),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22212_ (.CLK(net344),
    .D(net1952),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22213_ (.CLK(net345),
    .D(net1112),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22214_ (.CLK(net346),
    .D(net1899),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22215_ (.CLK(net347),
    .D(net2899),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22216_ (.CLK(net348),
    .D(net1799),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22217_ (.CLK(net349),
    .D(net2661),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22218_ (.CLK(net350),
    .D(net1528),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22219_ (.CLK(net351),
    .D(net2441),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22220_ (.CLK(net352),
    .D(net2303),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22221_ (.CLK(net353),
    .D(net2133),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22222_ (.CLK(net354),
    .D(net2673),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22223_ (.CLK(net355),
    .D(net1447),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22224_ (.CLK(net356),
    .D(net1984),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22225_ (.CLK(net357),
    .D(net2773),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22226_ (.CLK(net358),
    .D(net1503),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22227_ (.CLK(net359),
    .D(net2444),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22228_ (.CLK(net360),
    .D(net2099),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22229_ (.CLK(net361),
    .D(net1981),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22230_ (.CLK(net362),
    .D(net2327),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22231_ (.CLK(net363),
    .D(net2601),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22232_ (.CLK(net364),
    .D(net2516),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22233_ (.CLK(net365),
    .D(net830),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22234_ (.CLK(net366),
    .D(net2480),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22235_ (.CLK(net367),
    .D(net2549),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22236_ (.CLK(net368),
    .D(net2878),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22237_ (.CLK(net369),
    .D(net1517),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22238_ (.CLK(net370),
    .D(net1743),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22239_ (.CLK(net371),
    .D(net2006),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22240_ (.CLK(net372),
    .D(net1708),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22241_ (.CLK(net373),
    .D(net2136),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22242_ (.CLK(net374),
    .D(net1773),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22243_ (.CLK(net375),
    .D(net1203),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22244_ (.CLK(net376),
    .D(net2359),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22245_ (.CLK(net377),
    .D(net2242),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22246_ (.CLK(net378),
    .D(net2640),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22247_ (.CLK(net379),
    .D(net2526),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22248_ (.CLK(net380),
    .D(net2767),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22249_ (.CLK(net381),
    .D(net1429),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22250_ (.CLK(net382),
    .D(net1823),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22251_ (.CLK(net383),
    .D(net1867),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22252_ (.CLK(net384),
    .D(net2492),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22253_ (.CLK(net385),
    .D(net1208),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22254_ (.CLK(net386),
    .D(net1699),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22255_ (.CLK(net387),
    .D(net1682),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22256_ (.CLK(net388),
    .D(net2236),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22257_ (.CLK(net389),
    .D(net2003),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22258_ (.CLK(net390),
    .D(net1782),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22259_ (.CLK(net391),
    .D(net2127),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22260_ (.CLK(net392),
    .D(net1514),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22261_ (.CLK(net393),
    .D(net2047),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22262_ (.CLK(net394),
    .D(net2739),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22263_ (.CLK(net395),
    .D(net1063),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22264_ (.CLK(net396),
    .D(net2676),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22265_ (.CLK(net397),
    .D(net2312),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22266_ (.CLK(net398),
    .D(net2832),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22267_ (.CLK(net399),
    .D(net2019),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22268_ (.CLK(net400),
    .D(net2211),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22269_ (.CLK(net401),
    .D(net2463),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22270_ (.CLK(net402),
    .D(net2710),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22271_ (.CLK(net403),
    .D(net2398),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22272_ (.CLK(net404),
    .D(net1943),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22273_ (.CLK(net405),
    .D(net934),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22274_ (.CLK(net406),
    .D(net2255),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22275_ (.CLK(net407),
    .D(net2248),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22276_ (.CLK(net408),
    .D(net2764),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22277_ (.CLK(net409),
    .D(net2634),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22278_ (.CLK(net410),
    .D(net1556),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22279_ (.CLK(net411),
    .D(net2336),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22280_ (.CLK(net412),
    .D(net2454),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22281_ (.CLK(net413),
    .D(net2498),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22282_ (.CLK(net414),
    .D(net2863),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22283_ (.CLK(net415),
    .D(net1122),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22284_ (.CLK(net416),
    .D(net2627),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22285_ (.CLK(net417),
    .D(net2783),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22286_ (.CLK(net418),
    .D(net2059),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22287_ (.CLK(net419),
    .D(net2112),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22288_ (.CLK(net420),
    .D(net2722),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22289_ (.CLK(net421),
    .D(net2749),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22290_ (.CLK(net422),
    .D(net1490),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22291_ (.CLK(net423),
    .D(net2564),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22292_ (.CLK(net424),
    .D(net2165),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22293_ (.CLK(net425),
    .D(net2716),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22294_ (.CLK(net426),
    .D(net2387),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22295_ (.CLK(net427),
    .D(net2684),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22296_ (.CLK(net428),
    .D(net2697),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22297_ (.CLK(net429),
    .D(net2294),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22298_ (.CLK(net430),
    .D(net2109),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22299_ (.CLK(net431),
    .D(net1432),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22300_ (.CLK(net432),
    .D(net2145),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22301_ (.CLK(net433),
    .D(net2460),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22302_ (.CLK(net434),
    .D(net2065),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22303_ (.CLK(net435),
    .D(net1260),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22304_ (.CLK(net436),
    .D(net1975),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22305_ (.CLK(net437),
    .D(net2012),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22306_ (.CLK(net438),
    .D(net2042),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22307_ (.CLK(net439),
    .D(net2561),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22308_ (.CLK(net440),
    .D(net1479),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22309_ (.CLK(net441),
    .D(net2378),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22310_ (.CLK(net442),
    .D(net1843),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22311_ (.CLK(net443),
    .D(net2477),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22312_ (.CLK(net444),
    .D(net1779),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22313_ (.CLK(net445),
    .D(net1161),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22314_ (.CLK(net446),
    .D(net2056),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22315_ (.CLK(net447),
    .D(net2853),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22316_ (.CLK(net448),
    .D(net2904),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22317_ (.CLK(net449),
    .D(net1666),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22318_ (.CLK(net450),
    .D(net1761),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22319_ (.CLK(net451),
    .D(net2062),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22320_ (.CLK(net452),
    .D(net2670),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22321_ (.CLK(net453),
    .D(net2643),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22322_ (.CLK(net454),
    .D(net2447),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22323_ (.CLK(net455),
    .D(net1155),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22324_ (.CLK(net456),
    .D(net2847),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22325_ (.CLK(net457),
    .D(net2646),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22326_ (.CLK(net458),
    .D(net1820),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22327_ (.CLK(net459),
    .D(net2309),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22328_ (.CLK(net460),
    .D(net1553),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22329_ (.CLK(net461),
    .D(net2761),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22330_ (.CLK(net462),
    .D(net1679),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22331_ (.CLK(net463),
    .D(net2423),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22332_ (.CLK(net464),
    .D(net2306),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22333_ (.CLK(net465),
    .D(net1354),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22334_ (.CLK(net466),
    .D(net1734),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22335_ (.CLK(net467),
    .D(net2624),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22336_ (.CLK(net468),
    .D(net2171),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22337_ (.CLK(net469),
    .D(net2501),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22338_ (.CLK(net470),
    .D(net1426),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22339_ (.CLK(net471),
    .D(net2691),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22340_ (.CLK(net472),
    .D(net2850),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22341_ (.CLK(net473),
    .D(net1978),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22342_ (.CLK(net474),
    .D(net1725),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22343_ (.CLK(net475),
    .D(net1150),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22344_ (.CLK(net476),
    .D(net2420),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22345_ (.CLK(net477),
    .D(net2758),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22346_ (.CLK(net478),
    .D(net2507),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22347_ (.CLK(net479),
    .D(net2681),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22348_ (.CLK(net480),
    .D(net1474),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22349_ (.CLK(net481),
    .D(net2103),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22350_ (.CLK(net482),
    .D(net1955),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22351_ (.CLK(net483),
    .D(net1934),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22352_ (.CLK(net484),
    .D(net2339),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22353_ (.CLK(net485),
    .D(net2369),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22354_ (.CLK(net486),
    .D(net1455),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22355_ (.CLK(net487),
    .D(net2755),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22356_ (.CLK(net488),
    .D(net2725),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22357_ (.CLK(net489),
    .D(net2395),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22358_ (.CLK(net490),
    .D(net1460),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22359_ (.CLK(net491),
    .D(net2384),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22360_ (.CLK(net492),
    .D(net2081),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22361_ (.CLK(net493),
    .D(net2223),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22362_ (.CLK(net494),
    .D(net1902),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22363_ (.CLK(net495),
    .D(net1349),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22364_ (.CLK(net496),
    .D(net2701),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22365_ (.CLK(net497),
    .D(net2261),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22366_ (.CLK(net498),
    .D(net1685),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22367_ (.CLK(net499),
    .D(net2087),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22368_ (.CLK(net500),
    .D(net2730),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22369_ (.CLK(net501),
    .D(net1450),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22370_ (.CLK(net502),
    .D(net2704),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22371_ (.CLK(net503),
    .D(net2733),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22372_ (.CLK(net504),
    .D(net2829),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22373_ (.CLK(net505),
    .D(net997),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22374_ (.CLK(net506),
    .D(net2009),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22375_ (.CLK(net507),
    .D(net2330),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22376_ (.CLK(net508),
    .D(net1749),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22377_ (.CLK(net509),
    .D(net2375),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22378_ (.CLK(net510),
    .D(net2486),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22379_ (.CLK(net511),
    .D(net2857),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22380_ (.CLK(net512),
    .D(net2780),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22381_ (.CLK(net513),
    .D(net2558),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22382_ (.CLK(net514),
    .D(net2495),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22383_ (.CLK(net515),
    .D(net1181),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22384_ (.CLK(net516),
    .D(net2637),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22385_ (.CLK(net517),
    .D(net1776),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22386_ (.CLK(net518),
    .D(net2345),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22387_ (.CLK(net519),
    .D(net2570),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22388_ (.CLK(net520),
    .D(net1893),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22389_ (.CLK(net521),
    .D(net2520),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22390_ (.CLK(net522),
    .D(net2154),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22391_ (.CLK(net523),
    .D(net1994),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22392_ (.CLK(net524),
    .D(net1764),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22393_ (.CLK(net525),
    .D(net590),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22394_ (.CLK(net146),
    .D(net2084),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22395_ (.CLK(net147),
    .D(net2300),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22396_ (.CLK(net148),
    .D(net1855),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22397_ (.CLK(net149),
    .D(net2226),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22398_ (.CLK(net150),
    .D(net1630),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22399_ (.CLK(net151),
    .D(net2381),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22400_ (.CLK(net152),
    .D(net2407),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22401_ (.CLK(net153),
    .D(net2471),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22402_ (.CLK(net154),
    .D(net2068),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22403_ (.CLK(net155),
    .D(net1042),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22404_ (.CLK(net156),
    .D(net2139),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22405_ (.CLK(net157),
    .D(net2604),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22406_ (.CLK(net158),
    .D(net2365),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22407_ (.CLK(net159),
    .D(net2573),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22408_ (.CLK(net160),
    .D(net2752),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22409_ (.CLK(net161),
    .D(net2822),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22410_ (.CLK(net162),
    .D(net2576),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22411_ (.CLK(net163),
    .D(net2474),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22412_ (.CLK(net164),
    .D(net2429),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22413_ (.CLK(net165),
    .D(net1466),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22414_ (.CLK(net142),
    .D(net1837),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22415_ (.CLK(net143),
    .D(net2264),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22416_ (.CLK(net144),
    .D(net2649),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22417_ (.CLK(net145),
    .D(net2688),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22418_ (.CLK(clknet_leaf_66_i_clk),
    .D(net667),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22419_ (.CLK(clknet_leaf_66_i_clk),
    .D(net1082),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22420_ (.CLK(clknet_leaf_57_i_clk),
    .D(net4989),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _22421_ (.CLK(clknet_leaf_57_i_clk),
    .D(net4977),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _22422_ (.CLK(clknet_leaf_55_i_clk),
    .D(net5273),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22423_ (.CLK(clknet_leaf_55_i_clk),
    .D(net5336),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22424_ (.CLK(clknet_leaf_54_i_clk),
    .D(net5170),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22425_ (.CLK(clknet_leaf_50_i_clk),
    .D(net5426),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22426_ (.CLK(clknet_leaf_50_i_clk),
    .D(net5457),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _22427_ (.CLK(clknet_leaf_46_i_clk),
    .D(net4765),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _22428_ (.CLK(clknet_leaf_46_i_clk),
    .D(net4738),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _22429_ (.CLK(clknet_leaf_41_i_clk),
    .D(net4397),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _22430_ (.CLK(clknet_leaf_41_i_clk),
    .D(net4548),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _22431_ (.CLK(clknet_leaf_41_i_clk),
    .D(net4505),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22432_ (.CLK(clknet_leaf_40_i_clk),
    .D(net4544),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22433_ (.CLK(clknet_leaf_40_i_clk),
    .D(net4703),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22434_ (.CLK(clknet_leaf_40_i_clk),
    .D(net4940),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22435_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4471),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22436_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4651),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22437_ (.CLK(clknet_leaf_38_i_clk),
    .D(net4655),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22438_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4746),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22439_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4742),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22440_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4681),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22441_ (.CLK(clknet_leaf_39_i_clk),
    .D(net4707),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22442_ (.CLK(clknet_leaf_72_i_clk),
    .D(net4031),
    .Q(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22443_ (.CLK(clknet_leaf_72_i_clk),
    .D(net3536),
    .Q(\rbzero.trace_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22444_ (.CLK(clknet_leaf_72_i_clk),
    .D(net2984),
    .Q(\rbzero.trace_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22445_ (.CLK(clknet_leaf_51_i_clk),
    .D(net3982),
    .Q(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22446_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01615_),
    .Q(\reg_gpout[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22447_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01616_),
    .Q(\reg_gpout[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22448_ (.CLK(clknet_leaf_66_i_clk),
    .D(_01617_),
    .Q(\reg_gpout[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22449_ (.CLK(clknet_leaf_66_i_clk),
    .D(_01618_),
    .Q(\reg_gpout[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22450_ (.CLK(clknet_leaf_66_i_clk),
    .D(_01619_),
    .Q(\reg_gpout[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22451_ (.CLK(clknet_leaf_65_i_clk),
    .D(_01620_),
    .Q(\reg_gpout[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22452_ (.CLK(clknet_leaf_46_i_clk),
    .D(net651),
    .Q(reg_hsync));
 sky130_fd_sc_hd__dfxtp_1 _22453_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01622_),
    .Q(reg_vsync));
 sky130_fd_sc_hd__dfxtp_1 _22454_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01623_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22455_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01624_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22456_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01625_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22457_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01626_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22458_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01627_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22459_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01628_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22460_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01629_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22461_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01630_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22462_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01631_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22463_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01632_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22464_ (.CLK(clknet_leaf_57_i_clk),
    .D(_01633_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22465_ (.CLK(clknet_leaf_69_i_clk),
    .D(net659),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22466_ (.CLK(clknet_leaf_69_i_clk),
    .D(net1129),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22467_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4427),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22468_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4660),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22469_ (.CLK(clknet_leaf_79_i_clk),
    .D(net4808),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22470_ (.CLK(clknet_leaf_79_i_clk),
    .D(net4793),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22471_ (.CLK(clknet_leaf_81_i_clk),
    .D(net4441),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22472_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4624),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22473_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4907),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22474_ (.CLK(clknet_leaf_80_i_clk),
    .D(net4804),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22475_ (.CLK(clknet_leaf_77_i_clk),
    .D(net661),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22476_ (.CLK(clknet_3_5_0_i_clk),
    .D(net1922),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22477_ (.CLK(clknet_leaf_77_i_clk),
    .D(net655),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22478_ (.CLK(clknet_leaf_77_i_clk),
    .D(net1184),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22479_ (.CLK(clknet_leaf_67_i_clk),
    .D(net665),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22480_ (.CLK(clknet_leaf_67_i_clk),
    .D(net1137),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22481_ (.CLK(clknet_leaf_66_i_clk),
    .D(net663),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22482_ (.CLK(clknet_leaf_67_i_clk),
    .D(net1049),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03773_ (.A(_03773_),
    .X(clknet_0__03773_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03774_ (.A(_03774_),
    .X(clknet_0__03774_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03775_ (.A(_03775_),
    .X(clknet_0__03775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03776_ (.A(_03776_),
    .X(clknet_0__03776_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03777_ (.A(_03777_),
    .X(clknet_0__03777_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03778_ (.A(_03778_),
    .X(clknet_0__03778_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03779_ (.A(_03779_),
    .X(clknet_0__03779_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03780_ (.A(_03780_),
    .X(clknet_0__03780_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03781_ (.A(_03781_),
    .X(clknet_0__03781_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03980_ (.A(_03980_),
    .X(clknet_0__03980_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03981_ (.A(_03981_),
    .X(clknet_0__03981_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03982_ (.A(_03982_),
    .X(clknet_0__03982_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03983_ (.A(_03983_),
    .X(clknet_0__03983_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03984_ (.A(_03984_),
    .X(clknet_0__03984_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03985_ (.A(_03985_),
    .X(clknet_0__03985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03986_ (.A(_03986_),
    .X(clknet_0__03986_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03987_ (.A(_03987_),
    .X(clknet_0__03987_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03988_ (.A(_03988_),
    .X(clknet_0__03988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03989_ (.A(_03989_),
    .X(clknet_0__03989_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03990_ (.A(_03990_),
    .X(clknet_0__03990_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03991_ (.A(_03991_),
    .X(clknet_0__03991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03992_ (.A(_03992_),
    .X(clknet_0__03992_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03993_ (.A(_03993_),
    .X(clknet_0__03993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03994_ (.A(_03994_),
    .X(clknet_0__03994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03995_ (.A(_03995_),
    .X(clknet_0__03995_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03996_ (.A(_03996_),
    .X(clknet_0__03996_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03997_ (.A(_03997_),
    .X(clknet_0__03997_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03998_ (.A(_03998_),
    .X(clknet_0__03998_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03999_ (.A(_03999_),
    .X(clknet_0__03999_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04000_ (.A(_04000_),
    .X(clknet_0__04000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04001_ (.A(_04001_),
    .X(clknet_0__04001_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04002_ (.A(_04002_),
    .X(clknet_0__04002_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04003_ (.A(_04003_),
    .X(clknet_0__04003_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04004_ (.A(_04004_),
    .X(clknet_0__04004_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04005_ (.A(_04005_),
    .X(clknet_0__04005_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04006_ (.A(_04006_),
    .X(clknet_0__04006_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04007_ (.A(_04007_),
    .X(clknet_0__04007_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04008_ (.A(_04008_),
    .X(clknet_0__04008_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04009_ (.A(_04009_),
    .X(clknet_0__04009_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04010_ (.A(_04010_),
    .X(clknet_0__04010_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04011_ (.A(_04011_),
    .X(clknet_0__04011_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04012_ (.A(_04012_),
    .X(clknet_0__04012_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04800_ (.A(_04800_),
    .X(clknet_0__04800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05840_ (.A(_05840_),
    .X(clknet_0__05840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05891_ (.A(_05891_),
    .X(clknet_0__05891_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05942_ (.A(_05942_),
    .X(clknet_0__05942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05994_ (.A(_05994_),
    .X(clknet_0__05994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__06044_ (.A(_06044_),
    .X(clknet_0__06044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__06092_ (.A(_06092_),
    .X(clknet_0__06092_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03773_ (.A(clknet_0__03773_),
    .X(clknet_1_0__leaf__03773_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03774_ (.A(clknet_0__03774_),
    .X(clknet_1_0__leaf__03774_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03775_ (.A(clknet_0__03775_),
    .X(clknet_1_0__leaf__03775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03776_ (.A(clknet_0__03776_),
    .X(clknet_1_0__leaf__03776_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03777_ (.A(clknet_0__03777_),
    .X(clknet_1_0__leaf__03777_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03778_ (.A(clknet_0__03778_),
    .X(clknet_1_0__leaf__03778_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03779_ (.A(clknet_0__03779_),
    .X(clknet_1_0__leaf__03779_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03780_ (.A(clknet_0__03780_),
    .X(clknet_1_0__leaf__03780_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03781_ (.A(clknet_0__03781_),
    .X(clknet_1_0__leaf__03781_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03980_ (.A(clknet_0__03980_),
    .X(clknet_1_0__leaf__03980_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03981_ (.A(clknet_0__03981_),
    .X(clknet_1_0__leaf__03981_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03982_ (.A(clknet_0__03982_),
    .X(clknet_1_0__leaf__03982_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03983_ (.A(clknet_0__03983_),
    .X(clknet_1_0__leaf__03983_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03984_ (.A(clknet_0__03984_),
    .X(clknet_1_0__leaf__03984_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03985_ (.A(clknet_0__03985_),
    .X(clknet_1_0__leaf__03985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03986_ (.A(clknet_0__03986_),
    .X(clknet_1_0__leaf__03986_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03987_ (.A(clknet_0__03987_),
    .X(clknet_1_0__leaf__03987_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03988_ (.A(clknet_0__03988_),
    .X(clknet_1_0__leaf__03988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03989_ (.A(clknet_0__03989_),
    .X(clknet_1_0__leaf__03989_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03990_ (.A(clknet_0__03990_),
    .X(clknet_1_0__leaf__03990_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03991_ (.A(clknet_0__03991_),
    .X(clknet_1_0__leaf__03991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03992_ (.A(clknet_0__03992_),
    .X(clknet_1_0__leaf__03992_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03993_ (.A(clknet_0__03993_),
    .X(clknet_1_0__leaf__03993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03994_ (.A(clknet_0__03994_),
    .X(clknet_1_0__leaf__03994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03995_ (.A(clknet_0__03995_),
    .X(clknet_1_0__leaf__03995_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03996_ (.A(clknet_0__03996_),
    .X(clknet_1_0__leaf__03996_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03997_ (.A(clknet_0__03997_),
    .X(clknet_1_0__leaf__03997_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03998_ (.A(clknet_0__03998_),
    .X(clknet_1_0__leaf__03998_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03999_ (.A(clknet_0__03999_),
    .X(clknet_1_0__leaf__03999_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04000_ (.A(clknet_0__04000_),
    .X(clknet_1_0__leaf__04000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04001_ (.A(clknet_0__04001_),
    .X(clknet_1_0__leaf__04001_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04002_ (.A(clknet_0__04002_),
    .X(clknet_1_0__leaf__04002_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04003_ (.A(clknet_0__04003_),
    .X(clknet_1_0__leaf__04003_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04004_ (.A(clknet_0__04004_),
    .X(clknet_1_0__leaf__04004_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04005_ (.A(clknet_0__04005_),
    .X(clknet_1_0__leaf__04005_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04006_ (.A(clknet_0__04006_),
    .X(clknet_1_0__leaf__04006_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04007_ (.A(clknet_0__04007_),
    .X(clknet_1_0__leaf__04007_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04008_ (.A(clknet_0__04008_),
    .X(clknet_1_0__leaf__04008_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04009_ (.A(clknet_0__04009_),
    .X(clknet_1_0__leaf__04009_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04010_ (.A(clknet_0__04010_),
    .X(clknet_1_0__leaf__04010_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04011_ (.A(clknet_0__04011_),
    .X(clknet_1_0__leaf__04011_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04012_ (.A(clknet_0__04012_),
    .X(clknet_1_0__leaf__04012_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04800_ (.A(clknet_0__04800_),
    .X(clknet_1_0__leaf__04800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05840_ (.A(clknet_0__05840_),
    .X(clknet_1_0__leaf__05840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05891_ (.A(clknet_0__05891_),
    .X(clknet_1_0__leaf__05891_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05942_ (.A(clknet_0__05942_),
    .X(clknet_1_0__leaf__05942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05994_ (.A(clknet_0__05994_),
    .X(clknet_1_0__leaf__05994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__06044_ (.A(clknet_0__06044_),
    .X(clknet_1_0__leaf__06044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__06092_ (.A(clknet_0__06092_),
    .X(clknet_1_0__leaf__06092_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03773_ (.A(clknet_0__03773_),
    .X(clknet_1_1__leaf__03773_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03774_ (.A(clknet_0__03774_),
    .X(clknet_1_1__leaf__03774_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03775_ (.A(clknet_0__03775_),
    .X(clknet_1_1__leaf__03775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03776_ (.A(clknet_0__03776_),
    .X(clknet_1_1__leaf__03776_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03777_ (.A(clknet_0__03777_),
    .X(clknet_1_1__leaf__03777_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03778_ (.A(clknet_0__03778_),
    .X(clknet_1_1__leaf__03778_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03779_ (.A(clknet_0__03779_),
    .X(clknet_1_1__leaf__03779_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03780_ (.A(clknet_0__03780_),
    .X(clknet_1_1__leaf__03780_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03781_ (.A(clknet_0__03781_),
    .X(clknet_1_1__leaf__03781_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03980_ (.A(clknet_0__03980_),
    .X(clknet_1_1__leaf__03980_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03981_ (.A(clknet_0__03981_),
    .X(clknet_1_1__leaf__03981_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03982_ (.A(clknet_0__03982_),
    .X(clknet_1_1__leaf__03982_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03983_ (.A(clknet_0__03983_),
    .X(clknet_1_1__leaf__03983_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03984_ (.A(clknet_0__03984_),
    .X(clknet_1_1__leaf__03984_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03985_ (.A(clknet_0__03985_),
    .X(clknet_1_1__leaf__03985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03986_ (.A(clknet_0__03986_),
    .X(clknet_1_1__leaf__03986_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03987_ (.A(clknet_0__03987_),
    .X(clknet_1_1__leaf__03987_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03988_ (.A(clknet_0__03988_),
    .X(clknet_1_1__leaf__03988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03989_ (.A(clknet_0__03989_),
    .X(clknet_1_1__leaf__03989_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03990_ (.A(clknet_0__03990_),
    .X(clknet_1_1__leaf__03990_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03991_ (.A(clknet_0__03991_),
    .X(clknet_1_1__leaf__03991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03992_ (.A(clknet_0__03992_),
    .X(clknet_1_1__leaf__03992_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03993_ (.A(clknet_0__03993_),
    .X(clknet_1_1__leaf__03993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03994_ (.A(clknet_0__03994_),
    .X(clknet_1_1__leaf__03994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03995_ (.A(clknet_0__03995_),
    .X(clknet_1_1__leaf__03995_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03996_ (.A(clknet_0__03996_),
    .X(clknet_1_1__leaf__03996_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03997_ (.A(clknet_0__03997_),
    .X(clknet_1_1__leaf__03997_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03998_ (.A(clknet_0__03998_),
    .X(clknet_1_1__leaf__03998_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03999_ (.A(clknet_0__03999_),
    .X(clknet_1_1__leaf__03999_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04000_ (.A(clknet_0__04000_),
    .X(clknet_1_1__leaf__04000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04001_ (.A(clknet_0__04001_),
    .X(clknet_1_1__leaf__04001_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04002_ (.A(clknet_0__04002_),
    .X(clknet_1_1__leaf__04002_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04003_ (.A(clknet_0__04003_),
    .X(clknet_1_1__leaf__04003_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04004_ (.A(clknet_0__04004_),
    .X(clknet_1_1__leaf__04004_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04005_ (.A(clknet_0__04005_),
    .X(clknet_1_1__leaf__04005_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04006_ (.A(clknet_0__04006_),
    .X(clknet_1_1__leaf__04006_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04007_ (.A(clknet_0__04007_),
    .X(clknet_1_1__leaf__04007_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04008_ (.A(clknet_0__04008_),
    .X(clknet_1_1__leaf__04008_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04009_ (.A(clknet_0__04009_),
    .X(clknet_1_1__leaf__04009_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04010_ (.A(clknet_0__04010_),
    .X(clknet_1_1__leaf__04010_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04011_ (.A(clknet_0__04011_),
    .X(clknet_1_1__leaf__04011_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04012_ (.A(clknet_0__04012_),
    .X(clknet_1_1__leaf__04012_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04800_ (.A(clknet_0__04800_),
    .X(clknet_1_1__leaf__04800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05840_ (.A(clknet_0__05840_),
    .X(clknet_1_1__leaf__05840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05891_ (.A(clknet_0__05891_),
    .X(clknet_1_1__leaf__05891_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05942_ (.A(clknet_0__05942_),
    .X(clknet_1_1__leaf__05942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05994_ (.A(clknet_0__05994_),
    .X(clknet_1_1__leaf__05994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__06044_ (.A(clknet_0__06044_),
    .X(clknet_1_1__leaf__06044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__06092_ (.A(clknet_0__06092_),
    .X(clknet_1_1__leaf__06092_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_100_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_101_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_102_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net6321),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(net5709),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(net5711),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(net6542),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(net6544),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_01387_),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(net5720),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(net5722),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(net6228),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(net6230),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(net6231),
    .X(net1533));
 sky130_fd_sc_hd__buf_1 hold101 (.A(_03469_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(net6301),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(net6303),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_00808_),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(net7658),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_03420_),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(net4329),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(net6523),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(net6525),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_00812_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(net6548),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00954_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_03449_),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(_00940_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(net3099),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(_00916_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(net6042),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(net6044),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(net6045),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(net6577),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(net6579),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(_01497_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net6327),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(net5988),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(net5990),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_01447_),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(net5723),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(net5725),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(net6297),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_03430_),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(_00925_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\rbzero.spi_registers.buf_texadd2[14] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(net594),
    .X(net1563));
 sky130_fd_sc_hd__clkbuf_2 hold104 (.A(_02527_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_03414_),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(_00915_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(net6113),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(_03450_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_00941_),
    .X(net1568));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1045 (.A(net5779),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(net5781),
    .X(net1570));
 sky130_fd_sc_hd__buf_1 hold1047 (.A(net6270),
    .X(net1571));
 sky130_fd_sc_hd__buf_4 hold1048 (.A(_02986_),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(net5730),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00576_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(net6054),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(net6056),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_00922_),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(net6556),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_03979_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(_01266_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(net7627),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(net4724),
    .X(net1582));
 sky130_fd_sc_hd__buf_1 hold1059 (.A(net4468),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net823),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(net4470),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(net5713),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(net5715),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(net4614),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(net4616),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(net5735),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(net5737),
    .X(net1590));
 sky130_fd_sc_hd__buf_1 hold1067 (.A(net6057),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(net4225),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(net5742),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_03058_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(net5744),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(net6244),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(net6246),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(net6247),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(net4747),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(net4749),
    .X(net1599));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1076 (.A(net4264),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(net4864),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(net4866),
    .X(net1602));
 sky130_fd_sc_hd__buf_1 hold1079 (.A(net4274),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net4346),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(net6257),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(_03368_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_00882_),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(net3948),
    .X(net1607));
 sky130_fd_sc_hd__buf_4 hold1084 (.A(net3950),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(net5756),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(net6569),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(net6571),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_01333_),
    .X(net1612));
 sky130_fd_sc_hd__buf_1 hold1089 (.A(net6032),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net6315),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(net5764),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(net6558),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(net6560),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(_00810_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(net5749),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(net5751),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(net6597),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(net6599),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_01118_),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(net4728),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net6317),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(net4730),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(net6561),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_03378_),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(_00889_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(net6563),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(net6565),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_01567_),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(net6110),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_03453_),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(_00944_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_01362_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(net5782),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(_03082_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(net5997),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\rbzero.spi_registers.buf_texadd2[19] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(net1132),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(_03419_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_00920_),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(net6573),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(net6575),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(_01377_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net929),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(net6065),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(_03417_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_00918_),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(net6585),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_03377_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(_00888_),
    .X(net1649));
 sky130_fd_sc_hd__buf_1 hold1126 (.A(net5772),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(net5774),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(net6601),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(_03364_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_03059_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_00878_),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(net5794),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_03192_),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(net4228),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(net6617),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(net6619),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_01379_),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(net6232),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_03435_),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(_00930_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net5700),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(net6603),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(net6605),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_01486_),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(net6607),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_03366_),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(_00880_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(net6070),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(net6072),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(net6073),
    .X(net1672));
 sky130_fd_sc_hd__buf_1 hold1149 (.A(net4277),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net3285),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(net6663),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(_04432_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_01353_),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(net6703),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(net6705),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(_01499_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(net6581),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(net6583),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_01424_),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(net6879),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_03557_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(net5928),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(_01535_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(net6589),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(_03433_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_00928_),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(net7665),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_03438_),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(net6173),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(net6587),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(_03379_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net4676),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_00890_),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(net5757),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(net5759),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(net6849),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_04354_),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(_01423_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(net4671),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(net4673),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_00897_),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(net6299),
    .X(net1703));
 sky130_fd_sc_hd__buf_1 hold118 (.A(net6103),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_03363_),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(_00877_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(net6635),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(net6637),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_01409_),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(net6693),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_03432_),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(_00927_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(net6061),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(net6063),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_03021_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(net6064),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(net6655),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(net6657),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(_01339_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(net6649),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(_03447_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_00938_),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(net5787),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(net5789),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(net6651),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net4319),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(net6653),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(_01511_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(net6224),
    .X(net1726));
 sky130_fd_sc_hd__buf_4 hold1203 (.A(_03002_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(net5785),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(net6621),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_03385_),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(_00895_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(net6713),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(_04265_),
    .X(net1733));
 sky130_fd_sc_hd__buf_2 hold121 (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_01503_),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(net6289),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(net6291),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(net6292),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(net6613),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(net6615),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_01162_),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(net6767),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_04372_),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(_01407_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net4153),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(net6262),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(_03439_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_00934_),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(net6641),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(net6643),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(_01545_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(net7015),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(_04445_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_01341_),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(net6723),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net7659),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(net6725),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(_01154_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(net2172),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(_04485_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_01305_),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(net6743),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_04283_),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(_01487_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\rbzero.tex_r1[39] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(net5799),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_03444_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_01561_),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(net6677),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(net6679),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(_01371_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(net7667),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(_03386_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(net6105),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(net6645),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(net6647),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(_01411_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net5839),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(net6759),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(net6761),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_01554_),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(net6631),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(net6633),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(_01481_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(net5896),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(net5898),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_01427_),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\rbzero.spi_registers.buf_texadd2[16] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net4961),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(net1406),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(_03416_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_00917_),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(net6681),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_03398_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(_00903_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(net7674),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(_03250_),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(net6226),
    .X(net1792));
 sky130_fd_sc_hd__buf_1 hold1269 (.A(net7724),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net4963),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(net6791),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(net6793),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_01337_),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(net6683),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(net6685),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(_01385_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(net6695),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(_04509_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(_01283_),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(net6797),
    .X(net1803));
 sky130_fd_sc_hd__clkbuf_1 hold128 (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(net6799),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(_01113_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(net6255),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(_03406_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_00910_),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(net6775),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_04491_),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(_01299_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(net6961),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(net6963),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net4144),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_01369_),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(net6741),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(_04542_),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(_01160_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(net6827),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(net6829),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(_01495_),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(net6835),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_04359_),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_01419_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net4941),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(net6591),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(_04553_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_01150_),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(net5739),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(net5741),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(net6629),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(_03367_),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(_00881_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(net5847),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(net5849),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net4943),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(_01327_),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(net6901),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_04174_),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(_01583_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(net6707),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(net6709),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_01285_),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(net6673),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(net6675),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(_01479_),
    .X(net1843));
 sky130_fd_sc_hd__buf_1 hold132 (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(net6059),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(_03451_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(_00942_),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(net6721),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_03452_),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(_00943_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(net6669),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(net6671),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_01347_),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(net6687),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net4174),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(net6689),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(_01565_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(net6735),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(net5869),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_01308_),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(net7664),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_03383_),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(net6030),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\rbzero.spi_registers.buf_texadd3[20] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(_03455_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net4950),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(net4323),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(net6981),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(_04358_),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(_01420_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(net6739),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_03399_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_00904_),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(net6719),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_03434_),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(_00929_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net4952),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(net5889),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(net5891),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(_01269_),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(net6609),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(net6611),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_01367_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(net6757),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(_04508_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_01284_),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(net6235),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net4955),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_03402_),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(_00906_),
    .X(net1885));
 sky130_fd_sc_hd__clkbuf_2 hold1362 (.A(net7655),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(net4939),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(net6639),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(_04443_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_01343_),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(net6625),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(net6627),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(_01557_),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net4957),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(net6821),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(_04564_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_01140_),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(net6801),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_04398_),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(_01383_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(net6867),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(net6869),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_01531_),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(net6623),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net4958),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(_03431_),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_00926_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(net6691),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(_04531_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_01170_),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(net6567),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_03397_),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_00902_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(net6284),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(_03373_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net4960),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_00886_),
    .X(net1914));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1391 (.A(net5801),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(net5803),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(net6715),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(net6717),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(_01350_),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(net6554),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(_04155_),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_01645_),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(net7224),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net4964),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(net6737),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(_01307_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(net7070),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(_04452_),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_01335_),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(net2033),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_04528_),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(_01172_),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(net7017),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(net5805),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net4966),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_01520_),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(net6965),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(net6967),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(_01346_),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(net5984),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(net5986),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_01365_),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(net5930),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(net5932),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(_01441_),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net4944),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(net6665),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(net6667),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_01356_),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(net6731),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(net6733),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(_01123_),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(net6931),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_04400_),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(_01381_),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(net7003),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net4946),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_04248_),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(_01519_),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(net2023),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(net5835),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(_01364_),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(net7663),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(net4245),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(net6975),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(_04546_),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(_01156_),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\rbzero.pov.ready_buffer[55] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(net6659),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(_03436_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(_00931_),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(net2288),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(net5818),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(_01167_),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(net5952),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(net5954),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_01168_),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(net6701),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_03563_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(_04298_),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(_01473_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net7078),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(net7080),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_01510_),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(net6777),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_04382_),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(_01398_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(net2770),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(_04387_),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net4388),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(_01393_),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(net6891),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(_04442_),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(_01344_),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(\rbzero.spi_registers.buf_texadd3[12] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(net600),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(_03446_),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(_00937_),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(net5810),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(net5812),
    .X(net1993));
 sky130_fd_sc_hd__buf_1 hold147 (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(_01560_),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(net6877),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_04401_),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(_01380_),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_06626_),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(net7631),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(net4755),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(net2233),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(net5855),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(_01426_),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net4161),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(net6985),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(_04371_),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(_01408_),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(net6851),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(_04218_),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(_01543_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(net7057),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(_04297_),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(_01474_),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\rbzero.spi_registers.buf_texadd3[11] ),
    .X(net2013));
 sky130_fd_sc_hd__buf_1 hold149 (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(net597),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(_03445_),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(_00936_),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(net6751),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(net6753),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(_01436_),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(net6783),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(_03418_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(_00919_),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\rbzero.tex_g0[33] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net4168),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(net1956),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(_04421_),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(_01363_),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(net6871),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(net6873),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(_01142_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(net6947),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(net6949),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_01132_),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\rbzero.tex_b0[63] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\rbzero.pov.ready_buffer[70] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(net1929),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(_04527_),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(_01173_),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\rbzero.tex_b1[1] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(net5842),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(_01268_),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(net7068),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(_04296_),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(_01475_),
    .X(net2042));
 sky130_fd_sc_hd__clkbuf_2 hold1519 (.A(net5807),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_03514_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(net5809),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(net7033),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(_04347_),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(_01430_),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(net6769),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(_04425_),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(_01359_),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(net6955),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(_04558_),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(_01145_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net6183),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(net6711),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(_04287_),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_01483_),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(net6987),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(net6989),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(_01455_),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(net6795),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(_04282_),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_01488_),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(net6697),
    .X(net2063));
 sky130_fd_sc_hd__buf_1 hold154 (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(net6699),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(_01471_),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(net6817),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(net6819),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_01571_),
    .X(net2068));
 sky130_fd_sc_hd__clkbuf_2 hold1545 (.A(net4390),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(net7661),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(_03437_),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(net6165),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(net6745),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net4177),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(net6747),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(_01146_),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(net6853),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(_03365_),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_00879_),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(net6897),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(net6899),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(_01529_),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(net6847),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(_04196_),
    .X(net2083));
 sky130_fd_sc_hd__buf_1 hold156 (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_01563_),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\rbzero.tex_r1[14] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(net6881),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(_01536_),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(net3111),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(_00907_),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(net6169),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(_03370_),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_00884_),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\rbzero.spi_registers.buf_texadd2[13] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net4137),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(net591),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(_03412_),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_00914_),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(net5878),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(net5880),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(_01397_),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(\rbzero.tex_r0[59] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(net1472),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_04249_),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(_01518_),
    .X(net2103));
 sky130_fd_sc_hd__buf_1 hold158 (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(net6779),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(_04523_),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_01270_),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(net6823),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(net6825),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_01467_),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(net6915),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(net6917),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_01456_),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(net6661),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net4134),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(_03401_),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(_00905_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(net6979),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(_04446_),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(_01340_),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(net2196),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(net5866),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(_01294_),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(net4883),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(_03029_),
    .X(net2123));
 sky130_fd_sc_hd__buf_1 hold160 (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_00654_),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(net6889),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_04349_),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(_01428_),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(net7082),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(_04430_),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_01355_),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(net7011),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(_04390_),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(_01390_),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net4187),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(net6875),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(_04369_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_01410_),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(net6909),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_04185_),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(_01573_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(net6883),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(net5815),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(_01326_),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(net6991),
    .X(net2143));
 sky130_fd_sc_hd__clkbuf_1 hold162 (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_04303_),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(_01469_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(net6845),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(_04538_),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_01163_),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(net6763),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(net6765),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(_01320_),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(net2517),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_04200_),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net4180),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(_01559_),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(net5860),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_03448_),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(_00939_),
    .X(net2157));
 sky130_fd_sc_hd__buf_1 hold1634 (.A(net4678),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(net4680),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(net7037),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(net7039),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_01165_),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(net6921),
    .X(net2163));
 sky130_fd_sc_hd__buf_1 hold164 (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_04312_),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(_01461_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(net6925),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(_04506_),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_01286_),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(net7202),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(_04263_),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(_01505_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(\rbzero.tex_b1[39] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(net1756),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net4156),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(_04484_),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(_01306_),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(net5903),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(net5905),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(_01309_),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(net2411),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(net5901),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(_01290_),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(net5961),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(net5963),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(net4967),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(_01291_),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(net7053),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(_04495_),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(_01296_),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(net6749),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(_04479_),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_01310_),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(net5934),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(net5936),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(_01331_),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net4969),
    .X(net691));
 sky130_fd_sc_hd__buf_1 hold1670 (.A(net5851),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(net5853),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\rbzero.tex_b1[27] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(net2119),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_04498_),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(_01293_),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(net6841),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(_04476_),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(_01313_),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(net7047),
    .X(net2203));
 sky130_fd_sc_hd__buf_1 hold168 (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_04575_),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(_01130_),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(net6789),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(_04490_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(_01300_),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(net6929),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(_04339_),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(_01437_),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(net7118),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(net6885),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net4147),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(_01325_),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(net7009),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(_04589_),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(_01117_),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(net6939),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(_04410_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(_01373_),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(net7072),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_04232_),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(_01530_),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net4108),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(net6781),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(_04193_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(_01566_),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(net6911),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(_04489_),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(_01301_),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(net6036),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(net6038),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(net6039),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\rbzero.tex_g1[31] ),
    .X(net2233));
 sky130_fd_sc_hd__clkbuf_2 hold171 (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(net2001),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(_04352_),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(_01425_),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(net7027),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(_04418_),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(_01366_),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(net6855),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(net6857),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_01414_),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(net2448),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(net4131),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(_04458_),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(_01329_),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(net7074),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(net7076),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(_01444_),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(net7045),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(_04472_),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(_01317_),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\rbzero.tex_g1[48] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(net932),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net3087),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(_04331_),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(_01443_),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(net6179),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(_03372_),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(_00885_),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(net2698),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(_04228_),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(_01534_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(net7025),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(_04173_),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_03345_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(_01584_),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(net7094),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(_04409_),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(_01374_),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(net6951),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(net6953),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(_01126_),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(net7049),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(_04441_),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(_01345_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net4116),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(net6729),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(_03369_),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(_00883_),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(net6803),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(_04568_),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(_01136_),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(net4267),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(net4269),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(net6050),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(net6052),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(net7483),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(net6053),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(net6971),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(net6973),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(_01315_),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\rbzero.tex_b0[57] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(net1967),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(_04535_),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(_01166_),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(net7114),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(net7116),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net7613),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(_01466_),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(net6831),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(net6833),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(_01138_),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(net7043),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(_04195_),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(_01564_),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(net6997),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(net6999),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(_01389_),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(net4426),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(net6771),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(net6773),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(_01501_),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(net7172),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(_04273_),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(_01496_),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(net7100),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(net7102),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(_01434_),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(net6923),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(net5029),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_04423_),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(_01361_),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(net7178),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(_04549_),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(_01153_),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(net6859),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(_04518_),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(_01275_),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(net7041),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(_04473_),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net5031),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(_01316_),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(net7144),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(_04381_),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(_01399_),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(net6785),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(net6787),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(_01544_),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(net6837),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(net6839),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(_01143_),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net3421),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(net6903),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(_04326_),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(_01448_),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(net2366),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(_04246_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(_01521_),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(net6861),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(net6863),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(_01279_),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(net7055),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net4365),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(_04205_),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(_01555_),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(net7134),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(_04544_),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(_01158_),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(net6755),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(_04453_),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(_01334_),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(net7673),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(net5863),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(net4974),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(net6075),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(net6077),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(_00923_),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(net7051),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(_04365_),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(_01413_),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(net6843),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(_04431_),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(_01354_),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(net7152),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(net4976),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(net7154),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(_01575_),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(\rbzero.tex_r0[63] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(net2337),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(_04245_),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(_01522_),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(net6919),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(_04594_),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(_01112_),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(net6941),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net4545),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(_04215_),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(_01546_),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(net6865),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(_04293_),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(_01478_),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(net7005),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(_04190_),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(_01568_),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(\rbzero.tex_r1[6] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(net7090),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net4547),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(_01528_),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(net7065),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(net7067),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(_01463_),
    .X(net2387));
 sky130_fd_sc_hd__clkbuf_2 hold1864 (.A(net7650),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(net4825),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(net6727),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(_04552_),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(_01151_),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(net5885),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(net4394),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(net5887),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(_01526_),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(net2707),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(net5845),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(_01440_),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(net7029),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(_04555_),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(_01148_),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(net6913),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(_04424_),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(net4396),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(_01360_),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\rbzero.tex_r1[47] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(net7007),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(_01569_),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(net6983),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(_04590_),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(_01116_),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\rbzero.tex_b1[23] ),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(net2179),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(_04502_),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net3295),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(_01289_),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(net7086),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(_04530_),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(_01171_),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(net7242),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(_04254_),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(_01513_),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(net6935),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(_04269_),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(_01500_),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(net4516),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(net7112),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(_04413_),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(_01370_),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\rbzero.tex_r1[59] ),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(net5825),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(_01581_),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(net6933),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(_04567_),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(_01137_),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(net6813),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(net7614),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(net6815),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(_01318_),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(net7019),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(_04522_),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(_01271_),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(net7063),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(_04393_),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(_01388_),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(\rbzero.tex_g1[1] ),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(net5832),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net4659),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(_01396_),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(net6943),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(net6945),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(_01491_),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(\rbzero.tex_b1[63] ),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(net2243),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(_04457_),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(_01330_),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(net7156),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(_04325_),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net4986),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(_01449_),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(net6194),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(_03404_),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(_00908_),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(net7084),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(_04302_),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(_01470_),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(net7126),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(_04338_),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(_01438_),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net4988),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(net5871),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(net5873),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(_01295_),
    .X(net2466));
 sky130_fd_sc_hd__buf_1 hold1943 (.A(net5882),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(net5884),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(net6905),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(net6907),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(_01570_),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(net5827),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(net5829),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net7632),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(_01580_),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(net7035),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(_04291_),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(_01480_),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(net7104),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(_04376_),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(_01403_),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(net6805),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(net6807),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(_01133_),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net4642),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(net7208),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(_04213_),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(_01547_),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(net7194),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(_03381_),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(_00892_),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(net7182),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(_04357_),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(_01421_),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(net5980),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(net7621),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(net5982),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(_01551_),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(\rbzero.tex_g1[56] ),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(net7158),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(_01450_),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(net7232),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(_04262_),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(_01506_),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(net7122),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(_04545_),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net4522),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(_01157_),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(net7059),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(net7061),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(_01515_),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(net7200),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(_04494_),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(_01297_),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(net6969),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(_04578_),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(_01127_),
    .X(net2513));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold199 (.A(net7615),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(net6957),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(net6959),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(_01401_),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\rbzero.tex_r1[36] ),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(net2152),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(_04201_),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(_01558_),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(net7110),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(_04449_),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(_01338_),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(net4440),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(net6893),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(net6895),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(_01416_),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(net7031),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(_04428_),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(_01357_),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(net7013),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(_04550_),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(_01152_),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(net6201),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net3523),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(_03405_),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(_00909_),
    .X(net2535));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2012 (.A(net5875),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(net5877),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(net7142),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(_04408_),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(_01375_),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(net7672),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(_03267_),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(net6272),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_03518_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(net7214),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(_04475_),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(_01314_),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(net7021),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(net7023),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(_01404_),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(net6993),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(net6995),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(_01376_),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(net6274),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net6211),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(net6276),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(net6277),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(net7240),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(net5915),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(_01550_),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(net7220),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(_04295_),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(_01476_),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(net5910),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(net5912),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net6332),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(_01460_),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(net2577),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(_04464_),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(_01324_),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(net7140),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(_04204_),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(_01556_),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(net7160),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(_04182_),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(_01576_),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net6334),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(net2819),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(_04178_),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2052 (.A(_01579_),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(\rbzero.tex_b1[57] ),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(net2565),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(_04465_),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(_01323_),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(net6887),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(_04556_),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(_01147_),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_01119_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2060 (.A(net6937),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(_04512_),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2062 (.A(_01280_),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(net7106),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(_04487_),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(_01303_),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2066 (.A(net6293),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(net6295),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(net6296),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(net6927),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net3316),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(_03380_),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2071 (.A(_00891_),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(net7096),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(_04486_),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(_01304_),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(net7128),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2076 (.A(net7130),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2077 (.A(_01400_),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(net7180),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(_04184_),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net4636),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(_01574_),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2081 (.A(net6809),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(net6811),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(_01274_),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(net6977),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(_04581_),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(_01124_),
    .X(net2610));
 sky130_fd_sc_hd__buf_1 hold2087 (.A(net5968),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2088 (.A(net5970),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(net7293),
    .X(net2613));
 sky130_fd_sc_hd__buf_1 hold209 (.A(\rbzero.pov.ready_buffer[59] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(_04537_),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(_01164_),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(net7092),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(_04451_),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(_01336_),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(net7222),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(_04563_),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2097 (.A(_01141_),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(net7190),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(_04264_),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_03482_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(_01504_),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2101 (.A(net7166),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(_04320_),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(_01453_),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(\rbzero.pov.spi_counter[1] ),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2105 (.A(_03657_),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(_03662_),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(net4798),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2108 (.A(net7228),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(net5894),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net4336),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(_01446_),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(net7174),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2112 (.A(_04207_),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(_01553_),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(net7108),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(_04363_),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2116 (.A(_01415_),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2117 (.A(net7148),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(net7150),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(_01490_),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net4990),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(net7162),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(net7164),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2122 (.A(_01494_),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2123 (.A(net2685),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(_04172_),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(_01585_),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(net5923),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2127 (.A(net5925),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2128 (.A(_01111_),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(net7001),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net4992),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(_04520_),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(_01273_),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(net7210),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2133 (.A(_04577_),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(_01128_),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(net7098),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(_04395_),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(_01386_),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(net7244),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2139 (.A(_04405_),
    .X(net2663));
 sky130_fd_sc_hd__buf_1 hold214 (.A(net7616),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(_01378_),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(net7216),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(_04438_),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(_01348_),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(net7283),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2145 (.A(_04281_),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(_01489_),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(net7259),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(_04389_),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(_01391_),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net4623),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(net7226),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2151 (.A(_04343_),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(_01433_),
    .X(net2676));
 sky130_fd_sc_hd__clkbuf_2 hold2153 (.A(net5907),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(net5909),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(net7120),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(_04251_),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2157 (.A(_01516_),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2158 (.A(net7246),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(_04308_),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net3427),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(_01464_),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(\rbzero.tex_r1[63] ),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2162 (.A(net2647),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(_04171_),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(_01586_),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(net7192),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(_04260_),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(_01508_),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(net7218),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2169 (.A(_04586_),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(net4461),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(_01120_),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(net7234),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2172 (.A(net7236),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2173 (.A(_01465_),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(\rbzero.tex_r1[11] ),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(net2259),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(_04229_),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(_01533_),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(net7265),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2179 (.A(_04222_),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net5010),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(_01539_),
    .X(net2704));
 sky130_fd_sc_hd__clkbuf_2 hold2181 (.A(net5943),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(net5945),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(\rbzero.tex_g1[45] ),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2184 (.A(net2396),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(_04337_),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(_01439_),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(net7124),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(_04574_),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2189 (.A(_01131_),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(net5012),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(net7299),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2191 (.A(_04311_),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(_01462_),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(net7254),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(_04436_),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(_01349_),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(net2746),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2197 (.A(_04316_),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(_01457_),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2199 (.A(net7248),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\rbzero.pov.ready_buffer[68] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(_04238_),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(_01525_),
    .X(net2725));
 sky130_fd_sc_hd__clkbuf_2 hold2202 (.A(net5938),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(net5940),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(net7168),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(net7170),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(_01537_),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(net7196),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(net7198),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(_01540_),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_03506_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(net7136),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(net7138),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(_01122_),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(net7212),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(_04346_),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2215 (.A(_01431_),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(net7273),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(_04434_),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(_01351_),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(net7238),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net6156),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(_04469_),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(_01319_),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(\rbzero.tex_g1[63] ),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(net2720),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(_04315_),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(_01458_),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(net7271),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2227 (.A(_04180_),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(_01577_),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(net7277),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\rbzero.pov.ready_buffer[56] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(_04239_),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(_01524_),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2232 (.A(net7281),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(_04253_),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(_01514_),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(net7206),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(_04271_),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2237 (.A(_01498_),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(\rbzero.tex_g1[50] ),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(net7230),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_03567_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(_01445_),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(net7132),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2242 (.A(_04361_),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2243 (.A(_01417_),
    .X(net2767));
 sky130_fd_sc_hd__buf_1 hold2244 (.A(net5705),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2245 (.A(net5707),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(\rbzero.tex_g0[63] ),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(net1982),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(_04386_),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2249 (.A(_01394_),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net6214),
    .X(net749));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2250 (.A(net5965),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(net5967),
    .X(net2775));
 sky130_fd_sc_hd__buf_1 hold2252 (.A(net4648),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(net4650),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2254 (.A(net2854),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(_04211_),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(_01549_),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(net7176),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(_04319_),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2259 (.A(_01454_),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\rbzero.tex_g0[2] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(net7186),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(net7188),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2262 (.A(_01277_),
    .X(net2786));
 sky130_fd_sc_hd__buf_1 hold2263 (.A(net5745),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(net5747),
    .X(net2788));
 sky130_fd_sc_hd__clkbuf_2 hold2265 (.A(net5977),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(net5979),
    .X(net2790));
 sky130_fd_sc_hd__clkbuf_2 hold2267 (.A(net5946),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(net5948),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(net7263),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net5921),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(_04592_),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2271 (.A(_01114_),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(net7250),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(_04505_),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2274 (.A(_01287_),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(net7269),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2276 (.A(_04541_),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(_01161_),
    .X(net2801));
 sky130_fd_sc_hd__clkbuf_2 hold2278 (.A(net5917),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2279 (.A(net5919),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_01332_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(net7257),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2281 (.A(_04570_),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(_01134_),
    .X(net2806));
 sky130_fd_sc_hd__clkbuf_2 hold2283 (.A(net7653),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2284 (.A(net4878),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2285 (.A(net7275),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(_04585_),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(_01121_),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(net7310),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2289 (.A(_03508_),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net4994),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(_03510_),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(_00965_),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(net7184),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(_04580_),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(_01125_),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(\rbzero.tex_r1[56] ),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(net2574),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(_04179_),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(_01578_),
    .X(net2822));
 sky130_fd_sc_hd__clkbuf_2 hold2299 (.A(net5992),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(net4996),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2300 (.A(net5994),
    .X(net2824));
 sky130_fd_sc_hd__clkbuf_2 hold2301 (.A(net5949),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(net5951),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(net7279),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(_04220_),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(_01541_),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2306 (.A(net7287),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2307 (.A(_04341_),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(_01435_),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(net4775),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net5013),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2310 (.A(net4777),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(net3572),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2312 (.A(_03535_),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2313 (.A(_03536_),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(net6083),
    .X(net2838));
 sky130_fd_sc_hd__clkbuf_2 hold2315 (.A(net5972),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(net5974),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(net3944),
    .X(net2841));
 sky130_fd_sc_hd__buf_2 hold2318 (.A(net3946),
    .X(net2842));
 sky130_fd_sc_hd__clkbuf_4 hold2319 (.A(_03008_),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net5015),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(_00644_),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2321 (.A(net7289),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2322 (.A(_04276_),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(_01493_),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2324 (.A(net7291),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(_04259_),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2326 (.A(_01509_),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(net7261),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(_04286_),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(_01484_),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(net7492),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(\rbzero.tex_r1[26] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2331 (.A(net2778),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(_04212_),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2333 (.A(_01548_),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(net7267),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(_04517_),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2336 (.A(_01276_),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(net7303),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2338 (.A(net7305),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(_01451_),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net5060),
    .X(net758));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2340 (.A(net5958),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(net5960),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2342 (.A(net7252),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2343 (.A(_04511_),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2344 (.A(_01281_),
    .X(net2868));
 sky130_fd_sc_hd__buf_2 hold2345 (.A(net7888),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2346 (.A(net7301),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2347 (.A(_04416_),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(_01368_),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(net7666),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net5062),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(_03458_),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2351 (.A(net6034),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2352 (.A(net7285),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(_04374_),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2354 (.A(_01405_),
    .X(net2878));
 sky130_fd_sc_hd__clkbuf_2 hold2355 (.A(net6001),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(net6003),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(net7297),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(_04515_),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(_01278_),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net6336),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2360 (.A(net6221),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(net6223),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2362 (.A(_00600_),
    .X(net2886));
 sky130_fd_sc_hd__buf_1 hold2363 (.A(net7678),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2364 (.A(net4602),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(net3579),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(_03545_),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(net6128),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(net3359),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2369 (.A(_03556_),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(net6338),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2370 (.A(_00979_),
    .X(net2894));
 sky130_fd_sc_hd__buf_1 hold2371 (.A(net5998),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2372 (.A(net6000),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(net7295),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2374 (.A(_04397_),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2375 (.A(_01384_),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2376 (.A(net6019),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(net6021),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2378 (.A(net7308),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2379 (.A(_04285_),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_01272_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(_01485_),
    .X(net2904));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2381 (.A(net6004),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2382 (.A(net6006),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2383 (.A(net5490),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(net5492),
    .X(net2908));
 sky130_fd_sc_hd__buf_1 hold2385 (.A(net4743),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(net4745),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2387 (.A(net3364),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2388 (.A(_03534_),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(net4356),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net5006),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2390 (.A(\rbzero.pov.ready_buffer[51] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2391 (.A(_03549_),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(net4359),
    .X(net2916));
 sky130_fd_sc_hd__buf_1 hold2393 (.A(net6013),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2394 (.A(net6015),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2396 (.A(net6242),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(_00578_),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(net3610),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(_03541_),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(net5008),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2400 (.A(_00973_),
    .X(net2924));
 sky130_fd_sc_hd__buf_1 hold2401 (.A(net6016),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2402 (.A(net6018),
    .X(net2926));
 sky130_fd_sc_hd__buf_1 hold2403 (.A(\rbzero.pov.ready_buffer[65] ),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(_03497_),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(_03498_),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2406 (.A(net6131),
    .X(net2930));
 sky130_fd_sc_hd__buf_1 hold2407 (.A(net4739),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(net4741),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(net5462),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net5025),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(net5464),
    .X(net2934));
 sky130_fd_sc_hd__buf_2 hold2411 (.A(net7904),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2412 (.A(net6011),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(net7329),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(_03660_),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(net6177),
    .X(net2939));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2416 (.A(net4892),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2417 (.A(net4894),
    .X(net2941));
 sky130_fd_sc_hd__clkbuf_2 hold2418 (.A(net6096),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(net7733),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net5027),
    .X(net766));
 sky130_fd_sc_hd__buf_1 hold2420 (.A(\rbzero.pov.ready_buffer[64] ),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(_03494_),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(_03495_),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(net4301),
    .X(net2947));
 sky130_fd_sc_hd__buf_1 hold2424 (.A(net6046),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2425 (.A(_03025_),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2426 (.A(_00651_),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(\rbzero.spi_registers.buf_floor[3] ),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2428 (.A(net7328),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(_03101_),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net4606),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2430 (.A(_00697_),
    .X(net2954));
 sky130_fd_sc_hd__buf_2 hold2431 (.A(net4610),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2432 (.A(\rbzero.pov.ready_buffer[50] ),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(_03547_),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(net6192),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(net7736),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(_08244_),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(net4830),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(net4400),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2439 (.A(_00649_),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net4608),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(\rbzero.spi_registers.buf_sky[2] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2441 (.A(net7323),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2442 (.A(_03090_),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(_00690_),
    .X(net2967));
 sky130_fd_sc_hd__buf_1 hold2444 (.A(net4704),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(net4706),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(net3108),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(_03020_),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(_00647_),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(\rbzero.spi_registers.buf_floor[1] ),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net5071),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2450 (.A(net7326),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2451 (.A(_03098_),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(_00695_),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(\rbzero.spi_registers.sclk_buffer[2] ),
    .X(net2977));
 sky130_fd_sc_hd__buf_2 hold2454 (.A(_02524_),
    .X(net2978));
 sky130_fd_sc_hd__clkbuf_2 hold2455 (.A(_02989_),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(_03024_),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(_00650_),
    .X(net2981));
 sky130_fd_sc_hd__clkbuf_2 hold2458 (.A(net6167),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(_04131_),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(net5073),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(net6252),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(net7726),
    .X(net2985));
 sky130_fd_sc_hd__buf_2 hold2462 (.A(net4890),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2463 (.A(_04854_),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2464 (.A(_03951_),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(net6026),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(\rbzero.pov.ready_buffer[48] ),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(_03543_),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2468 (.A(net4295),
    .X(net2992));
 sky130_fd_sc_hd__clkbuf_2 hold2469 (.A(net6022),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net5002),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(_00487_),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2471 (.A(net7366),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2472 (.A(_03092_),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2473 (.A(_03093_),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(_00692_),
    .X(net2998));
 sky130_fd_sc_hd__buf_1 hold2475 (.A(\rbzero.pov.ready_buffer[66] ),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2476 (.A(_03499_),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(_03500_),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(net6200),
    .X(net3002));
 sky130_fd_sc_hd__clkbuf_2 hold2479 (.A(net6126),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net5004),
    .X(net772));
 sky130_fd_sc_hd__buf_1 hold2480 (.A(_09522_),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(net4309),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(net4788),
    .X(net3007));
 sky130_fd_sc_hd__clkbuf_2 hold2484 (.A(net6129),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2485 (.A(_09643_),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(\rbzero.spi_registers.buf_texadd1[10] ),
    .X(net3010));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2487 (.A(net618),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(_03376_),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(_00887_),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net7676),
    .X(net773));
 sky130_fd_sc_hd__buf_4 hold2490 (.A(net4531),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(net4533),
    .X(net3015));
 sky130_fd_sc_hd__clkbuf_2 hold2492 (.A(net4316),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(net7792),
    .X(net3017));
 sky130_fd_sc_hd__buf_1 hold2494 (.A(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(net6320),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(_00614_),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2497 (.A(net6234),
    .X(net3021));
 sky130_fd_sc_hd__buf_2 hold2498 (.A(net612),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2499 (.A(_00639_),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net7517),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 hold2500 (.A(net6081),
    .X(net3024));
 sky130_fd_sc_hd__buf_1 hold2501 (.A(_09285_),
    .X(net3025));
 sky130_fd_sc_hd__clkbuf_4 hold2502 (.A(net4682),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(net4684),
    .X(net3027));
 sky130_fd_sc_hd__clkbuf_4 hold2504 (.A(net6198),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2505 (.A(net7447),
    .X(net3029));
 sky130_fd_sc_hd__buf_1 hold2506 (.A(\rbzero.pov.ready_buffer[62] ),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(_03490_),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2508 (.A(_03491_),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2509 (.A(net4339),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net4978),
    .X(net775));
 sky130_fd_sc_hd__buf_1 hold2510 (.A(net6308),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(net6310),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(_00598_),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .X(net3037));
 sky130_fd_sc_hd__clkbuf_4 hold2514 (.A(net616),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2515 (.A(_00640_),
    .X(net3039));
 sky130_fd_sc_hd__clkbuf_2 hold2516 (.A(net4343),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2517 (.A(net7823),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(net7907),
    .X(net3042));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2519 (.A(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net4980),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(_02701_),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2521 (.A(net4813),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(net7480),
    .X(net3046));
 sky130_fd_sc_hd__buf_1 hold2523 (.A(net7547),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(_08220_),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2525 (.A(net6283),
    .X(net3049));
 sky130_fd_sc_hd__clkbuf_2 hold2526 (.A(net6163),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(_00635_),
    .X(net3051));
 sky130_fd_sc_hd__buf_1 hold2528 (.A(net6197),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2529 (.A(_00637_),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net5052),
    .X(net777));
 sky130_fd_sc_hd__buf_1 hold2530 (.A(net4535),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(_08225_),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(net4785),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(net4352),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2534 (.A(net3741),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2535 (.A(_02475_),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(_02482_),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2537 (.A(_02483_),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2538 (.A(_02484_),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(net5683),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net5054),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2540 (.A(net5685),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2541 (.A(net7828),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2542 (.A(net4928),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(_08216_),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2544 (.A(net6280),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .X(net3069));
 sky130_fd_sc_hd__buf_2 hold2546 (.A(net910),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(_00642_),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2548 (.A(net6028),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(_00645_),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net4982),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_2 hold2550 (.A(net7311),
    .X(net3074));
 sky130_fd_sc_hd__buf_2 hold2551 (.A(_02493_),
    .X(net3075));
 sky130_fd_sc_hd__clkbuf_2 hold2552 (.A(_03251_),
    .X(net3076));
 sky130_fd_sc_hd__buf_2 hold2553 (.A(_03252_),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(_03254_),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2555 (.A(_03255_),
    .X(net3079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(_00809_),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2557 (.A(\rbzero.pov.ready_buffer[57] ),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(_03570_),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2559 (.A(_03572_),
    .X(net3083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net4984),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2560 (.A(_00983_),
    .X(net3084));
 sky130_fd_sc_hd__clkbuf_2 hold2561 (.A(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(net3085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2562 (.A(net4872),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .X(net3087));
 sky130_fd_sc_hd__clkbuf_4 hold2564 (.A(net697),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2565 (.A(_00641_),
    .X(net3089));
 sky130_fd_sc_hd__clkbuf_2 hold2566 (.A(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2567 (.A(_02918_),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2568 (.A(net4819),
    .X(net3092));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2569 (.A(net6171),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net5033),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2570 (.A(_00636_),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2571 (.A(net6196),
    .X(net3095));
 sky130_fd_sc_hd__buf_4 hold2572 (.A(net3052),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2573 (.A(_03010_),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(_00638_),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .X(net3099));
 sky130_fd_sc_hd__clkbuf_4 hold2576 (.A(net1546),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2577 (.A(_00643_),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2578 (.A(net7795),
    .X(net3102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(net7916),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net5035),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(net3939),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(_03248_),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2582 (.A(_03249_),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(_00806_),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(net6145),
    .X(net3108));
 sky130_fd_sc_hd__clkbuf_2 hold2585 (.A(net2970),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2586 (.A(_00646_),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .X(net3111));
 sky130_fd_sc_hd__clkbuf_4 hold2588 (.A(net2088),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(_00634_),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net5037),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2590 (.A(net7489),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2591 (.A(net7817),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(\rbzero.spi_registers.buf_floor[5] ),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2593 (.A(_03262_),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(_03263_),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(_00813_),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(net7813),
    .X(net3120));
 sky130_fd_sc_hd__clkbuf_1 hold2597 (.A(_04618_),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2598 (.A(net4733),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(net3932),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net5039),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2600 (.A(_03257_),
    .X(net3124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2601 (.A(_03258_),
    .X(net3125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2602 (.A(_00811_),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(net4379),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(\rbzero.color_floor[5] ),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2605 (.A(_03103_),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(_03104_),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2607 (.A(_00699_),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(\rbzero.side_hot ),
    .X(net3480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2609 (.A(_02806_),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net7472),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2610 (.A(net4628),
    .X(net3134));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2611 (.A(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(net7321),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(_00612_),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2614 (.A(net7781),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(\rbzero.pov.ready_buffer[39] ),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(net7351),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2617 (.A(_03592_),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(_00991_),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(net7788),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net5044),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(\rbzero.color_sky[0] ),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2621 (.A(_03085_),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(_03086_),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2623 (.A(_00688_),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2624 (.A(net4392),
    .X(net3148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(net7595),
    .X(net3149));
 sky130_fd_sc_hd__clkbuf_2 hold2626 (.A(net7338),
    .X(net3150));
 sky130_fd_sc_hd__buf_2 hold2627 (.A(_02494_),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2628 (.A(_03460_),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(_03461_),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(net5046),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(_00949_),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(net4402),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2632 (.A(\rbzero.pov.ready_buffer[73] ),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(_03526_),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2634 (.A(_03527_),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(_03528_),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2636 (.A(_00969_),
    .X(net3160));
 sky130_fd_sc_hd__buf_1 hold2637 (.A(net4404),
    .X(net3161));
 sky130_fd_sc_hd__buf_1 hold2638 (.A(net7494),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(net7757),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net5067),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(net6068),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2641 (.A(_00606_),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2642 (.A(net3473),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(_08227_),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(net4583),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(net7744),
    .X(net3169));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2646 (.A(net4416),
    .X(net3170));
 sky130_fd_sc_hd__clkbuf_2 hold2647 (.A(net4713),
    .X(net3171));
 sky130_fd_sc_hd__clkbuf_2 hold2648 (.A(net4715),
    .X(net3172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(net7742),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net5069),
    .X(net789));
 sky130_fd_sc_hd__buf_1 hold2650 (.A(net4428),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(net3346),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(_03628_),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2653 (.A(_03629_),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(_01012_),
    .X(net3178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(net4436),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(net3956),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(_03245_),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(_03246_),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2659 (.A(_00804_),
    .X(net3183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(net5090),
    .X(net790));
 sky130_fd_sc_hd__buf_1 hold2660 (.A(net4452),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(net4430),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2662 (.A(net3577),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2663 (.A(_08222_),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(net6261),
    .X(net3188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2665 (.A(\rbzero.pov.ready_buffer[5] ),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(_03794_),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(_03795_),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(_01180_),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(net7826),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(net5092),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(net7147),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(_00590_),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(net6305),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(_00592_),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(net3794),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(_08213_),
    .X(net3201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(_00421_),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(\rbzero.row_render.size[7] ),
    .X(net3551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net5056),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(net6079),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(_00579_),
    .X(net3205));
 sky130_fd_sc_hd__clkbuf_2 hold2682 (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(net6153),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(_00417_),
    .X(net3208));
 sky130_fd_sc_hd__buf_1 hold2685 (.A(net4457),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(net4450),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(net3912),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(_02509_),
    .X(net3212));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2689 (.A(_02522_),
    .X(net3213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net5058),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2690 (.A(_02525_),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(_00574_),
    .X(net3215));
 sky130_fd_sc_hd__clkbuf_2 hold2692 (.A(net4718),
    .X(net3216));
 sky130_fd_sc_hd__buf_1 hold2693 (.A(net4454),
    .X(net3217));
 sky130_fd_sc_hd__buf_1 hold2694 (.A(\rbzero.row_render.wall[1] ),
    .X(net3218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(net7319),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(_00522_),
    .X(net3220));
 sky130_fd_sc_hd__buf_1 hold2697 (.A(net7530),
    .X(net3221));
 sky130_fd_sc_hd__clkbuf_2 hold2698 (.A(net684),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(net6099),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net7617),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(_00428_),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(\rbzero.pov.spi_counter[0] ),
    .X(net3225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(_03654_),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(_03656_),
    .X(net3227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(_01029_),
    .X(net3228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(\rbzero.pov.ready_buffer[18] ),
    .X(net3229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(_03824_),
    .X(net3230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(_03825_),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(_01193_),
    .X(net3232));
 sky130_fd_sc_hd__buf_1 hold2709 (.A(net4537),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net4216),
    .X(net795));
 sky130_fd_sc_hd__buf_1 hold2710 (.A(_02406_),
    .X(net3234));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2711 (.A(_02416_),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(_02422_),
    .X(net3236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(net6085),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(_00580_),
    .X(net3239));
 sky130_fd_sc_hd__buf_1 hold2716 (.A(net4466),
    .X(net3240));
 sky130_fd_sc_hd__clkbuf_2 hold2717 (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(net3241));
 sky130_fd_sc_hd__clkbuf_4 hold2718 (.A(_02572_),
    .X(net3242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(_03631_),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(net4325),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(_03632_),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(_01014_),
    .X(net3245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(net6088),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(_00601_),
    .X(net3248));
 sky130_fd_sc_hd__buf_1 hold2725 (.A(net6175),
    .X(net3249));
 sky130_fd_sc_hd__buf_4 hold2726 (.A(_03800_),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(_03943_),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(_03944_),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(_01248_),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_03323_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2730 (.A(\rbzero.spi_registers.buf_sky[0] ),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(_03242_),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2732 (.A(_03243_),
    .X(net3256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2733 (.A(_00802_),
    .X(net3257));
 sky130_fd_sc_hd__buf_1 hold2734 (.A(\rbzero.pov.ready_buffer[61] ),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(_03918_),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(_03919_),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(_01236_),
    .X(net3261));
 sky130_fd_sc_hd__buf_2 hold2738 (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(net6125),
    .X(net3263));
 sky130_fd_sc_hd__buf_2 hold274 (.A(_03324_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2740 (.A(_00419_),
    .X(net3264));
 sky130_fd_sc_hd__clkbuf_2 hold2741 (.A(\rbzero.wall_tracer.mapX[5] ),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(net6142),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(_00620_),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(net5570),
    .X(net3268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(_03783_),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(_03784_),
    .X(net3270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(_01175_),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(net7372),
    .X(net3272));
 sky130_fd_sc_hd__buf_1 hold2749 (.A(_08266_),
    .X(net3273));
 sky130_fd_sc_hd__clkbuf_4 hold275 (.A(_03339_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2750 (.A(net5449),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(net1239),
    .X(net3275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2752 (.A(_03890_),
    .X(net3276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(_03891_),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(_01223_),
    .X(net3278));
 sky130_fd_sc_hd__clkbuf_4 hold2755 (.A(net7256),
    .X(net3279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(_02744_),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2757 (.A(_02745_),
    .X(net3281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2758 (.A(_00597_),
    .X(net3282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(net4926),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net5122),
    .X(net800));
 sky130_fd_sc_hd__buf_1 hold2760 (.A(net7535),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2761 (.A(\rbzero.pov.ready_buffer[54] ),
    .X(net3285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(net639),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(_03903_),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(_03904_),
    .X(net3288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(_01229_),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(net5602),
    .X(net3290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(net1272),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2768 (.A(_03830_),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2769 (.A(_03831_),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(net5131),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2770 (.A(_01196_),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(\rbzero.pov.ready_buffer[23] ),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(net713),
    .X(net3296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(_03834_),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2774 (.A(_03835_),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(_01198_),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(\rbzero.pov.ready_buffer[42] ),
    .X(net3300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(net935),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2778 (.A(_03876_),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2779 (.A(_03877_),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(net5133),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2780 (.A(_01217_),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(\rbzero.pov.ready_buffer[41] ),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2782 (.A(_03874_),
    .X(net3306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(_03875_),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2784 (.A(_01216_),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(\rbzero.pov.ready_buffer[72] ),
    .X(net3309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(net1034),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2787 (.A(_03941_),
    .X(net3311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2788 (.A(_03942_),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2789 (.A(_01247_),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net4998),
    .X(net803));
 sky130_fd_sc_hd__buf_1 hold2790 (.A(net7532),
    .X(net3314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(net7820),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2792 (.A(\rbzero.pov.ready_buffer[9] ),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(net731),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(_03804_),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(_03805_),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(_01184_),
    .X(net3320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2797 (.A(net4482),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(\rbzero.pov.ready_buffer[17] ),
    .X(net3322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2799 (.A(net1251),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(net5000),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2800 (.A(_03821_),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(_03822_),
    .X(net3325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(_01192_),
    .X(net3326));
 sky130_fd_sc_hd__buf_1 hold2803 (.A(net4474),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(net7324),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(_03665_),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(_03666_),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(_01032_),
    .X(net3331));
 sky130_fd_sc_hd__clkbuf_2 hold2808 (.A(net4726),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net5041),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2810 (.A(net6091),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(_00416_),
    .X(net3335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2812 (.A(\rbzero.pov.ready_buffer[40] ),
    .X(net3336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2813 (.A(net845),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2814 (.A(_03872_),
    .X(net3338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(_03873_),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(_01215_),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(\rbzero.pov.spi_buffer[50] ),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(net1343),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2819 (.A(_03894_),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net5043),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2820 (.A(_03895_),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2821 (.A(_01225_),
    .X(net3345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(\rbzero.pov.ready_buffer[16] ),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(net3175),
    .X(net3347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(_03819_),
    .X(net3348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(_03820_),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(_01191_),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(\rbzero.pov.ready_buffer[20] ),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(net1226),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(_03828_),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net5064),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(_03829_),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(_01195_),
    .X(net3355));
 sky130_fd_sc_hd__clkbuf_2 hold2832 (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(net6144),
    .X(net3357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(_00418_),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2835 (.A(\rbzero.pov.ready_buffer[53] ),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(net2892),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(_03900_),
    .X(net3361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2838 (.A(_03901_),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(_01228_),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net5066),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2840 (.A(\rbzero.pov.ready_buffer[44] ),
    .X(net3364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(net2911),
    .X(net3365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(_03881_),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(_03882_),
    .X(net3367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(_01219_),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2845 (.A(net4498),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2847 (.A(net6094),
    .X(net3371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(_00586_),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(net7544),
    .X(net3373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net5196),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(net3968),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(_02983_),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(_02984_),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(_00626_),
    .X(net3377));
 sky130_fd_sc_hd__buf_2 hold2854 (.A(\rbzero.row_render.wall[0] ),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(net6498),
    .X(net3379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(_00521_),
    .X(net3380));
 sky130_fd_sc_hd__buf_1 hold2857 (.A(net4496),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(\rbzero.pov.spi_buffer[70] ),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2859 (.A(net1220),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(net5198),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(_03937_),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2861 (.A(_03938_),
    .X(net3385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2862 (.A(_01245_),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2863 (.A(\rbzero.pov.ready_buffer[14] ),
    .X(net3387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2864 (.A(net949),
    .X(net3388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2865 (.A(_03815_),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2866 (.A(_03816_),
    .X(net3390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2867 (.A(_01189_),
    .X(net3391));
 sky130_fd_sc_hd__clkbuf_2 hold2868 (.A(net7468),
    .X(net3392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2869 (.A(_02392_),
    .X(net3393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net5105),
    .X(net811));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2870 (.A(_02400_),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2871 (.A(_02405_),
    .X(net3395));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2872 (.A(_02408_),
    .X(net3396));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2873 (.A(net3418),
    .X(net3397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2874 (.A(_10060_),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2875 (.A(_10069_),
    .X(net3399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2876 (.A(_10075_),
    .X(net3400));
 sky130_fd_sc_hd__buf_1 hold2877 (.A(_10078_),
    .X(net3401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2878 (.A(net4908),
    .X(net3402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2879 (.A(_04625_),
    .X(net3403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net5107),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2880 (.A(net4948),
    .X(net3404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2882 (.A(_02589_),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2883 (.A(net4693),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2885 (.A(net6101),
    .X(net3409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2886 (.A(_00608_),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2887 (.A(net5687),
    .X(net3411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2888 (.A(net1314),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2889 (.A(_03861_),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net5021),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2890 (.A(_03862_),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2891 (.A(_01210_),
    .X(net3415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2892 (.A(net4927),
    .X(net3416));
 sky130_fd_sc_hd__clkbuf_2 hold2893 (.A(net3066),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2894 (.A(net7475),
    .X(net3418));
 sky130_fd_sc_hd__buf_1 hold2895 (.A(net3397),
    .X(net3419));
 sky130_fd_sc_hd__buf_1 hold2896 (.A(net4529),
    .X(net3420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2897 (.A(\rbzero.pov.ready_buffer[34] ),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2898 (.A(net705),
    .X(net3422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2899 (.A(_03859_),
    .X(net3423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(net5023),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2900 (.A(_03860_),
    .X(net3424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2901 (.A(_01209_),
    .X(net3425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2902 (.A(net7540),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2903 (.A(\rbzero.pov.ready_buffer[6] ),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2904 (.A(net740),
    .X(net3428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2905 (.A(_03796_),
    .X(net3429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2906 (.A(_03797_),
    .X(net3430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2907 (.A(_01181_),
    .X(net3431));
 sky130_fd_sc_hd__buf_1 hold2908 (.A(net4500),
    .X(net3432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2909 (.A(net4512),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net5200),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2910 (.A(net5693),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2911 (.A(net1395),
    .X(net3435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2912 (.A(_03896_),
    .X(net3436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2913 (.A(_03897_),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2914 (.A(_01226_),
    .X(net3438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2915 (.A(\rbzero.pov.ready_buffer[43] ),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2916 (.A(net927),
    .X(net3440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2917 (.A(_03878_),
    .X(net3441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2918 (.A(_03879_),
    .X(net3442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2919 (.A(_01218_),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(net5202),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2921 (.A(_02889_),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2922 (.A(net4760),
    .X(net3446));
 sky130_fd_sc_hd__buf_1 hold2923 (.A(net4506),
    .X(net3447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2924 (.A(\rbzero.pov.ready_buffer[19] ),
    .X(net3448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2925 (.A(net1366),
    .X(net3449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2926 (.A(_03826_),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2927 (.A(_03827_),
    .X(net3451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2928 (.A(_01194_),
    .X(net3452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2929 (.A(\rbzero.pov.ready_buffer[15] ),
    .X(net3453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(net5098),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2930 (.A(_03817_),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2931 (.A(_03818_),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2932 (.A(_01190_),
    .X(net3456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2934 (.A(net6108),
    .X(net3458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2935 (.A(_00602_),
    .X(net3459));
 sky130_fd_sc_hd__buf_1 hold2936 (.A(net4539),
    .X(net3460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2937 (.A(net4925),
    .X(net3461));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2938 (.A(net3283),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2939 (.A(_08211_),
    .X(net3463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(net5100),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2940 (.A(net6205),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2941 (.A(net5663),
    .X(net3465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2942 (.A(net1177),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2943 (.A(_03812_),
    .X(net3467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2944 (.A(_03813_),
    .X(net3468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2945 (.A(_01188_),
    .X(net3469));
 sky130_fd_sc_hd__buf_1 hold2946 (.A(net4569),
    .X(net3470));
 sky130_fd_sc_hd__buf_1 hold2947 (.A(net4565),
    .X(net3471));
 sky130_fd_sc_hd__buf_1 hold2948 (.A(net4557),
    .X(net3472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2949 (.A(net7551),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net5075),
    .X(net819));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2950 (.A(net3166),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2951 (.A(net4853),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2952 (.A(net1175),
    .X(net3476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2953 (.A(_03916_),
    .X(net3477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2954 (.A(_03917_),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2955 (.A(_01235_),
    .X(net3479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2957 (.A(_02902_),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2958 (.A(net4664),
    .X(net3482));
 sky130_fd_sc_hd__buf_1 hold2959 (.A(\rbzero.pov.ready_buffer[58] ),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net5077),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2960 (.A(_03912_),
    .X(net3484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2961 (.A(_03913_),
    .X(net3485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2962 (.A(_01233_),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2963 (.A(net5770),
    .X(net3487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2964 (.A(net1247),
    .X(net3488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2965 (.A(_03914_),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2966 (.A(_03915_),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2967 (.A(_01234_),
    .X(net3491));
 sky130_fd_sc_hd__buf_1 hold2968 (.A(net4578),
    .X(net3492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2969 (.A(net4555),
    .X(net3493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net5109),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2970 (.A(net4527),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2971 (.A(net4855),
    .X(net3495));
 sky130_fd_sc_hd__buf_1 hold2972 (.A(net1411),
    .X(net3496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2973 (.A(_03935_),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2974 (.A(_03936_),
    .X(net3498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2975 (.A(_01244_),
    .X(net3499));
 sky130_fd_sc_hd__buf_1 hold2976 (.A(net4559),
    .X(net3500));
 sky130_fd_sc_hd__buf_1 hold2977 (.A(net4572),
    .X(net3501));
 sky130_fd_sc_hd__buf_1 hold2978 (.A(net4574),
    .X(net3502));
 sky130_fd_sc_hd__buf_1 hold2979 (.A(net4567),
    .X(net3503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(net5111),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2980 (.A(net7467),
    .X(net3504));
 sky130_fd_sc_hd__buf_1 hold2981 (.A(net3392),
    .X(net3505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2982 (.A(net4929),
    .X(net3506));
 sky130_fd_sc_hd__clkbuf_2 hold2983 (.A(_04619_),
    .X(net3507));
 sky130_fd_sc_hd__buf_4 hold2984 (.A(_06390_),
    .X(net3508));
 sky130_fd_sc_hd__buf_1 hold2985 (.A(_08286_),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2986 (.A(_08291_),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2987 (.A(_08292_),
    .X(net3511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2988 (.A(_00464_),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2989 (.A(net4858),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\rbzero.spi_registers.buf_mapdx[3] ),
    .X(net823));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2990 (.A(net1360),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2991 (.A(_03933_),
    .X(net3515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2992 (.A(_03934_),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2993 (.A(_01243_),
    .X(net3517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2994 (.A(net7751),
    .X(net3518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2995 (.A(\rbzero.pov.ready_buffer[37] ),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2996 (.A(_03865_),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2997 (.A(_03866_),
    .X(net3521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2998 (.A(_01212_),
    .X(net3522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2999 (.A(\rbzero.pov.ready_buffer[71] ),
    .X(net3523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net630),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3000 (.A(net725),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3001 (.A(_03939_),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3002 (.A(_03940_),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3003 (.A(_01246_),
    .X(net3527));
 sky130_fd_sc_hd__buf_1 hold3004 (.A(net4585),
    .X(net3528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3005 (.A(net5667),
    .X(net3529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3006 (.A(net1413),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3007 (.A(_03870_),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3008 (.A(_03871_),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3009 (.A(_01214_),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net7313),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3010 (.A(net4025),
    .X(net3534));
 sky130_fd_sc_hd__buf_2 hold3011 (.A(_04819_),
    .X(net3535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3012 (.A(_01612_),
    .X(net3536));
 sky130_fd_sc_hd__buf_1 hold3013 (.A(net4592),
    .X(net3537));
 sky130_fd_sc_hd__buf_2 hold3015 (.A(net6122),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3016 (.A(_08198_),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3017 (.A(_00414_),
    .X(net3541));
 sky130_fd_sc_hd__buf_1 hold3018 (.A(net4590),
    .X(net3542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3019 (.A(net3605),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(net5116),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3020 (.A(_03621_),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3021 (.A(_03622_),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3022 (.A(_01007_),
    .X(net3546));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3023 (.A(\rbzero.pov.ready_buffer[26] ),
    .X(net3547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3024 (.A(_03841_),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3025 (.A(_03842_),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3026 (.A(_01201_),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3028 (.A(_02672_),
    .X(net3552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3029 (.A(net4769),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net5118),
    .X(net827));
 sky130_fd_sc_hd__buf_1 hold3030 (.A(net4612),
    .X(net3554));
 sky130_fd_sc_hd__buf_1 hold3031 (.A(net4598),
    .X(net3555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3032 (.A(\rbzero.pov.spi_buffer[27] ),
    .X(net3556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3033 (.A(net1409),
    .X(net3557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3034 (.A(_03843_),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3035 (.A(_03844_),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(_01202_),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3037 (.A(net4843),
    .X(net3561));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3038 (.A(_03652_),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3039 (.A(net7331),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(net6342),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3040 (.A(_01034_),
    .X(net3564));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3041 (.A(net4604),
    .X(net3565));
 sky130_fd_sc_hd__buf_1 hold3042 (.A(net4596),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3043 (.A(net5790),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3044 (.A(net1316),
    .X(net3568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3045 (.A(_03909_),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3046 (.A(_03910_),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3047 (.A(_01232_),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3048 (.A(\rbzero.pov.ready_buffer[45] ),
    .X(net3572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3049 (.A(net2835),
    .X(net3573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net6344),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3050 (.A(_03883_),
    .X(net3574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3051 (.A(_03884_),
    .X(net3575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3052 (.A(_01220_),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3053 (.A(net7558),
    .X(net3577));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3054 (.A(net3186),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3055 (.A(\rbzero.pov.ready_buffer[49] ),
    .X(net3579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3056 (.A(net2889),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3057 (.A(_03892_),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3058 (.A(_03893_),
    .X(net3582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3059 (.A(_01224_),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_01402_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3060 (.A(net5474),
    .X(net3584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3061 (.A(net1125),
    .X(net3585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3062 (.A(_03802_),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3063 (.A(_03803_),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3064 (.A(_01183_),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3065 (.A(net5611),
    .X(net3589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3066 (.A(net1170),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3067 (.A(_03787_),
    .X(net3591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3068 (.A(_03788_),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3069 (.A(_01177_),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(net5078),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3071 (.A(net6116),
    .X(net3595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3072 (.A(_00582_),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3073 (.A(net5766),
    .X(net3597));
 sky130_fd_sc_hd__buf_1 hold3074 (.A(net1362),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3075 (.A(_03905_),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3076 (.A(_03906_),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3077 (.A(_01230_),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3079 (.A(_02615_),
    .X(net3603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(net5080),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3080 (.A(net4669),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3081 (.A(\rbzero.pov.ready_buffer[11] ),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3082 (.A(net3543),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3083 (.A(_03808_),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3084 (.A(_03809_),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3085 (.A(_01186_),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3086 (.A(\rbzero.pov.ready_buffer[47] ),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3087 (.A(net2922),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3088 (.A(_03887_),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3089 (.A(_03888_),
    .X(net3613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net5094),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3090 (.A(_01222_),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3091 (.A(\rbzero.pov.ready_buffer[4] ),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3092 (.A(_03642_),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3093 (.A(_03643_),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3094 (.A(_01022_),
    .X(net3618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3095 (.A(net5698),
    .X(net3619));
 sky130_fd_sc_hd__buf_1 hold3096 (.A(_04893_),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3097 (.A(_06215_),
    .X(net3621));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3098 (.A(_06258_),
    .X(net3622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3099 (.A(_08285_),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net5096),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3100 (.A(_08287_),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3101 (.A(_08288_),
    .X(net3625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3102 (.A(_00463_),
    .X(net3626));
 sky130_fd_sc_hd__clkbuf_2 hold3103 (.A(net652),
    .X(net3627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3104 (.A(net6149),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3105 (.A(_00429_),
    .X(net3629));
 sky130_fd_sc_hd__buf_1 hold3106 (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(net3630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3107 (.A(_08230_),
    .X(net3631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3108 (.A(_00427_),
    .X(net3632));
 sky130_fd_sc_hd__clkbuf_2 hold3109 (.A(net682),
    .X(net3633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net5160),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3110 (.A(net6135),
    .X(net3634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3111 (.A(_00432_),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3112 (.A(\rbzero.pov.ready_buffer[7] ),
    .X(net3636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3113 (.A(_03798_),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3114 (.A(_03799_),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3115 (.A(_01182_),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3116 (.A(\rbzero.pov.spi_buffer[1] ),
    .X(net3640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3117 (.A(net1237),
    .X(net3641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3118 (.A(_03785_),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3119 (.A(_03786_),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net5162),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3120 (.A(_01176_),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3121 (.A(net5778),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3122 (.A(net1322),
    .X(net3646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3123 (.A(_03907_),
    .X(net3647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3124 (.A(_03908_),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3125 (.A(_01231_),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3126 (.A(net5617),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3127 (.A(net1438),
    .X(net3651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3128 (.A(_03846_),
    .X(net3652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3129 (.A(_03847_),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(net5086),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3130 (.A(_01203_),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3132 (.A(net7333),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3133 (.A(_03608_),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3134 (.A(_01000_),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3135 (.A(net5600),
    .X(net3659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3136 (.A(net1230),
    .X(net3660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3137 (.A(_03810_),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3138 (.A(_03811_),
    .X(net3662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3139 (.A(_01187_),
    .X(net3663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(net5088),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3140 (.A(net5671),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3141 (.A(net1370),
    .X(net3665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3142 (.A(_03863_),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3143 (.A(_03864_),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3144 (.A(_01211_),
    .X(net3668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3145 (.A(\rbzero.pov.spi_buffer[66] ),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3146 (.A(net1241),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3147 (.A(_03929_),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3148 (.A(_03930_),
    .X(net3672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3149 (.A(_01241_),
    .X(net3673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\rbzero.traced_texa[-10] ),
    .X(net839));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3150 (.A(\rbzero.pov.ready_buffer[3] ),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3151 (.A(_03640_),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3152 (.A(_03641_),
    .X(net3676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3153 (.A(_01021_),
    .X(net3677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3154 (.A(net4856),
    .X(net3678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3155 (.A(net1199),
    .X(net3679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3156 (.A(_03931_),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3157 (.A(_03932_),
    .X(net3681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3158 (.A(_01242_),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3159 (.A(net5530),
    .X(net3683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net7514),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3160 (.A(net1224),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3161 (.A(_03806_),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3162 (.A(_03807_),
    .X(net3686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3163 (.A(_01185_),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3165 (.A(_02685_),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3166 (.A(net4698),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3167 (.A(net3779),
    .X(net3691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3168 (.A(_08242_),
    .X(net3692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3169 (.A(net4781),
    .X(net3693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net5215),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3170 (.A(\rbzero.pov.ready_buffer[33] ),
    .X(net3694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3171 (.A(net857),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3172 (.A(_03856_),
    .X(net3696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3173 (.A(_03857_),
    .X(net3697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3174 (.A(_01208_),
    .X(net3698));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3175 (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(net3699));
 sky130_fd_sc_hd__buf_2 hold3176 (.A(_02790_),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3177 (.A(_03647_),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3178 (.A(_03648_),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3179 (.A(_01025_),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(net5217),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3180 (.A(\rbzero.pov.spi_buffer[62] ),
    .X(net3704));
 sky130_fd_sc_hd__buf_1 hold3181 (.A(net1253),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3182 (.A(_03920_),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3183 (.A(_03921_),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3184 (.A(_01237_),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3185 (.A(\rbzero.pov.ready_buffer[32] ),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3186 (.A(_03854_),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3187 (.A(_03855_),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3188 (.A(_01207_),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3189 (.A(\rbzero.pov.ready_buffer[46] ),
    .X(net3713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net5242),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3190 (.A(_03885_),
    .X(net3714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3191 (.A(_03886_),
    .X(net3715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3192 (.A(_01221_),
    .X(net3716));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3193 (.A(net4618),
    .X(net3717));
 sky130_fd_sc_hd__clkbuf_2 hold3194 (.A(net671),
    .X(net3718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3195 (.A(net6151),
    .X(net3719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3196 (.A(_00430_),
    .X(net3720));
 sky130_fd_sc_hd__clkbuf_4 hold3198 (.A(net6133),
    .X(net3722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3199 (.A(_08194_),
    .X(net3723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(net5244),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3200 (.A(_00413_),
    .X(net3724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3202 (.A(net6119),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3203 (.A(_00604_),
    .X(net3727));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3204 (.A(\rbzero.pov.ready_buffer[24] ),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3205 (.A(_03837_),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3206 (.A(_03838_),
    .X(net3730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3207 (.A(_01199_),
    .X(net3731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3208 (.A(net6007),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3209 (.A(_03922_),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net3336),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3210 (.A(_03923_),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3211 (.A(_01238_),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3212 (.A(net5507),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3213 (.A(net1243),
    .X(net3737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3214 (.A(_03792_),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3215 (.A(_03793_),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3216 (.A(_01179_),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3217 (.A(net7524),
    .X(net3741));
 sky130_fd_sc_hd__buf_1 hold3218 (.A(net3058),
    .X(net3742));
 sky130_fd_sc_hd__buf_1 hold3219 (.A(\rbzero.pov.ready_buffer[25] ),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(net4646),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3220 (.A(net7341),
    .X(net3744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3221 (.A(_03606_),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3222 (.A(_00999_),
    .X(net3746));
 sky130_fd_sc_hd__buf_1 hold3223 (.A(net7359),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3224 (.A(_02968_),
    .X(net3748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3225 (.A(_02969_),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3226 (.A(_00621_),
    .X(net3750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3227 (.A(\rbzero.pov.spi_buffer[65] ),
    .X(net3751));
 sky130_fd_sc_hd__buf_1 hold3228 (.A(net1355),
    .X(net3752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3229 (.A(_03927_),
    .X(net3753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net5171),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3230 (.A(_03928_),
    .X(net3754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3231 (.A(_01240_),
    .X(net3755));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3232 (.A(\rbzero.pov.ready_buffer[22] ),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3233 (.A(_03832_),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3234 (.A(_03833_),
    .X(net3758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3235 (.A(_01197_),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3236 (.A(net7352),
    .X(net3760));
 sky130_fd_sc_hd__buf_1 hold3237 (.A(_04813_),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3238 (.A(_05355_),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3239 (.A(_00476_),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(net5173),
    .X(net848));
 sky130_fd_sc_hd__buf_1 hold3240 (.A(\rbzero.pov.ready_buffer[31] ),
    .X(net3764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3241 (.A(_03852_),
    .X(net3765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3242 (.A(_03853_),
    .X(net3766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3243 (.A(_01206_),
    .X(net3767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3245 (.A(net7335),
    .X(net3769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3246 (.A(_03612_),
    .X(net3770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3247 (.A(_01003_),
    .X(net3771));
 sky130_fd_sc_hd__clkbuf_2 hold3248 (.A(net678),
    .X(net3772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3249 (.A(net6147),
    .X(net3773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(net5221),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3250 (.A(_00431_),
    .X(net3774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3251 (.A(\rbzero.pov.ready_buffer[38] ),
    .X(net3775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3252 (.A(_03868_),
    .X(net3776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3253 (.A(_03869_),
    .X(net3777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3254 (.A(_01213_),
    .X(net3778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3255 (.A(net7767),
    .X(net3779));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3256 (.A(net3691),
    .X(net3780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3257 (.A(\rbzero.pov.spi_buffer[30] ),
    .X(net3781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3258 (.A(net1381),
    .X(net3782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3259 (.A(_03850_),
    .X(net3783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net5223),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3260 (.A(_03851_),
    .X(net3784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3261 (.A(_01205_),
    .X(net3785));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3262 (.A(\rbzero.debug_overlay.facingX[-1] ),
    .X(net3786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3263 (.A(_03595_),
    .X(net3787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3264 (.A(_03596_),
    .X(net3788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3265 (.A(_00993_),
    .X(net3789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3267 (.A(net6138),
    .X(net3791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3268 (.A(_00415_),
    .X(net3792));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3269 (.A(net4638),
    .X(net3793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(net4735),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3270 (.A(net4973),
    .X(net3794));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3271 (.A(net3200),
    .X(net3795));
 sky130_fd_sc_hd__clkbuf_2 hold3272 (.A(\rbzero.wall_tracer.rayAddendX[2] ),
    .X(net3796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3273 (.A(net6326),
    .X(net3797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3274 (.A(_00584_),
    .X(net3798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3275 (.A(net5636),
    .X(net3799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3276 (.A(net1306),
    .X(net3800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3277 (.A(_03898_),
    .X(net3801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3278 (.A(_03899_),
    .X(net3802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3279 (.A(_01227_),
    .X(net3803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net4737),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_4 hold3280 (.A(\rbzero.map_rom.b6 ),
    .X(net3804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3281 (.A(net6189),
    .X(net3805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3282 (.A(_00595_),
    .X(net3806));
 sky130_fd_sc_hd__buf_2 hold3283 (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(net3807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3284 (.A(_03644_),
    .X(net3808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3285 (.A(_03645_),
    .X(net3809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3286 (.A(_01023_),
    .X(net3810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3287 (.A(net4847),
    .X(net3811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3288 (.A(net1483),
    .X(net3812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3289 (.A(_03925_),
    .X(net3813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(net5154),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3290 (.A(_03926_),
    .X(net3814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3291 (.A(_01239_),
    .X(net3815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3292 (.A(net5556),
    .X(net3816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3293 (.A(net1328),
    .X(net3817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3294 (.A(_03789_),
    .X(net3818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3295 (.A(_03790_),
    .X(net3819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3296 (.A(_01178_),
    .X(net3820));
 sky130_fd_sc_hd__buf_2 hold3297 (.A(net6154),
    .X(net3821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3298 (.A(_02945_),
    .X(net3822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3299 (.A(_02946_),
    .X(net3823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net5156),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3300 (.A(_00615_),
    .X(net3824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3301 (.A(net7347),
    .X(net3825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3302 (.A(_03668_),
    .X(net3826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3303 (.A(_03669_),
    .X(net3827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3304 (.A(_01033_),
    .X(net3828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3306 (.A(net7337),
    .X(net3830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3307 (.A(_03604_),
    .X(net3831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3308 (.A(_00998_),
    .X(net3832));
 sky130_fd_sc_hd__buf_1 hold3309 (.A(\rbzero.pov.ready_buffer[29] ),
    .X(net3833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net5017),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3310 (.A(_03848_),
    .X(net3834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3311 (.A(_03849_),
    .X(net3835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3312 (.A(_01204_),
    .X(net3836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3313 (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(net3837));
 sky130_fd_sc_hd__clkbuf_4 hold3314 (.A(_05406_),
    .X(net3838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3315 (.A(_03626_),
    .X(net3839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3316 (.A(_03627_),
    .X(net3840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3317 (.A(_01011_),
    .X(net3841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3318 (.A(net5568),
    .X(net3842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3319 (.A(net1339),
    .X(net3843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(net5019),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3320 (.A(_03839_),
    .X(net3844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3321 (.A(_03840_),
    .X(net3845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3322 (.A(_01200_),
    .X(net3846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3324 (.A(net7345),
    .X(net3848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3325 (.A(_03590_),
    .X(net3849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3326 (.A(_00990_),
    .X(net3850));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3327 (.A(net4688),
    .X(net3851));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3328 (.A(net4686),
    .X(net3852));
 sky130_fd_sc_hd__clkbuf_4 hold3329 (.A(net7346),
    .X(net3853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(net3694),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3330 (.A(_02960_),
    .X(net3854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3331 (.A(_02961_),
    .X(net3855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3332 (.A(_00619_),
    .X(net3856));
 sky130_fd_sc_hd__clkbuf_2 hold3333 (.A(\rbzero.debug_overlay.facingY[0] ),
    .X(net3857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3334 (.A(_03617_),
    .X(net3858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3335 (.A(_03618_),
    .X(net3859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3336 (.A(_01005_),
    .X(net3860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3338 (.A(_02832_),
    .X(net3862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3339 (.A(net4711),
    .X(net3863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net4632),
    .X(net858));
 sky130_fd_sc_hd__buf_1 hold3340 (.A(\rbzero.spi_registers.buf_vinf ),
    .X(net3864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3341 (.A(_03299_),
    .X(net3865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3342 (.A(_03300_),
    .X(net3866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3343 (.A(_00836_),
    .X(net3867));
 sky130_fd_sc_hd__buf_2 hold3344 (.A(net4048),
    .X(net3868));
 sky130_fd_sc_hd__clkbuf_2 hold3345 (.A(_04719_),
    .X(net3869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3346 (.A(_04720_),
    .X(net3870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3347 (.A(_00473_),
    .X(net3871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3349 (.A(net7349),
    .X(net3873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net5167),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3350 (.A(_03588_),
    .X(net3874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3351 (.A(_00989_),
    .X(net3875));
 sky130_fd_sc_hd__buf_2 hold3352 (.A(\rbzero.debug_overlay.facingY[10] ),
    .X(net3876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3353 (.A(_03619_),
    .X(net3877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3354 (.A(_03620_),
    .X(net3878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3355 (.A(_01006_),
    .X(net3879));
 sky130_fd_sc_hd__buf_2 hold3356 (.A(net4674),
    .X(net3880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3357 (.A(_06232_),
    .X(net3881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3358 (.A(_02733_),
    .X(net3882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3359 (.A(_02734_),
    .X(net3883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net5169),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3360 (.A(_00594_),
    .X(net3884));
 sky130_fd_sc_hd__buf_1 hold3361 (.A(net7358),
    .X(net3885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3362 (.A(_02980_),
    .X(net3886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3363 (.A(_02981_),
    .X(net3887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3364 (.A(_00625_),
    .X(net3888));
 sky130_fd_sc_hd__buf_1 hold3365 (.A(net7354),
    .X(net3889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3366 (.A(_02971_),
    .X(net3890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3367 (.A(_02972_),
    .X(net3891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3368 (.A(_00622_),
    .X(net3892));
 sky130_fd_sc_hd__clkbuf_4 hold3369 (.A(net6212),
    .X(net3893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(net5139),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3370 (.A(_02741_),
    .X(net3894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3371 (.A(_02742_),
    .X(net3895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3372 (.A(_00596_),
    .X(net3896));
 sky130_fd_sc_hd__buf_2 hold3373 (.A(net6264),
    .X(net3897));
 sky130_fd_sc_hd__buf_1 hold3374 (.A(_03030_),
    .X(net3898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3375 (.A(net6331),
    .X(net3899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3377 (.A(net7343),
    .X(net3901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3378 (.A(_03600_),
    .X(net3902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3379 (.A(_00996_),
    .X(net3903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(net5141),
    .X(net862));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3380 (.A(net7356),
    .X(net3904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3381 (.A(_02977_),
    .X(net3905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3382 (.A(_02978_),
    .X(net3906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3383 (.A(_00624_),
    .X(net3907));
 sky130_fd_sc_hd__clkbuf_2 hold3384 (.A(net6024),
    .X(net3908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3385 (.A(_05331_),
    .X(net3909));
 sky130_fd_sc_hd__buf_1 hold3386 (.A(_05332_),
    .X(net3910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3387 (.A(_00475_),
    .X(net3911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3388 (.A(\rbzero.spi_registers.spi_counter[2] ),
    .X(net3912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3389 (.A(net3211),
    .X(net3913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net4904),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3390 (.A(_02974_),
    .X(net3914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3391 (.A(_02975_),
    .X(net3915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3392 (.A(_00623_),
    .X(net3916));
 sky130_fd_sc_hd__clkbuf_4 hold3393 (.A(net6206),
    .X(net3917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3394 (.A(_02729_),
    .X(net3918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3395 (.A(_02730_),
    .X(net3919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3396 (.A(_00593_),
    .X(net3920));
 sky130_fd_sc_hd__clkbuf_4 hold3397 (.A(net6209),
    .X(net3921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3398 (.A(_02957_),
    .X(net3922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3399 (.A(net6218),
    .X(net3923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net4906),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3400 (.A(_00618_),
    .X(net3924));
 sky130_fd_sc_hd__buf_1 hold3401 (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .X(net3925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3402 (.A(_03466_),
    .X(net3926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3403 (.A(_03467_),
    .X(net3927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3404 (.A(_00952_),
    .X(net3928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3405 (.A(net6040),
    .X(net3929));
 sky130_fd_sc_hd__buf_4 hold3406 (.A(_05827_),
    .X(net3930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3407 (.A(_01262_),
    .X(net3931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3408 (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(net3932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3409 (.A(net3123),
    .X(net3933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(net5282),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3410 (.A(_02998_),
    .X(net3934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3411 (.A(_00631_),
    .X(net3935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3412 (.A(net6219),
    .X(net3936));
 sky130_fd_sc_hd__buf_4 hold3413 (.A(_05828_),
    .X(net3937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3414 (.A(_01263_),
    .X(net3938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3415 (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(net3939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3416 (.A(net3104),
    .X(net3940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3417 (.A(_03000_),
    .X(net3941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3418 (.A(_03003_),
    .X(net3942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3419 (.A(_00633_),
    .X(net3943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net5284),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3420 (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .X(net3944));
 sky130_fd_sc_hd__buf_1 hold3421 (.A(net2841),
    .X(net3945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3422 (.A(_02987_),
    .X(net3946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3423 (.A(_00632_),
    .X(net3947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3424 (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(net3948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3425 (.A(net1607),
    .X(net3949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3426 (.A(_02994_),
    .X(net3950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3427 (.A(_00629_),
    .X(net3951));
 sky130_fd_sc_hd__buf_2 hold3428 (.A(\rbzero.debug_overlay.playerY[5] ),
    .X(net3952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3429 (.A(_03575_),
    .X(net3953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net5123),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3430 (.A(_03576_),
    .X(net3954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3431 (.A(_00984_),
    .X(net3955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3432 (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(net3956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3433 (.A(net3180),
    .X(net3957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3434 (.A(_02996_),
    .X(net3958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3435 (.A(_00630_),
    .X(net3959));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3436 (.A(net7314),
    .X(net3960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3437 (.A(_03464_),
    .X(net3961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3438 (.A(_03465_),
    .X(net3962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3439 (.A(_00951_),
    .X(net3963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net5125),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_4 hold3440 (.A(net6286),
    .X(net3964));
 sky130_fd_sc_hd__clkbuf_4 hold3441 (.A(_05824_),
    .X(net3965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3442 (.A(_03958_),
    .X(net3966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3443 (.A(_01255_),
    .X(net3967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3444 (.A(\rbzero.spi_registers.spi_counter[5] ),
    .X(net3968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3445 (.A(net3374),
    .X(net3969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3446 (.A(_02519_),
    .X(net3970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3447 (.A(net88),
    .X(net3971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3448 (.A(_03459_),
    .X(net3972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3449 (.A(_03462_),
    .X(net3973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net7502),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3450 (.A(_03463_),
    .X(net3974));
 sky130_fd_sc_hd__clkbuf_1 hold3451 (.A(net6313),
    .X(net3975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3452 (.A(_09914_),
    .X(net3976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3453 (.A(_09915_),
    .X(net3977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3454 (.A(_09916_),
    .X(net3978));
 sky130_fd_sc_hd__buf_2 hold3455 (.A(_09917_),
    .X(net3979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3456 (.A(_04127_),
    .X(net3980));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3457 (.A(_04128_),
    .X(net3981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3458 (.A(_01614_),
    .X(net3982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3459 (.A(\rbzero.map_rom.f2 ),
    .X(net3983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net5177),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_4 hold3460 (.A(_06212_),
    .X(net3984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3461 (.A(_02954_),
    .X(net3985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3462 (.A(_00617_),
    .X(net3986));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3463 (.A(net6048),
    .X(net3987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3464 (.A(_04810_),
    .X(net3988));
 sky130_fd_sc_hd__clkbuf_2 hold3465 (.A(_04811_),
    .X(net3989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3466 (.A(_00474_),
    .X(net3990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3467 (.A(net6312),
    .X(net3991));
 sky130_fd_sc_hd__clkbuf_4 hold3468 (.A(net3975),
    .X(net3992));
 sky130_fd_sc_hd__buf_4 hold3469 (.A(_04163_),
    .X(net3993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(net5179),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3470 (.A(net6314),
    .X(net3994));
 sky130_fd_sc_hd__buf_2 hold3471 (.A(\rbzero.debug_overlay.playerX[1] ),
    .X(net3995));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3472 (.A(_04828_),
    .X(net3996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3473 (.A(_02948_),
    .X(net3997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3474 (.A(_02949_),
    .X(net3998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3475 (.A(net6250),
    .X(net3999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3476 (.A(_00616_),
    .X(net4000));
 sky130_fd_sc_hd__buf_2 hold3477 (.A(net5956),
    .X(net4001));
 sky130_fd_sc_hd__buf_4 hold3478 (.A(_05829_),
    .X(net4002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3479 (.A(_01261_),
    .X(net4003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(net5333),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 hold3480 (.A(net7361),
    .X(net4004));
 sky130_fd_sc_hd__clkbuf_2 hold3481 (.A(net4042),
    .X(net4005));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3482 (.A(_05444_),
    .X(net4006));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3483 (.A(_05445_),
    .X(net4007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3484 (.A(_00458_),
    .X(net4008));
 sky130_fd_sc_hd__clkbuf_4 hold3485 (.A(net7364),
    .X(net4009));
 sky130_fd_sc_hd__clkbuf_2 hold3486 (.A(_04613_),
    .X(net4010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3487 (.A(_05348_),
    .X(net4011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3488 (.A(_00477_),
    .X(net4012));
 sky130_fd_sc_hd__clkbuf_2 hold3489 (.A(net6329),
    .X(net4013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(net5335),
    .X(net873));
 sky130_fd_sc_hd__buf_2 hold3490 (.A(_04889_),
    .X(net4014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3491 (.A(_03950_),
    .X(net4015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3492 (.A(_03955_),
    .X(net4016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3493 (.A(_03956_),
    .X(net4017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3494 (.A(_03957_),
    .X(net4018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3495 (.A(_01254_),
    .X(net4019));
 sky130_fd_sc_hd__clkbuf_2 hold3496 (.A(net7307),
    .X(net4020));
 sky130_fd_sc_hd__buf_4 hold3497 (.A(_05817_),
    .X(net4021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3498 (.A(_03963_),
    .X(net4022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3499 (.A(_03964_),
    .X(net4023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(net5127),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3500 (.A(_01256_),
    .X(net4024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3501 (.A(\rbzero.trace_state[0] ),
    .X(net4025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3502 (.A(net3534),
    .X(net4026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3503 (.A(_04627_),
    .X(net4027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3504 (.A(_04126_),
    .X(net4028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3505 (.A(_04129_),
    .X(net4029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3506 (.A(_04130_),
    .X(net4030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3507 (.A(_01611_),
    .X(net4031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3508 (.A(\gpout0.vpos[4] ),
    .X(net4032));
 sky130_fd_sc_hd__clkbuf_4 hold3509 (.A(_04805_),
    .X(net4033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net5129),
    .X(net875));
 sky130_fd_sc_hd__buf_2 hold3510 (.A(_05194_),
    .X(net4034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3511 (.A(_01258_),
    .X(net4035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3512 (.A(net4069),
    .X(net4036));
 sky130_fd_sc_hd__clkbuf_2 hold3513 (.A(_04598_),
    .X(net4037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3514 (.A(_05326_),
    .X(net4038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3515 (.A(_09922_),
    .X(net4039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3516 (.A(_00478_),
    .X(net4040));
 sky130_fd_sc_hd__clkbuf_2 hold3517 (.A(net4051),
    .X(net4041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3518 (.A(_05199_),
    .X(net4042));
 sky130_fd_sc_hd__buf_4 hold3519 (.A(net4005),
    .X(net4043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(net5229),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3520 (.A(_05202_),
    .X(net4044));
 sky130_fd_sc_hd__clkbuf_4 hold3521 (.A(_05531_),
    .X(net4045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3522 (.A(_08278_),
    .X(net4046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3523 (.A(_00459_),
    .X(net4047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3524 (.A(\gpout0.hpos[0] ),
    .X(net4048));
 sky130_fd_sc_hd__buf_2 hold3525 (.A(net3868),
    .X(net4049));
 sky130_fd_sc_hd__clkbuf_2 hold3526 (.A(_04159_),
    .X(net4050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3527 (.A(\gpout0.hpos[7] ),
    .X(net4051));
 sky130_fd_sc_hd__clkbuf_2 hold3528 (.A(net4041),
    .X(net4052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3529 (.A(_04164_),
    .X(net4053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(net5231),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3530 (.A(_09924_),
    .X(net4054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3531 (.A(_09926_),
    .X(net4055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3532 (.A(_09927_),
    .X(net4056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3533 (.A(_00480_),
    .X(net4057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3534 (.A(net4098),
    .X(net4058));
 sky130_fd_sc_hd__clkbuf_4 hold3535 (.A(_04804_),
    .X(net4059));
 sky130_fd_sc_hd__buf_4 hold3536 (.A(_05193_),
    .X(net4060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3537 (.A(_03967_),
    .X(net4061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3538 (.A(_01260_),
    .X(net4062));
 sky130_fd_sc_hd__buf_2 hold3539 (.A(net6190),
    .X(net4063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(net5082),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3540 (.A(_04845_),
    .X(net4064));
 sky130_fd_sc_hd__buf_1 hold3541 (.A(_04859_),
    .X(net4065));
 sky130_fd_sc_hd__clkbuf_4 hold3542 (.A(_05615_),
    .X(net4066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3543 (.A(_08280_),
    .X(net4067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3544 (.A(_00460_),
    .X(net4068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3545 (.A(\gpout0.hpos[6] ),
    .X(net4069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3546 (.A(net4036),
    .X(net4070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3547 (.A(_05327_),
    .X(net4071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3548 (.A(_05334_),
    .X(net4072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3549 (.A(_05352_),
    .X(net4073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net5084),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3550 (.A(_05353_),
    .X(net4074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3551 (.A(_09923_),
    .X(net4075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3552 (.A(net5995),
    .X(net4076));
 sky130_fd_sc_hd__clkbuf_4 hold3553 (.A(_05187_),
    .X(net4077));
 sky130_fd_sc_hd__clkbuf_4 hold3554 (.A(_05779_),
    .X(net4078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3555 (.A(_08282_),
    .X(net4079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3556 (.A(_00462_),
    .X(net4080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3557 (.A(\rbzero.color_sky[4] ),
    .X(net4081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3558 (.A(_05691_),
    .X(net4082));
 sky130_fd_sc_hd__clkbuf_4 hold3559 (.A(_05698_),
    .X(net4083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(net5270),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3560 (.A(_08281_),
    .X(net4084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3561 (.A(_00461_),
    .X(net4085));
 sky130_fd_sc_hd__buf_2 hold3562 (.A(net3480),
    .X(net4086));
 sky130_fd_sc_hd__clkbuf_2 hold3563 (.A(_04646_),
    .X(net4087));
 sky130_fd_sc_hd__clkbuf_4 hold3564 (.A(_08293_),
    .X(net4088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3565 (.A(_00465_),
    .X(net4089));
 sky130_fd_sc_hd__buf_2 hold3566 (.A(net6181),
    .X(net4090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3567 (.A(_04825_),
    .X(net4091));
 sky130_fd_sc_hd__buf_1 hold3568 (.A(_04841_),
    .X(net4092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3569 (.A(_04907_),
    .X(net4093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(net5272),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3570 (.A(_04908_),
    .X(net4094));
 sky130_fd_sc_hd__buf_4 hold3571 (.A(_05203_),
    .X(net4095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3572 (.A(_08277_),
    .X(net4096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3573 (.A(_00457_),
    .X(net4097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3574 (.A(\gpout0.vpos[5] ),
    .X(net4098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3575 (.A(net4058),
    .X(net4099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3576 (.A(_03968_),
    .X(net4100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3577 (.A(_03969_),
    .X(net4101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3578 (.A(\rbzero.vga_sync.vsync ),
    .X(net4102));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3579 (.A(net1451),
    .X(net4103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(net5185),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3580 (.A(_04620_),
    .X(net4104));
 sky130_fd_sc_hd__clkbuf_2 hold3581 (.A(net4218),
    .X(net4105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3582 (.A(_09909_),
    .X(net4106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3583 (.A(_09910_),
    .X(net4107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3584 (.A(\rbzero.row_render.size[10] ),
    .X(net4108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3585 (.A(net694),
    .X(net4109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3586 (.A(net7482),
    .X(net4110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3587 (.A(net700),
    .X(net4111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3588 (.A(net7624),
    .X(net4112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3589 (.A(_00790_),
    .X(net4113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(net5187),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3590 (.A(net602),
    .X(net4114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3591 (.A(net7620),
    .X(net4115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3592 (.A(_00866_),
    .X(net4116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3593 (.A(net699),
    .X(net4117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3594 (.A(net7622),
    .X(net4118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3595 (.A(_00789_),
    .X(net4119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3596 (.A(net599),
    .X(net4120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3597 (.A(net7623),
    .X(net4121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3598 (.A(_00717_),
    .X(net4122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3599 (.A(net605),
    .X(net4123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(net5309),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3600 (.A(net7628),
    .X(net4124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3601 (.A(_00740_),
    .X(net4125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3602 (.A(net620),
    .X(net4126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3603 (.A(net7625),
    .X(net4127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3604 (.A(_00720_),
    .X(net4128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3605 (.A(net608),
    .X(net4129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3606 (.A(net7633),
    .X(net4130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3607 (.A(_00508_),
    .X(net4131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3608 (.A(net696),
    .X(net4132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3609 (.A(net7573),
    .X(net4133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(net5311),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3610 (.A(_00518_),
    .X(net4134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3611 (.A(net683),
    .X(net4135));
 sky130_fd_sc_hd__buf_1 hold3612 (.A(net7537),
    .X(net4136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3613 (.A(_00519_),
    .X(net4137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3614 (.A(net681),
    .X(net4138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3615 (.A(net7491),
    .X(net4139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3616 (.A(net757),
    .X(net4140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3617 (.A(net7471),
    .X(net4141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3618 (.A(net785),
    .X(net4142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3619 (.A(net7637),
    .X(net4143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(net5225),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3620 (.A(_00515_),
    .X(net4144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3621 (.A(net653),
    .X(net4145));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3622 (.A(net7635),
    .X(net4146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3623 (.A(_00507_),
    .X(net4147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3624 (.A(net693),
    .X(net4148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3625 (.A(net7634),
    .X(net4149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3626 (.A(_00718_),
    .X(net4150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3627 (.A(net611),
    .X(net4151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3628 (.A(\rbzero.traced_texa[-4] ),
    .X(net4152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3629 (.A(net7619),
    .X(net4153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(net5227),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3630 (.A(net646),
    .X(net4154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3631 (.A(\rbzero.traced_texa[10] ),
    .X(net4155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3632 (.A(net7555),
    .X(net4156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3633 (.A(net689),
    .X(net4157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3634 (.A(net7486),
    .X(net4158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3635 (.A(net924),
    .X(net4159));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3636 (.A(net7643),
    .X(net4160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3637 (.A(_00516_),
    .X(net4161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3638 (.A(net672),
    .X(net4162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3639 (.A(net7501),
    .X(net4163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(net7638),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3640 (.A(net869),
    .X(net4164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3641 (.A(net7499),
    .X(net4165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3642 (.A(net923),
    .X(net4166));
 sky130_fd_sc_hd__buf_1 hold3643 (.A(net7644),
    .X(net4167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3644 (.A(_00510_),
    .X(net4168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3645 (.A(net674),
    .X(net4169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3646 (.A(net7636),
    .X(net4170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3647 (.A(_00773_),
    .X(net4171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3648 (.A(net1134),
    .X(net4172));
 sky130_fd_sc_hd__buf_1 hold3649 (.A(net7641),
    .X(net4173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net4420),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3650 (.A(_00509_),
    .X(net4174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3651 (.A(net657),
    .X(net4175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3652 (.A(net7642),
    .X(net4176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3653 (.A(_00517_),
    .X(net4177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3654 (.A(net679),
    .X(net4178));
 sky130_fd_sc_hd__buf_1 hold3655 (.A(\rbzero.traced_texa[1] ),
    .X(net4179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3656 (.A(net7553),
    .X(net4180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3657 (.A(net687),
    .X(net4181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3658 (.A(net7497),
    .X(net4182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3659 (.A(net1010),
    .X(net4183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\rbzero.traced_texa[-8] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3660 (.A(net7448),
    .X(net4184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3661 (.A(net1060),
    .X(net4185));
 sky130_fd_sc_hd__buf_1 hold3662 (.A(net7648),
    .X(net4186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3663 (.A(_00514_),
    .X(net4187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3664 (.A(net685),
    .X(net4188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3665 (.A(net7711),
    .X(net4189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3666 (.A(net1072),
    .X(net4190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3667 (.A(net7646),
    .X(net4191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3668 (.A(_00754_),
    .X(net4192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3669 (.A(net1085),
    .X(net4193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(net7507),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3670 (.A(net7649),
    .X(net4194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3671 (.A(_00777_),
    .X(net4195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3672 (.A(net1117),
    .X(net4196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3673 (.A(net7651),
    .X(net4197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3674 (.A(_00683_),
    .X(net4198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3675 (.A(net1143),
    .X(net4199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3676 (.A(net7717),
    .X(net4200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3677 (.A(net1257),
    .X(net4201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3679 (.A(net7506),
    .X(net4203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(net5157),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3680 (.A(net891),
    .X(net4204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3681 (.A(net7654),
    .X(net4205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3682 (.A(_00770_),
    .X(net4206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3683 (.A(net1408),
    .X(net4207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3684 (.A(net7656),
    .X(net4208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3685 (.A(_00769_),
    .X(net4209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3686 (.A(net1216),
    .X(net4210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3687 (.A(net7657),
    .X(net4211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3688 (.A(_00760_),
    .X(net4212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3689 (.A(net1219),
    .X(net4213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(net5159),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3690 (.A(net4222),
    .X(net4214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3691 (.A(_03166_),
    .X(net4215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3692 (.A(_00746_),
    .X(net4216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3693 (.A(net795),
    .X(net4217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3694 (.A(\rbzero.debug_overlay.playerX[-1] ),
    .X(net4218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3695 (.A(net4105),
    .X(net4219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3696 (.A(_00963_),
    .X(net4220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3697 (.A(net1015),
    .X(net4221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3698 (.A(\rbzero.spi_registers.buf_texadd1[16] ),
    .X(net4222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3699 (.A(net4214),
    .X(net4223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(net5235),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3700 (.A(_03382_),
    .X(net4224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3701 (.A(_00893_),
    .X(net4225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3702 (.A(net1592),
    .X(net4226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3703 (.A(net7660),
    .X(net4227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3704 (.A(_00766_),
    .X(net4228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3705 (.A(net1657),
    .X(net4229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3706 (.A(net7721),
    .X(net4230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3707 (.A(net1500),
    .X(net4231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3709 (.A(net7513),
    .X(net4233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net5237),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3710 (.A(net840),
    .X(net4234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3711 (.A(net4242),
    .X(net4235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3712 (.A(_03410_),
    .X(net4236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3713 (.A(_00912_),
    .X(net4237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3714 (.A(net613),
    .X(net4238));
 sky130_fd_sc_hd__clkbuf_2 hold3715 (.A(net7679),
    .X(net4239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3716 (.A(_00494_),
    .X(net4240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3717 (.A(net1423),
    .X(net4241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3718 (.A(\rbzero.spi_registers.buf_texadd2[11] ),
    .X(net4242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3719 (.A(net4235),
    .X(net4243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(net5146),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3720 (.A(_03191_),
    .X(net4244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3721 (.A(_00765_),
    .X(net4245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3722 (.A(net1960),
    .X(net4246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3723 (.A(\rbzero.spi_registers.texadd0[13] ),
    .X(net4247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3724 (.A(net1023),
    .X(net4248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3725 (.A(_00719_),
    .X(net4249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3726 (.A(net1024),
    .X(net4250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3728 (.A(net7516),
    .X(net4252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3729 (.A(net774),
    .X(net4253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(net5148),
    .X(net897));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3730 (.A(net7662),
    .X(net4254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3731 (.A(_00498_),
    .X(net4255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3732 (.A(net1496),
    .X(net4256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3733 (.A(net7669),
    .X(net4257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3734 (.A(_03409_),
    .X(net4258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3735 (.A(_00911_),
    .X(net4259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3736 (.A(net615),
    .X(net4260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3737 (.A(net7668),
    .X(net4261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3738 (.A(_00767_),
    .X(net4262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3739 (.A(net593),
    .X(net4263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(net5189),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3740 (.A(net7845),
    .X(net4264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3741 (.A(net1600),
    .X(net4265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3742 (.A(_00486_),
    .X(net4266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3743 (.A(\rbzero.spi_registers.texadd2[10] ),
    .X(net4267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3744 (.A(net2280),
    .X(net4268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3745 (.A(_00764_),
    .X(net4269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3746 (.A(net2281),
    .X(net4270));
 sky130_fd_sc_hd__buf_1 hold3747 (.A(net7671),
    .X(net4271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3748 (.A(_00495_),
    .X(net4272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3749 (.A(net1190),
    .X(net4273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(net5191),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3750 (.A(net7846),
    .X(net4274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3751 (.A(net1603),
    .X(net4275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3752 (.A(_00483_),
    .X(net4276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3753 (.A(net7942),
    .X(net4277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3754 (.A(net1673),
    .X(net4278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3755 (.A(_00485_),
    .X(net4279));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3756 (.A(net7670),
    .X(net4280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3757 (.A(_00497_),
    .X(net4281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3758 (.A(net1394),
    .X(net4282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3759 (.A(net7723),
    .X(net4283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(net5258),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3760 (.A(net1793),
    .X(net4284));
 sky130_fd_sc_hd__clkbuf_1 hold3761 (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(net4285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3762 (.A(_00512_),
    .X(net4286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3763 (.A(net1101),
    .X(net4287));
 sky130_fd_sc_hd__clkbuf_2 hold3764 (.A(\rbzero.debug_overlay.playerY[-1] ),
    .X(net4288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3765 (.A(_00978_),
    .X(net4289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3766 (.A(net1020),
    .X(net4290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3767 (.A(net7675),
    .X(net4291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3768 (.A(_00768_),
    .X(net4292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3769 (.A(net596),
    .X(net4293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(net5260),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_2 hold3770 (.A(net7379),
    .X(net4294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3771 (.A(_00974_),
    .X(net4295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3772 (.A(net2992),
    .X(net4296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3774 (.A(net7519),
    .X(net4298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3775 (.A(net1012),
    .X(net4299));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3776 (.A(net7427),
    .X(net4300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3777 (.A(_00960_),
    .X(net4301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3778 (.A(net2947),
    .X(net4302));
 sky130_fd_sc_hd__clkbuf_2 hold3779 (.A(net7677),
    .X(net4303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(net5142),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3780 (.A(_00496_),
    .X(net4304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3781 (.A(net1305),
    .X(net4305));
 sky130_fd_sc_hd__clkbuf_2 hold3782 (.A(net7752),
    .X(net4306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3783 (.A(_00956_),
    .X(net4307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3784 (.A(net1158),
    .X(net4308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3785 (.A(net7804),
    .X(net4309));
 sky130_fd_sc_hd__buf_1 hold3786 (.A(net3005),
    .X(net4310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3787 (.A(_08049_),
    .X(net4311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3788 (.A(net7739),
    .X(net4312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3789 (.A(net1304),
    .X(net4313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(net5144),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3790 (.A(net7791),
    .X(net4314));
 sky130_fd_sc_hd__buf_1 hold3791 (.A(net3017),
    .X(net4315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3792 (.A(\rbzero.row_render.size[1] ),
    .X(net4316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3793 (.A(net3016),
    .X(net4317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3794 (.A(net4321),
    .X(net4318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3795 (.A(_00648_),
    .X(net4319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3796 (.A(net644),
    .X(net4320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3797 (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .X(net4321));
 sky130_fd_sc_hd__clkbuf_2 hold3798 (.A(net4318),
    .X(net4322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3799 (.A(_00945_),
    .X(net4323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(net5321),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3800 (.A(net1864),
    .X(net4324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3801 (.A(\rbzero.spi_registers.spi_done ),
    .X(net4325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3802 (.A(net796),
    .X(net4326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3803 (.A(_03357_),
    .X(net4327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3804 (.A(_03391_),
    .X(net4328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3805 (.A(_00921_),
    .X(net4329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3806 (.A(net1539),
    .X(net4330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3807 (.A(net7906),
    .X(net4331));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3808 (.A(net3042),
    .X(net4332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3809 (.A(net7822),
    .X(net4333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net5323),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3810 (.A(net3041),
    .X(net4334));
 sky130_fd_sc_hd__buf_4 hold3811 (.A(net7369),
    .X(net4335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3812 (.A(_00955_),
    .X(net4336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3813 (.A(net735),
    .X(net4337));
 sky130_fd_sc_hd__clkbuf_2 hold3814 (.A(net7731),
    .X(net4338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3815 (.A(_00958_),
    .X(net4339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3816 (.A(net3033),
    .X(net4340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3817 (.A(net7735),
    .X(net4341));
 sky130_fd_sc_hd__buf_1 hold3818 (.A(net2959),
    .X(net4342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3819 (.A(net3551),
    .X(net4343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(net5246),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3820 (.A(net3040),
    .X(net4344));
 sky130_fd_sc_hd__clkbuf_2 hold3821 (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .X(net4345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3822 (.A(_00669_),
    .X(net4346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3823 (.A(net632),
    .X(net4347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3824 (.A(net7479),
    .X(net4348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3825 (.A(net3046),
    .X(net4349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3826 (.A(net7880),
    .X(net4350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3827 (.A(net1189),
    .X(net4351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3828 (.A(net7800),
    .X(net4352));
 sky130_fd_sc_hd__buf_1 hold3829 (.A(net3057),
    .X(net4353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(net5248),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3830 (.A(_08118_),
    .X(net4354));
 sky130_fd_sc_hd__buf_2 hold3831 (.A(net7999),
    .X(net4355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3832 (.A(_00970_),
    .X(net4356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3833 (.A(net2913),
    .X(net4357));
 sky130_fd_sc_hd__clkbuf_4 hold3834 (.A(net7445),
    .X(net4358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3835 (.A(_00977_),
    .X(net4359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3836 (.A(net2916),
    .X(net4360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3837 (.A(net7827),
    .X(net4361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3838 (.A(net3065),
    .X(net4362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(net4790),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3840 (.A(_03584_),
    .X(net4364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3841 (.A(_00986_),
    .X(net4365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3842 (.A(net706),
    .X(net4366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3843 (.A(net7915),
    .X(net4367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3844 (.A(net3103),
    .X(net4368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3845 (.A(net7794),
    .X(net4369));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3846 (.A(net3102),
    .X(net4370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3847 (.A(net7488),
    .X(net4371));
 sky130_fd_sc_hd__buf_1 hold3848 (.A(net3114),
    .X(net4372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3849 (.A(net7816),
    .X(net4373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(net4792),
    .X(net909));
 sky130_fd_sc_hd__buf_1 hold3850 (.A(net3115),
    .X(net4374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3851 (.A(net7900),
    .X(net4375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3852 (.A(net1422),
    .X(net4376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3853 (.A(net7812),
    .X(net4377));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3854 (.A(net3120),
    .X(net4378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3855 (.A(net7892),
    .X(net4379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3856 (.A(net3127),
    .X(net4380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3857 (.A(net7780),
    .X(net4381));
 sky130_fd_sc_hd__buf_1 hold3858 (.A(net3138),
    .X(net4382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3859 (.A(net7737),
    .X(net4383));
 sky130_fd_sc_hd__buf_1 hold386 (.A(net3069),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3860 (.A(net1393),
    .X(net4384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3861 (.A(net7787),
    .X(net4385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3862 (.A(net3143),
    .X(net4386));
 sky130_fd_sc_hd__buf_2 hold3863 (.A(\rbzero.debug_overlay.playerY[2] ),
    .X(net4387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3864 (.A(_00981_),
    .X(net4388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3865 (.A(net670),
    .X(net4389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3866 (.A(\rbzero.row_render.size[8] ),
    .X(net4390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3867 (.A(net2069),
    .X(net4391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3868 (.A(net7450),
    .X(net4392));
 sky130_fd_sc_hd__buf_1 hold3869 (.A(net3148),
    .X(net4393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_03346_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3870 (.A(\rbzero.texV[-2] ),
    .X(net4394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3871 (.A(net711),
    .X(net4395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3872 (.A(_01598_),
    .X(net4396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3873 (.A(net712),
    .X(net4397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3874 (.A(net7594),
    .X(net4398));
 sky130_fd_sc_hd__buf_1 hold3875 (.A(net3149),
    .X(net4399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3876 (.A(net6074),
    .X(net4400));
 sky130_fd_sc_hd__clkbuf_2 hold3877 (.A(net2962),
    .X(net4401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3878 (.A(net7747),
    .X(net4402));
 sky130_fd_sc_hd__buf_1 hold3879 (.A(net3155),
    .X(net4403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(net5351),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3880 (.A(net7839),
    .X(net4404));
 sky130_fd_sc_hd__buf_1 hold3881 (.A(net3161),
    .X(net4405));
 sky130_fd_sc_hd__clkbuf_2 hold3882 (.A(\rbzero.debug_overlay.facingX[10] ),
    .X(net4406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3883 (.A(_03598_),
    .X(net4407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3884 (.A(_00995_),
    .X(net4408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3885 (.A(net928),
    .X(net4409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3886 (.A(net7493),
    .X(net4410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3887 (.A(net3162),
    .X(net4411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3889 (.A(_03609_),
    .X(net4413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(net4805),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3890 (.A(_01001_),
    .X(net4414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3891 (.A(net1099),
    .X(net4415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3892 (.A(net7811),
    .X(net4416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3893 (.A(net3170),
    .X(net4417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3895 (.A(_03610_),
    .X(net4419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3896 (.A(_01002_),
    .X(net4420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3897 (.A(net889),
    .X(net4421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3898 (.A(net7743),
    .X(net4422));
 sky130_fd_sc_hd__buf_1 hold3899 (.A(net3169),
    .X(net4423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(net4807),
    .X(net914));
 sky130_fd_sc_hd__buf_2 hold3900 (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(net4424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3901 (.A(_02533_),
    .X(net4425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3902 (.A(_01636_),
    .X(net4426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3903 (.A(net702),
    .X(net4427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3904 (.A(net7528),
    .X(net4428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3905 (.A(net3174),
    .X(net4429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3906 (.A(net7918),
    .X(net4430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3907 (.A(net3185),
    .X(net4431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3908 (.A(net7741),
    .X(net4432));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3909 (.A(net3173),
    .X(net4433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(net5329),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3910 (.A(net7825),
    .X(net4434));
 sky130_fd_sc_hd__buf_1 hold3911 (.A(net3193),
    .X(net4435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3912 (.A(net7521),
    .X(net4436));
 sky130_fd_sc_hd__buf_1 hold3913 (.A(net3179),
    .X(net4437));
 sky130_fd_sc_hd__buf_2 hold3914 (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(net4438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3915 (.A(_02753_),
    .X(net4439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3916 (.A(_01640_),
    .X(net4440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3917 (.A(net724),
    .X(net4441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3919 (.A(_03585_),
    .X(net4443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(net5331),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3920 (.A(_00987_),
    .X(net4444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3921 (.A(net952),
    .X(net4445));
 sky130_fd_sc_hd__buf_2 hold3922 (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(net4446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3923 (.A(_03624_),
    .X(net4447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3924 (.A(_01009_),
    .X(net4448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3925 (.A(net1299),
    .X(net4449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3926 (.A(net7806),
    .X(net4450));
 sky130_fd_sc_hd__buf_1 hold3927 (.A(net3210),
    .X(net4451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3928 (.A(net7533),
    .X(net4452));
 sky130_fd_sc_hd__buf_1 hold3929 (.A(net3184),
    .X(net4453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(net5164),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3930 (.A(net7838),
    .X(net4454));
 sky130_fd_sc_hd__buf_1 hold3931 (.A(net3217),
    .X(net4455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3932 (.A(_08060_),
    .X(net4456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3933 (.A(net7542),
    .X(net4457));
 sky130_fd_sc_hd__buf_1 hold3934 (.A(net3209),
    .X(net4458));
 sky130_fd_sc_hd__clkbuf_4 hold3935 (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(net4459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3936 (.A(_03646_),
    .X(net4460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3937 (.A(_01024_),
    .X(net4461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3938 (.A(net741),
    .X(net4462));
 sky130_fd_sc_hd__clkbuf_4 hold3939 (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(net4463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(net5166),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3940 (.A(_03630_),
    .X(net4464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3941 (.A(_01013_),
    .X(net4465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3942 (.A(net7523),
    .X(net4466));
 sky130_fd_sc_hd__buf_1 hold3943 (.A(net3240),
    .X(net4467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3944 (.A(\rbzero.texV[4] ),
    .X(net4468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3945 (.A(net1583),
    .X(net4469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3946 (.A(_01604_),
    .X(net4470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3947 (.A(net1584),
    .X(net4471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3948 (.A(net7819),
    .X(net4472));
 sky130_fd_sc_hd__buf_1 hold3949 (.A(net3315),
    .X(net4473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(net5294),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3950 (.A(net7459),
    .X(net4474));
 sky130_fd_sc_hd__buf_1 hold3951 (.A(net3327),
    .X(net4475));
 sky130_fd_sc_hd__buf_2 hold3952 (.A(net4492),
    .X(net4476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3953 (.A(_02539_),
    .X(net4477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3954 (.A(_02540_),
    .X(net4478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3955 (.A(_02544_),
    .X(net4479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3956 (.A(_00577_),
    .X(net4480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3957 (.A(net1077),
    .X(net4481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3958 (.A(net7481),
    .X(net4482));
 sky130_fd_sc_hd__clkbuf_2 hold3959 (.A(net3321),
    .X(net4483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(net5296),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3960 (.A(net7534),
    .X(net4484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3961 (.A(net3284),
    .X(net4485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3962 (.A(net7531),
    .X(net4486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3963 (.A(net3314),
    .X(net4487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3964 (.A(net7529),
    .X(net4488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3965 (.A(net3221),
    .X(net4489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3966 (.A(net7543),
    .X(net4490));
 sky130_fd_sc_hd__buf_1 hold3967 (.A(net3373),
    .X(net4491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3968 (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(net4492));
 sky130_fd_sc_hd__clkbuf_2 hold3969 (.A(net4476),
    .X(net4493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net5101),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3970 (.A(_03625_),
    .X(net4494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3971 (.A(_01010_),
    .X(net4495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3972 (.A(net7453),
    .X(net4496));
 sky130_fd_sc_hd__buf_1 hold3973 (.A(net3381),
    .X(net4497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3974 (.A(net7545),
    .X(net4498));
 sky130_fd_sc_hd__buf_1 hold3975 (.A(net3369),
    .X(net4499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3976 (.A(net7525),
    .X(net4500));
 sky130_fd_sc_hd__buf_1 hold3977 (.A(net3432),
    .X(net4501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3978 (.A(\rbzero.texV[0] ),
    .X(net4502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3979 (.A(net1166),
    .X(net4503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(net5103),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3980 (.A(_01600_),
    .X(net4504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3981 (.A(net1167),
    .X(net4505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3982 (.A(net7522),
    .X(net4506));
 sky130_fd_sc_hd__buf_1 hold3983 (.A(net3447),
    .X(net4507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3984 (.A(net7887),
    .X(net4508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3985 (.A(net2869),
    .X(net4509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3986 (.A(net7539),
    .X(net4510));
 sky130_fd_sc_hd__buf_1 hold3987 (.A(net3426),
    .X(net4511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3988 (.A(net7527),
    .X(net4512));
 sky130_fd_sc_hd__buf_1 hold3989 (.A(net3433),
    .X(net4513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(net7500),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3991 (.A(_03601_),
    .X(net4515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3992 (.A(_00997_),
    .X(net4516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3993 (.A(net714),
    .X(net4517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3994 (.A(net7753),
    .X(net4518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3995 (.A(net1495),
    .X(net4519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3997 (.A(_03586_),
    .X(net4521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3998 (.A(_00988_),
    .X(net4522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3999 (.A(net722),
    .X(net4523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(net7487),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_2 hold4000 (.A(net3630),
    .X(net4524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4001 (.A(_00513_),
    .X(net4525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4002 (.A(net1145),
    .X(net4526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4003 (.A(net7548),
    .X(net4527));
 sky130_fd_sc_hd__buf_1 hold4004 (.A(net3494),
    .X(net4528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4005 (.A(net7814),
    .X(net4529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4006 (.A(net3420),
    .X(net4530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4007 (.A(\rbzero.row_render.side ),
    .X(net4531));
 sky130_fd_sc_hd__buf_2 hold4008 (.A(net3014),
    .X(net4532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4009 (.A(_00482_),
    .X(net4533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(net5135),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4010 (.A(net3015),
    .X(net4534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4011 (.A(net7536),
    .X(net4535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4012 (.A(net3054),
    .X(net4536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4013 (.A(net7538),
    .X(net4537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4014 (.A(net3233),
    .X(net4538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4015 (.A(net7541),
    .X(net4539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4016 (.A(net3460),
    .X(net4540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4017 (.A(\rbzero.texV[1] ),
    .X(net4541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4018 (.A(net1456),
    .X(net4542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4019 (.A(_01601_),
    .X(net4543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(net5137),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4020 (.A(net1457),
    .X(net4544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4021 (.A(\rbzero.texV[-1] ),
    .X(net4545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4022 (.A(net709),
    .X(net4546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4023 (.A(_01599_),
    .X(net4547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4024 (.A(net710),
    .X(net4548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4025 (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(net4549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4026 (.A(_02761_),
    .X(net4550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4027 (.A(_02763_),
    .X(net4551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4028 (.A(_02764_),
    .X(net4552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4029 (.A(_00599_),
    .X(net4553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(net3439),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4030 (.A(net1092),
    .X(net4554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4031 (.A(net7549),
    .X(net4555));
 sky130_fd_sc_hd__buf_1 hold4032 (.A(net3493),
    .X(net4556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4033 (.A(net7408),
    .X(net4557));
 sky130_fd_sc_hd__buf_1 hold4034 (.A(net3472),
    .X(net4558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4035 (.A(net7550),
    .X(net4559));
 sky130_fd_sc_hd__buf_1 hold4036 (.A(net3500),
    .X(net4560));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4037 (.A(\rbzero.debug_overlay.facingX[0] ),
    .X(net4561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4038 (.A(_03597_),
    .X(net4562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4039 (.A(_00994_),
    .X(net4563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(net4408),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4040 (.A(net936),
    .X(net4564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4041 (.A(net7762),
    .X(net4565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4042 (.A(net3471),
    .X(net4566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4043 (.A(net7460),
    .X(net4567));
 sky130_fd_sc_hd__buf_1 hold4044 (.A(net3503),
    .X(net4568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4045 (.A(net7834),
    .X(net4569));
 sky130_fd_sc_hd__buf_1 hold4046 (.A(net3470),
    .X(net4570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4047 (.A(_08252_),
    .X(net4571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4048 (.A(net7490),
    .X(net4572));
 sky130_fd_sc_hd__buf_1 hold4049 (.A(net3501),
    .X(net4573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\rbzero.spi_registers.buf_mapdx[4] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4050 (.A(net7914),
    .X(net4574));
 sky130_fd_sc_hd__buf_1 hold4051 (.A(net3502),
    .X(net4575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4052 (.A(net7750),
    .X(net4576));
 sky130_fd_sc_hd__clkbuf_2 hold4053 (.A(net3518),
    .X(net4577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4054 (.A(net7807),
    .X(net4578));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4055 (.A(net3492),
    .X(net4579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4056 (.A(_08251_),
    .X(net4580));
 sky130_fd_sc_hd__buf_2 hold4057 (.A(net4285),
    .X(net4581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4058 (.A(_08228_),
    .X(net4582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4059 (.A(_00426_),
    .X(net4583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(net636),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4060 (.A(net3168),
    .X(net4584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4061 (.A(net7899),
    .X(net4585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4062 (.A(net3528),
    .X(net4586));
 sky130_fd_sc_hd__buf_2 hold4063 (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(net4587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4064 (.A(_03634_),
    .X(net4588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4065 (.A(_01016_),
    .X(net4589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4066 (.A(net7557),
    .X(net4590));
 sky130_fd_sc_hd__buf_1 hold4067 (.A(net3542),
    .X(net4591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4068 (.A(net7924),
    .X(net4592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4069 (.A(net3537),
    .X(net4593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(net7316),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4070 (.A(net7546),
    .X(net4594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4071 (.A(net3047),
    .X(net4595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4072 (.A(net7560),
    .X(net4596));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4073 (.A(net3566),
    .X(net4597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4074 (.A(net7432),
    .X(net4598));
 sky130_fd_sc_hd__buf_1 hold4075 (.A(net3555),
    .X(net4599));
 sky130_fd_sc_hd__clkbuf_2 hold4076 (.A(\rbzero.debug_overlay.facingY[-1] ),
    .X(net4600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4077 (.A(_03615_),
    .X(net4601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4078 (.A(_01004_),
    .X(net4602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4079 (.A(net2888),
    .X(net4603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(net2252),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4080 (.A(net7902),
    .X(net4604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4081 (.A(net3565),
    .X(net4605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4082 (.A(\rbzero.spi_registers.buf_texadd0[20] ),
    .X(net4606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4083 (.A(net767),
    .X(net4607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4084 (.A(_00873_),
    .X(net4608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4085 (.A(net768),
    .X(net4609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4086 (.A(net7748),
    .X(net4610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4087 (.A(net2955),
    .X(net4611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4088 (.A(net7526),
    .X(net4612));
 sky130_fd_sc_hd__buf_1 hold4089 (.A(net3554),
    .X(net4613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_04334_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4090 (.A(\rbzero.pov.ready_buffer[0] ),
    .X(net4614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4091 (.A(net1587),
    .X(net4615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4092 (.A(_01018_),
    .X(net4616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4093 (.A(net1588),
    .X(net4617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4094 (.A(\rbzero.wall_tracer.stepDistX[8] ),
    .X(net4618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4095 (.A(net3717),
    .X(net4619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4096 (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(net4620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4097 (.A(_02754_),
    .X(net4621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4098 (.A(_04150_),
    .X(net4622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4099 (.A(_01641_),
    .X(net4623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_01442_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4100 (.A(net739),
    .X(net4624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4101 (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(net4625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4102 (.A(_02799_),
    .X(net4626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4103 (.A(_02802_),
    .X(net4627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4104 (.A(net7577),
    .X(net4628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4105 (.A(net3134),
    .X(net4629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4107 (.A(_03583_),
    .X(net4631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4108 (.A(_00985_),
    .X(net4632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4109 (.A(net858),
    .X(net4633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(net3300),
    .X(net935));
 sky130_fd_sc_hd__buf_2 hold4110 (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(net4634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4111 (.A(_03650_),
    .X(net4635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4112 (.A(_01027_),
    .X(net4636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4113 (.A(net732),
    .X(net4637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4114 (.A(net7797),
    .X(net4638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4115 (.A(net3793),
    .X(net4639));
 sky130_fd_sc_hd__buf_2 hold4116 (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(net4640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4117 (.A(_03639_),
    .X(net4641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4118 (.A(_01020_),
    .X(net4642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4119 (.A(net720),
    .X(net4643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(net4563),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4121 (.A(_03593_),
    .X(net4645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4122 (.A(_00992_),
    .X(net4646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4123 (.A(net846),
    .X(net4647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4124 (.A(\rbzero.texV[5] ),
    .X(net4648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4125 (.A(net2776),
    .X(net4649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4126 (.A(_01605_),
    .X(net4650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4127 (.A(net2777),
    .X(net4651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4128 (.A(\rbzero.texV[6] ),
    .X(net4652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4129 (.A(net1504),
    .X(net4653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(net5254),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4130 (.A(_01606_),
    .X(net4654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4131 (.A(net1505),
    .X(net4655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4132 (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(net4656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4133 (.A(_02534_),
    .X(net4657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4134 (.A(_04144_),
    .X(net4658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4135 (.A(_01637_),
    .X(net4659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4136 (.A(net716),
    .X(net4660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4138 (.A(_02877_),
    .X(net4662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4139 (.A(_02892_),
    .X(net4663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(net5256),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4140 (.A(_00610_),
    .X(net4664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4141 (.A(net3482),
    .X(net4665));
 sky130_fd_sc_hd__buf_2 hold4142 (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(net4666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4143 (.A(_02601_),
    .X(net4667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4144 (.A(_02604_),
    .X(net4668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4145 (.A(_00583_),
    .X(net4669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4146 (.A(net3604),
    .X(net4670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4147 (.A(\rbzero.spi_registers.buf_texadd1[20] ),
    .X(net4671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4148 (.A(net1700),
    .X(net4672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4149 (.A(_03387_),
    .X(net4673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(net5317),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4150 (.A(\rbzero.debug_overlay.playerY[1] ),
    .X(net4674));
 sky130_fd_sc_hd__clkbuf_2 hold4151 (.A(net3880),
    .X(net4675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4152 (.A(_00980_),
    .X(net4676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4153 (.A(net641),
    .X(net4677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4154 (.A(\rbzero.texV[9] ),
    .X(net4678));
 sky130_fd_sc_hd__buf_1 hold4155 (.A(net2158),
    .X(net4679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4156 (.A(_01609_),
    .X(net4680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4157 (.A(net2159),
    .X(net4681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4158 (.A(\rbzero.row_render.vinf ),
    .X(net4682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4159 (.A(net3026),
    .X(net4683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(net5319),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4160 (.A(_00665_),
    .X(net4684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4161 (.A(net3027),
    .X(net4685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4162 (.A(net7561),
    .X(net4686));
 sky130_fd_sc_hd__buf_1 hold4163 (.A(net3852),
    .X(net4687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4164 (.A(net7562),
    .X(net4688));
 sky130_fd_sc_hd__buf_1 hold4165 (.A(net3851),
    .X(net4689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4166 (.A(net4771),
    .X(net4690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4167 (.A(_02582_),
    .X(net4691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4168 (.A(_02585_),
    .X(net4692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4169 (.A(_00581_),
    .X(net4693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(net7629),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4170 (.A(net3407),
    .X(net4694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4172 (.A(_02660_),
    .X(net4696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4173 (.A(_02674_),
    .X(net4697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4174 (.A(_00588_),
    .X(net4698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4175 (.A(net3690),
    .X(net4699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4176 (.A(\rbzero.texV[2] ),
    .X(net4700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4177 (.A(net1364),
    .X(net4701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4178 (.A(_01602_),
    .X(net4702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4179 (.A(net1365),
    .X(net4703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(net4803),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4180 (.A(\rbzero.texV[10] ),
    .X(net4704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4181 (.A(net2968),
    .X(net4705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4182 (.A(_01610_),
    .X(net4706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4183 (.A(net2969),
    .X(net4707));
 sky130_fd_sc_hd__clkbuf_2 hold4184 (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(net4708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4185 (.A(_02818_),
    .X(net4709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4186 (.A(_02821_),
    .X(net4710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4187 (.A(_00605_),
    .X(net4711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4188 (.A(net3863),
    .X(net4712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4189 (.A(net7451),
    .X(net4713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(net5274),
    .X(net943));
 sky130_fd_sc_hd__buf_1 hold4190 (.A(net3171),
    .X(net4714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4191 (.A(net7606),
    .X(net4715));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4192 (.A(net3172),
    .X(net4716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4193 (.A(_08257_),
    .X(net4717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4194 (.A(net7840),
    .X(net4718));
 sky130_fd_sc_hd__buf_1 hold4195 (.A(net3216),
    .X(net4719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4197 (.A(_02855_),
    .X(net4721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4198 (.A(_02859_),
    .X(net4722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4199 (.A(_02861_),
    .X(net4723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(net5276),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4200 (.A(_00607_),
    .X(net4724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4201 (.A(net1582),
    .X(net4725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4202 (.A(net7844),
    .X(net4726));
 sky130_fd_sc_hd__buf_1 hold4203 (.A(net3332),
    .X(net4727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4204 (.A(\rbzero.pov.ready_buffer[1] ),
    .X(net4728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4205 (.A(net1623),
    .X(net4729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4206 (.A(_01019_),
    .X(net4730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4207 (.A(net1624),
    .X(net4731));
 sky130_fd_sc_hd__clkbuf_1 hold4208 (.A(net3121),
    .X(net4732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4209 (.A(net7583),
    .X(net4733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net5378),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4210 (.A(net3122),
    .X(net4734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4211 (.A(\rbzero.texV[-3] ),
    .X(net4735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4212 (.A(net851),
    .X(net4736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4213 (.A(_01597_),
    .X(net4737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4214 (.A(net852),
    .X(net4738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4215 (.A(\rbzero.texV[8] ),
    .X(net4739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4216 (.A(net2931),
    .X(net4740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4217 (.A(_01608_),
    .X(net4741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4218 (.A(net2932),
    .X(net4742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4219 (.A(\rbzero.texV[7] ),
    .X(net4743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net5380),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4220 (.A(net2909),
    .X(net4744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4221 (.A(_01607_),
    .X(net4745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4222 (.A(net2910),
    .X(net4746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4223 (.A(\rbzero.pov.ready_buffer[8] ),
    .X(net4747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4224 (.A(net1598),
    .X(net4748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4225 (.A(_01026_),
    .X(net4749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4226 (.A(net1599),
    .X(net4750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4228 (.A(_02638_),
    .X(net4752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4229 (.A(_02642_),
    .X(net4753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(net5355),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4230 (.A(_02644_),
    .X(net4754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4231 (.A(_00585_),
    .X(net4755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4232 (.A(net2000),
    .X(net4756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4234 (.A(_02881_),
    .X(net4758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4235 (.A(_02882_),
    .X(net4759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4236 (.A(_00609_),
    .X(net4760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4237 (.A(net3446),
    .X(net4761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4238 (.A(\rbzero.texV[-4] ),
    .X(net4762));
 sky130_fd_sc_hd__buf_1 hold4239 (.A(net979),
    .X(net4763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(net5357),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4240 (.A(_01596_),
    .X(net4764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4241 (.A(net980),
    .X(net4765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4243 (.A(_02664_),
    .X(net4767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4244 (.A(_02665_),
    .X(net4768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4245 (.A(_00587_),
    .X(net4769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4246 (.A(net3553),
    .X(net4770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4247 (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(net4771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4248 (.A(net4690),
    .X(net4772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4249 (.A(_03633_),
    .X(net4773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net3387),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4250 (.A(_01015_),
    .X(net4774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4251 (.A(\rbzero.pov.ready_buffer[12] ),
    .X(net4775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4252 (.A(net2833),
    .X(net4776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4253 (.A(_01008_),
    .X(net4777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4254 (.A(net2834),
    .X(net4778));
 sky130_fd_sc_hd__buf_4 hold4255 (.A(net680),
    .X(net4779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4256 (.A(_08243_),
    .X(net4780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4257 (.A(_00433_),
    .X(net4781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4258 (.A(net3693),
    .X(net4782));
 sky130_fd_sc_hd__clkbuf_2 hold4259 (.A(net686),
    .X(net4783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(net4495),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4260 (.A(_08226_),
    .X(net4784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4261 (.A(_00425_),
    .X(net4785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4262 (.A(net3056),
    .X(net4786));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4263 (.A(net3006),
    .X(net4787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4264 (.A(_00591_),
    .X(net4788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4265 (.A(net3007),
    .X(net4789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4266 (.A(\rbzero.wall_tracer.rayAddendX[-6] ),
    .X(net4790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4267 (.A(net908),
    .X(net4791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4268 (.A(_01639_),
    .X(net4792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4269 (.A(net909),
    .X(net4793));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold427 (.A(net7647),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4270 (.A(net4836),
    .X(net4794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4271 (.A(_03653_),
    .X(net4795));
 sky130_fd_sc_hd__buf_1 hold4272 (.A(_03655_),
    .X(net4796));
 sky130_fd_sc_hd__buf_1 hold4273 (.A(_03658_),
    .X(net4797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4274 (.A(_01030_),
    .X(net4798));
 sky130_fd_sc_hd__buf_2 hold4275 (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(net4799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4276 (.A(_02759_),
    .X(net4800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4277 (.A(_04153_),
    .X(net4801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4278 (.A(_04154_),
    .X(net4802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4279 (.A(_01643_),
    .X(net4803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(net4444),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4280 (.A(net942),
    .X(net4804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4281 (.A(\rbzero.wall_tracer.rayAddendX[-7] ),
    .X(net4805));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4282 (.A(net913),
    .X(net4806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4283 (.A(_01638_),
    .X(net4807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4284 (.A(net914),
    .X(net4808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4286 (.A(_02689_),
    .X(net4810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4287 (.A(_02690_),
    .X(net4811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4288 (.A(_02691_),
    .X(net4812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4289 (.A(_00589_),
    .X(net4813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(net5597),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4290 (.A(net3045),
    .X(net4814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4292 (.A(_02906_),
    .X(net4816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4293 (.A(_02907_),
    .X(net4817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4294 (.A(_02908_),
    .X(net4818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4295 (.A(_00611_),
    .X(net4819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4296 (.A(net3092),
    .X(net4820));
 sky130_fd_sc_hd__buf_2 hold4297 (.A(net6112),
    .X(net4821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4298 (.A(_06199_),
    .X(net4822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4299 (.A(_06200_),
    .X(net4823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_03680_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4300 (.A(_06201_),
    .X(net4824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4301 (.A(_00386_),
    .X(net4825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4302 (.A(net2389),
    .X(net4826));
 sky130_fd_sc_hd__buf_1 hold4303 (.A(net688),
    .X(net4827));
 sky130_fd_sc_hd__clkbuf_4 hold4304 (.A(_06256_),
    .X(net4828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4305 (.A(_08245_),
    .X(net4829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4306 (.A(_00434_),
    .X(net4830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4307 (.A(net2961),
    .X(net4831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4308 (.A(\rbzero.pov.spi_buffer[63] ),
    .X(net4832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4309 (.A(net1209),
    .X(net4833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(net5599),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4310 (.A(_01099_),
    .X(net4834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4311 (.A(net1210),
    .X(net4835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4312 (.A(\rbzero.pov.sclk_buffer[2] ),
    .X(net4836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4313 (.A(net4794),
    .X(net4837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4314 (.A(_03677_),
    .X(net4838));
 sky130_fd_sc_hd__clkbuf_2 hold4315 (.A(_03757_),
    .X(net4839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4316 (.A(_03764_),
    .X(net4840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4317 (.A(_01101_),
    .X(net4841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4318 (.A(net1356),
    .X(net4842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4319 (.A(\rbzero.pov.ss_buffer[1] ),
    .X(net4843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(net5297),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4320 (.A(net3561),
    .X(net4844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4321 (.A(_03674_),
    .X(net4845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4322 (.A(_01102_),
    .X(net4846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4323 (.A(\rbzero.pov.spi_buffer[64] ),
    .X(net4847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4324 (.A(_01100_),
    .X(net4848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4325 (.A(net4859),
    .X(net4849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4326 (.A(net1282),
    .X(net4850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4327 (.A(_03760_),
    .X(net4851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4328 (.A(_01098_),
    .X(net4852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4329 (.A(\rbzero.pov.spi_buffer[60] ),
    .X(net4853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(net5299),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4330 (.A(_01096_),
    .X(net4854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4331 (.A(\rbzero.pov.spi_buffer[69] ),
    .X(net4855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4332 (.A(\rbzero.pov.spi_buffer[67] ),
    .X(net4856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4333 (.A(_01103_),
    .X(net4857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4334 (.A(\rbzero.pov.spi_buffer[68] ),
    .X(net4858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4335 (.A(\rbzero.pov.spi_buffer[61] ),
    .X(net4859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4336 (.A(\rbzero.pov.spi_buffer[73] ),
    .X(net4860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4337 (.A(net1187),
    .X(net4861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4338 (.A(_01109_),
    .X(net4862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4339 (.A(net1188),
    .X(net4863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net5181),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4340 (.A(\rbzero.pov.spi_counter[2] ),
    .X(net4864));
 sky130_fd_sc_hd__buf_1 hold4341 (.A(net1601),
    .X(net4865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4342 (.A(_01031_),
    .X(net4866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4343 (.A(\rbzero.pov.spi_buffer[72] ),
    .X(net4867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4344 (.A(net1508),
    .X(net4868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4345 (.A(_01108_),
    .X(net4869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4346 (.A(net1509),
    .X(net4870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4348 (.A(_00613_),
    .X(net4872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4349 (.A(net3086),
    .X(net4873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net5183),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 hold4350 (.A(net6158),
    .X(net4874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4351 (.A(_09958_),
    .X(net4875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4352 (.A(_09959_),
    .X(net4876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4353 (.A(_09961_),
    .X(net4877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4354 (.A(_00523_),
    .X(net4878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4355 (.A(net2808),
    .X(net4879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4356 (.A(\rbzero.pov.spi_buffer[71] ),
    .X(net4880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4357 (.A(net1302),
    .X(net4881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4358 (.A(_01107_),
    .X(net4882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4359 (.A(\rbzero.pov.sclk_buffer[1] ),
    .X(net4883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(net5374),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4360 (.A(net2122),
    .X(net4884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4361 (.A(_01106_),
    .X(net4885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4362 (.A(\rbzero.wall_tracer.mapY[8] ),
    .X(net4886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4363 (.A(net1130),
    .X(net4887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4364 (.A(_00388_),
    .X(net4888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4365 (.A(net1131),
    .X(net4889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4366 (.A(\gpout0.hpos[1] ),
    .X(net4890));
 sky130_fd_sc_hd__clkbuf_4 hold4367 (.A(net2986),
    .X(net4891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4368 (.A(\rbzero.debug_overlay.playerY[-7] ),
    .X(net4892));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4369 (.A(net2940),
    .X(net4893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(net5376),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4370 (.A(_00972_),
    .X(net4894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4371 (.A(net2941),
    .X(net4895));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4372 (.A(net6288),
    .X(net4896));
 sky130_fd_sc_hd__clkbuf_2 hold4373 (.A(_06227_),
    .X(net4897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4374 (.A(_06261_),
    .X(net4898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4375 (.A(_06267_),
    .X(net4899));
 sky130_fd_sc_hd__clkbuf_2 hold4376 (.A(_06268_),
    .X(net4900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4377 (.A(_09963_),
    .X(net4901));
 sky130_fd_sc_hd__clkbuf_4 hold4378 (.A(_09964_),
    .X(net4902));
 sky130_fd_sc_hd__buf_4 hold4379 (.A(_10039_),
    .X(net4903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(net5359),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4380 (.A(\rbzero.wall_tracer.rayAddendY[-7] ),
    .X(net4904));
 sky130_fd_sc_hd__buf_1 hold4381 (.A(net863),
    .X(net4905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4382 (.A(_01642_),
    .X(net4906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4383 (.A(net864),
    .X(net4907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4384 (.A(net7353),
    .X(net4908));
 sky130_fd_sc_hd__buf_2 hold4385 (.A(net3402),
    .X(net4909));
 sky130_fd_sc_hd__buf_1 hold4386 (.A(_04629_),
    .X(net4910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4387 (.A(_06203_),
    .X(net4911));
 sky130_fd_sc_hd__buf_1 hold4388 (.A(net6269),
    .X(net4912));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold4389 (.A(_06245_),
    .X(net4913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(net5361),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4390 (.A(_06347_),
    .X(net4914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4391 (.A(_06348_),
    .X(net4915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4392 (.A(_06359_),
    .X(net4916));
 sky130_fd_sc_hd__buf_1 hold4393 (.A(_06383_),
    .X(net4917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4394 (.A(_06389_),
    .X(net4918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4395 (.A(_06391_),
    .X(net4919));
 sky130_fd_sc_hd__clkbuf_2 hold4396 (.A(_02337_),
    .X(net4920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4397 (.A(\rbzero.wall_tracer.mapX[8] ),
    .X(net4921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4398 (.A(net1249),
    .X(net4922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4399 (.A(_00525_),
    .X(net4923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(net5313),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4400 (.A(net1250),
    .X(net4924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4401 (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .X(net4925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4402 (.A(net3461),
    .X(net4926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4403 (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .X(net4927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4404 (.A(net3416),
    .X(net4928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4405 (.A(\rbzero.trace_state[1] ),
    .X(net4929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4406 (.A(net3506),
    .X(net4930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4407 (.A(_04626_),
    .X(net4931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4408 (.A(_08247_),
    .X(net4932));
 sky130_fd_sc_hd__clkbuf_2 hold4409 (.A(_08248_),
    .X(net4933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net5315),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4410 (.A(_08267_),
    .X(net4934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4411 (.A(\rbzero.traced_texa[3] ),
    .X(net4935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4412 (.A(net1144),
    .X(net4936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4413 (.A(_04088_),
    .X(net4937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4414 (.A(_04092_),
    .X(net4938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4415 (.A(_01603_),
    .X(net4939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4416 (.A(net1887),
    .X(net4940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4417 (.A(\gpout2.clk_div[0] ),
    .X(net4941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4418 (.A(net654),
    .X(net4942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4419 (.A(_01646_),
    .X(net4943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net5341),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4420 (.A(\gpout5.clk_div[0] ),
    .X(net4944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4421 (.A(net666),
    .X(net4945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4422 (.A(_01587_),
    .X(net4946));
 sky130_fd_sc_hd__buf_4 hold4423 (.A(_04636_),
    .X(net4947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4424 (.A(_00000_),
    .X(net4948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4425 (.A(net3404),
    .X(net4949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4426 (.A(\gpout0.clk_div[0] ),
    .X(net4950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4427 (.A(net658),
    .X(net4951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4428 (.A(_01634_),
    .X(net4952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(net5343),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_4 hold4430 (.A(_08661_),
    .X(net4954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4431 (.A(\gpout1.clk_div[0] ),
    .X(net4955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4432 (.A(net660),
    .X(net4956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4433 (.A(_01644_),
    .X(net4957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4434 (.A(\gpout4.clk_div[0] ),
    .X(net4958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4435 (.A(net662),
    .X(net4959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4436 (.A(_01650_),
    .X(net4960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4437 (.A(\rbzero.hsync ),
    .X(net4961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4438 (.A(net650),
    .X(net4962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4439 (.A(_01621_),
    .X(net4963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\rbzero.spi_registers.buf_texadd0[12] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4440 (.A(\gpout3.clk_div[0] ),
    .X(net4964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4441 (.A(net664),
    .X(net4965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4442 (.A(_01648_),
    .X(net4966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4443 (.A(\rbzero.pov.spi_counter[6] ),
    .X(net4967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4444 (.A(net690),
    .X(net4968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4445 (.A(_01035_),
    .X(net4969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4446 (.A(net691),
    .X(net4970));
 sky130_fd_sc_hd__buf_1 hold4447 (.A(\gpout0.vpos[6] ),
    .X(net4971));
 sky130_fd_sc_hd__clkbuf_4 hold4448 (.A(_04801_),
    .X(net4972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4449 (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .X(net4973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(net609),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4450 (.A(\rbzero.texV[-10] ),
    .X(net4974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4451 (.A(net707),
    .X(net4975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4452 (.A(_01590_),
    .X(net4976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4453 (.A(net708),
    .X(net4977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4454 (.A(\rbzero.spi_registers.texadd3[21] ),
    .X(net4978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4455 (.A(net775),
    .X(net4979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4456 (.A(_00799_),
    .X(net4980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4457 (.A(net776),
    .X(net4981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4458 (.A(\rbzero.spi_registers.texadd1[9] ),
    .X(net4982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4459 (.A(net779),
    .X(net4983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net7339),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4460 (.A(_00739_),
    .X(net4984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4461 (.A(net780),
    .X(net4985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4462 (.A(\rbzero.texV[-11] ),
    .X(net4986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4463 (.A(net717),
    .X(net4987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4464 (.A(_01589_),
    .X(net4988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4465 (.A(net718),
    .X(net4989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4466 (.A(\rbzero.spi_registers.buf_texadd0[17] ),
    .X(net4990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4467 (.A(net736),
    .X(net4991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4468 (.A(_00870_),
    .X(net4992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4469 (.A(net737),
    .X(net4993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net5266),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4470 (.A(\rbzero.spi_registers.texadd1[8] ),
    .X(net4994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4471 (.A(net753),
    .X(net4995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4472 (.A(_00738_),
    .X(net4996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4473 (.A(net754),
    .X(net4997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4474 (.A(\rbzero.spi_registers.texadd3[10] ),
    .X(net4998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4475 (.A(net803),
    .X(net4999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4476 (.A(_00788_),
    .X(net5000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4477 (.A(net804),
    .X(net5001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4478 (.A(\rbzero.spi_registers.texadd3[17] ),
    .X(net5002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4479 (.A(net771),
    .X(net5003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(net5268),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4480 (.A(_00795_),
    .X(net5004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4481 (.A(net772),
    .X(net5005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4482 (.A(\rbzero.spi_registers.texadd1[18] ),
    .X(net5006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4483 (.A(net763),
    .X(net5007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4484 (.A(_00748_),
    .X(net5008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4485 (.A(net764),
    .X(net5009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4486 (.A(\rbzero.spi_registers.buf_texadd0[15] ),
    .X(net5010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4487 (.A(net742),
    .X(net5011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4488 (.A(_00868_),
    .X(net5012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4489 (.A(\rbzero.spi_registers.buf_mapdy[3] ),
    .X(net5013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(net5278),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4490 (.A(net755),
    .X(net5014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4491 (.A(_00846_),
    .X(net5015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4492 (.A(net756),
    .X(net5016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4493 (.A(\rbzero.spi_registers.texadd3[16] ),
    .X(net5017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4494 (.A(net855),
    .X(net5018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4495 (.A(_00794_),
    .X(net5019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4496 (.A(net856),
    .X(net5020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4497 (.A(\rbzero.spi_registers.texadd1[7] ),
    .X(net5021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4498 (.A(net813),
    .X(net5022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4499 (.A(_00737_),
    .X(net5023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(net5280),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4500 (.A(net814),
    .X(net5024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4501 (.A(\rbzero.spi_registers.texadd1[6] ),
    .X(net5025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4502 (.A(net765),
    .X(net5026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4503 (.A(_00736_),
    .X(net5027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4504 (.A(net766),
    .X(net5028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4505 (.A(\rbzero.spi_registers.buf_texadd0[10] ),
    .X(net5029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4506 (.A(net703),
    .X(net5030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4507 (.A(_00863_),
    .X(net5031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4508 (.A(net704),
    .X(net5032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4509 (.A(\rbzero.spi_registers.buf_texadd0[21] ),
    .X(net5033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net5345),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4510 (.A(net781),
    .X(net5034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4511 (.A(_00874_),
    .X(net5035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4512 (.A(net782),
    .X(net5036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4513 (.A(\rbzero.spi_registers.buf_texadd0[23] ),
    .X(net5037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4514 (.A(net783),
    .X(net5038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4515 (.A(_00876_),
    .X(net5039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4516 (.A(net784),
    .X(net5040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4517 (.A(\rbzero.spi_registers.texadd0[20] ),
    .X(net5041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4518 (.A(net805),
    .X(net5042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4519 (.A(_00726_),
    .X(net5043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(net5347),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4520 (.A(\rbzero.spi_registers.buf_othery[3] ),
    .X(net5044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4521 (.A(net786),
    .X(net5045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4522 (.A(_00828_),
    .X(net5046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4523 (.A(net787),
    .X(net5047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4524 (.A(\rbzero.pov.spi_buffer[32] ),
    .X(net5048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4525 (.A(net1274),
    .X(net5049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4526 (.A(_01068_),
    .X(net5050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4527 (.A(net1275),
    .X(net5051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4528 (.A(\rbzero.spi_registers.texadd1[15] ),
    .X(net5052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4529 (.A(net777),
    .X(net5053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(net5419),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4530 (.A(_00745_),
    .X(net5054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4531 (.A(net778),
    .X(net5055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4532 (.A(\rbzero.spi_registers.buf_texadd0[4] ),
    .X(net5056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4533 (.A(net792),
    .X(net5057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4534 (.A(_00857_),
    .X(net5058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4535 (.A(net793),
    .X(net5059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4536 (.A(\rbzero.spi_registers.buf_texadd0[16] ),
    .X(net5060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4537 (.A(net758),
    .X(net5061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4538 (.A(_00869_),
    .X(net5062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4539 (.A(net759),
    .X(net5063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net5421),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4540 (.A(\rbzero.spi_registers.buf_mapdy[0] ),
    .X(net5064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4541 (.A(net807),
    .X(net5065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4542 (.A(_00843_),
    .X(net5066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4543 (.A(\rbzero.color_sky[3] ),
    .X(net5067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4544 (.A(net788),
    .X(net5068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4545 (.A(_00691_),
    .X(net5069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4546 (.A(net789),
    .X(net5070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4547 (.A(\rbzero.spi_registers.buf_texadd0[1] ),
    .X(net5071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4548 (.A(net769),
    .X(net5072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4549 (.A(_00854_),
    .X(net5073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net4762),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4550 (.A(net770),
    .X(net5074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4551 (.A(\rbzero.spi_registers.texadd0[21] ),
    .X(net5075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4552 (.A(net819),
    .X(net5076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4553 (.A(_00727_),
    .X(net5077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4554 (.A(\rbzero.spi_registers.buf_mapdy[5] ),
    .X(net5078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4555 (.A(net831),
    .X(net5079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4556 (.A(_00848_),
    .X(net5080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4557 (.A(net832),
    .X(net5081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4558 (.A(\rbzero.spi_registers.texadd1[14] ),
    .X(net5082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4559 (.A(net878),
    .X(net5083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(net4764),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4560 (.A(_00744_),
    .X(net5084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4561 (.A(net879),
    .X(net5085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4562 (.A(\rbzero.spi_registers.buf_texadd0[0] ),
    .X(net5086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4563 (.A(net837),
    .X(net5087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4564 (.A(_00853_),
    .X(net5088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4565 (.A(net838),
    .X(net5089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4566 (.A(\rbzero.spi_registers.texadd3[23] ),
    .X(net5090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4567 (.A(net790),
    .X(net5091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4568 (.A(_00801_),
    .X(net5092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4569 (.A(net791),
    .X(net5093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(net5366),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4570 (.A(\rbzero.spi_registers.buf_texadd0[22] ),
    .X(net5094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4571 (.A(net833),
    .X(net5095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4572 (.A(_00875_),
    .X(net5096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4573 (.A(net834),
    .X(net5097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4574 (.A(\rbzero.spi_registers.buf_mapdx[5] ),
    .X(net5098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4575 (.A(net817),
    .X(net5099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4576 (.A(_00842_),
    .X(net5100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4577 (.A(\rbzero.spi_registers.texadd3[9] ),
    .X(net5101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4578 (.A(net921),
    .X(net5102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4579 (.A(_00787_),
    .X(net5103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net5368),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4580 (.A(net922),
    .X(net5104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4581 (.A(\rbzero.spi_registers.texadd3[20] ),
    .X(net5105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4582 (.A(net811),
    .X(net5106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4583 (.A(_00798_),
    .X(net5107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4584 (.A(net812),
    .X(net5108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4585 (.A(\rbzero.spi_registers.buf_otherx[3] ),
    .X(net5109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4586 (.A(net821),
    .X(net5110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4587 (.A(_00823_),
    .X(net5111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4588 (.A(net822),
    .X(net5112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4589 (.A(\rbzero.pov.spi_buffer[31] ),
    .X(net5113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(net5290),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4590 (.A(net1278),
    .X(net5114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4591 (.A(_01067_),
    .X(net5115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4592 (.A(\rbzero.color_sky[1] ),
    .X(net5116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4593 (.A(net826),
    .X(net5117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4594 (.A(_00689_),
    .X(net5118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4595 (.A(net827),
    .X(net5119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4596 (.A(\rbzero.spi_registers.buf_texadd0[11] ),
    .X(net5120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4597 (.A(net603),
    .X(net5121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4598 (.A(_00864_),
    .X(net5122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4599 (.A(\rbzero.spi_registers.buf_othery[2] ),
    .X(net5123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(net5292),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4600 (.A(net867),
    .X(net5124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4601 (.A(_00827_),
    .X(net5125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4602 (.A(net868),
    .X(net5126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4603 (.A(\rbzero.spi_registers.texadd0[6] ),
    .X(net5127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4604 (.A(net874),
    .X(net5128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4605 (.A(_00712_),
    .X(net5129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4606 (.A(net875),
    .X(net5130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4607 (.A(\rbzero.spi_registers.buf_mapdx[0] ),
    .X(net5131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4608 (.A(net801),
    .X(net5132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4609 (.A(_00837_),
    .X(net5133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net5470),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4610 (.A(net802),
    .X(net5134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4611 (.A(\rbzero.spi_registers.texadd1[5] ),
    .X(net5135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4612 (.A(net925),
    .X(net5136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4613 (.A(_00735_),
    .X(net5137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4614 (.A(net926),
    .X(net5138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4615 (.A(\rbzero.spi_registers.buf_texadd0[18] ),
    .X(net5139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4616 (.A(net861),
    .X(net5140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4617 (.A(_00871_),
    .X(net5141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4618 (.A(\rbzero.spi_registers.texadd3[15] ),
    .X(net5142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4619 (.A(net902),
    .X(net5143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(net5472),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4620 (.A(_00793_),
    .X(net5144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4621 (.A(net903),
    .X(net5145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4622 (.A(\rbzero.spi_registers.texadd3[1] ),
    .X(net5146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4623 (.A(net896),
    .X(net5147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4624 (.A(_00779_),
    .X(net5148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4625 (.A(net897),
    .X(net5149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4626 (.A(\rbzero.color_floor[4] ),
    .X(net5150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4627 (.A(net987),
    .X(net5151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4628 (.A(_00698_),
    .X(net5152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4629 (.A(net988),
    .X(net5153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(net5150),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4630 (.A(\rbzero.spi_registers.buf_mapdx[2] ),
    .X(net5154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4631 (.A(net853),
    .X(net5155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4632 (.A(_00839_),
    .X(net5156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4633 (.A(\rbzero.spi_registers.texadd1[20] ),
    .X(net5157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4634 (.A(net892),
    .X(net5158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4635 (.A(_00750_),
    .X(net5159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4636 (.A(\rbzero.spi_registers.buf_texadd0[19] ),
    .X(net5160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4637 (.A(net835),
    .X(net5161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4638 (.A(_00872_),
    .X(net5162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4639 (.A(net836),
    .X(net5163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(net5152),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4640 (.A(\rbzero.spi_registers.texadd0[17] ),
    .X(net5164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4641 (.A(net917),
    .X(net5165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4642 (.A(_00723_),
    .X(net5166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4643 (.A(\rbzero.texV[-7] ),
    .X(net5167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4644 (.A(net859),
    .X(net5168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4645 (.A(_01593_),
    .X(net5169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4646 (.A(net860),
    .X(net5170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4647 (.A(\rbzero.spi_registers.texadd0[10] ),
    .X(net5171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4648 (.A(net847),
    .X(net5172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4649 (.A(_00716_),
    .X(net5173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(net5262),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4650 (.A(net5494),
    .X(net5174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4651 (.A(net1470),
    .X(net5175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4652 (.A(_01066_),
    .X(net5176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4653 (.A(\rbzero.spi_registers.buf_vshift[3] ),
    .X(net5177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4654 (.A(net870),
    .X(net5178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4655 (.A(_00833_),
    .X(net5179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4656 (.A(net871),
    .X(net5180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4657 (.A(\rbzero.spi_registers.texadd1[12] ),
    .X(net5181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4658 (.A(net958),
    .X(net5182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4659 (.A(_00742_),
    .X(net5183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net5264),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4660 (.A(net959),
    .X(net5184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4661 (.A(\rbzero.spi_registers.buf_mapdy[4] ),
    .X(net5185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4662 (.A(net882),
    .X(net5186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4663 (.A(_00847_),
    .X(net5187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4664 (.A(net883),
    .X(net5188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4665 (.A(\rbzero.spi_registers.buf_mapdx[1] ),
    .X(net5189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4666 (.A(net898),
    .X(net5190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4667 (.A(_00838_),
    .X(net5191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4668 (.A(\rbzero.pov.spi_buffer[44] ),
    .X(net5192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4669 (.A(net1290),
    .X(net5193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net5301),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4670 (.A(_01080_),
    .X(net5194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4671 (.A(net1291),
    .X(net5195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4672 (.A(\rbzero.spi_registers.buf_texadd0[6] ),
    .X(net5196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4673 (.A(net809),
    .X(net5197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4674 (.A(_00859_),
    .X(net5198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4675 (.A(net810),
    .X(net5199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4676 (.A(\rbzero.spi_registers.buf_texadd0[7] ),
    .X(net5200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4677 (.A(net815),
    .X(net5201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4678 (.A(_00860_),
    .X(net5202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4679 (.A(net816),
    .X(net5203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(net5303),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4680 (.A(\rbzero.pov.spi_buffer[46] ),
    .X(net5204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4681 (.A(net1375),
    .X(net5205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4682 (.A(_01082_),
    .X(net5206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4683 (.A(net1376),
    .X(net5207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4684 (.A(\rbzero.pov.spi_buffer[9] ),
    .X(net5208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4685 (.A(net1245),
    .X(net5209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4686 (.A(_01045_),
    .X(net5210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4687 (.A(\rbzero.pov.spi_buffer[43] ),
    .X(net5211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4688 (.A(net1228),
    .X(net5212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4689 (.A(_01079_),
    .X(net5213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net5370),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4690 (.A(net1229),
    .X(net5214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4691 (.A(\rbzero.spi_registers.buf_mapdy[2] ),
    .X(net5215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4692 (.A(net841),
    .X(net5216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4693 (.A(_00845_),
    .X(net5217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4694 (.A(\rbzero.pov.spi_buffer[47] ),
    .X(net5218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4695 (.A(net1324),
    .X(net5219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4696 (.A(_01083_),
    .X(net5220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4697 (.A(\rbzero.spi_registers.buf_texadd0[8] ),
    .X(net5221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4698 (.A(net849),
    .X(net5222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4699 (.A(_00861_),
    .X(net5223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net5372),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4700 (.A(net850),
    .X(net5224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4701 (.A(\rbzero.spi_registers.buf_texadd0[2] ),
    .X(net5225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4702 (.A(net886),
    .X(net5226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4703 (.A(_00855_),
    .X(net5227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4704 (.A(net887),
    .X(net5228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4705 (.A(\rbzero.spi_registers.texadd0[7] ),
    .X(net5229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4706 (.A(net876),
    .X(net5230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4707 (.A(_00713_),
    .X(net5231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4708 (.A(\rbzero.pov.spi_buffer[33] ),
    .X(net5232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4709 (.A(net1433),
    .X(net5233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(net6358),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4710 (.A(_01069_),
    .X(net5234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4711 (.A(\rbzero.spi_registers.buf_texadd0[3] ),
    .X(net5235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4712 (.A(net894),
    .X(net5236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4713 (.A(_00856_),
    .X(net5237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4714 (.A(net895),
    .X(net5238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4715 (.A(\rbzero.pov.spi_buffer[45] ),
    .X(net5239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4716 (.A(net1270),
    .X(net5240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4717 (.A(_01081_),
    .X(net5241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4718 (.A(\rbzero.spi_registers.buf_mapdyw[0] ),
    .X(net5242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4719 (.A(net843),
    .X(net5243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(net6360),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4720 (.A(_00851_),
    .X(net5244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4721 (.A(net844),
    .X(net5245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4722 (.A(\rbzero.spi_registers.buf_vshift[0] ),
    .X(net5246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4723 (.A(net906),
    .X(net5247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4724 (.A(_00830_),
    .X(net5248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4725 (.A(net907),
    .X(net5249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4726 (.A(\rbzero.pov.spi_buffer[6] ),
    .X(net5250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4727 (.A(net1232),
    .X(net5251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4728 (.A(_01042_),
    .X(net5252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4729 (.A(net1233),
    .X(net5253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_01542_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4730 (.A(\rbzero.spi_registers.buf_otherx[0] ),
    .X(net5254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4731 (.A(net937),
    .X(net5255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4732 (.A(_00820_),
    .X(net5256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4733 (.A(net938),
    .X(net5257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4734 (.A(\rbzero.spi_registers.texadd1[11] ),
    .X(net5258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4735 (.A(net900),
    .X(net5259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4736 (.A(_00741_),
    .X(net5260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4737 (.A(net901),
    .X(net5261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4738 (.A(\rbzero.spi_registers.texadd3[0] ),
    .X(net5262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4739 (.A(net989),
    .X(net5263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(net5423),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4740 (.A(_00778_),
    .X(net5264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4741 (.A(net990),
    .X(net5265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4742 (.A(\rbzero.spi_registers.texadd1[2] ),
    .X(net5266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4743 (.A(net971),
    .X(net5267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4744 (.A(_00732_),
    .X(net5268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4745 (.A(net972),
    .X(net5269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4746 (.A(\rbzero.texV[-9] ),
    .X(net5270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4747 (.A(net880),
    .X(net5271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4748 (.A(_01591_),
    .X(net5272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4749 (.A(net881),
    .X(net5273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(net5425),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4750 (.A(\rbzero.spi_registers.texadd1[19] ),
    .X(net5274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4751 (.A(net943),
    .X(net5275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4752 (.A(_00749_),
    .X(net5276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4753 (.A(net944),
    .X(net5277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4754 (.A(\rbzero.spi_registers.buf_mapdyw[1] ),
    .X(net5278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4755 (.A(net973),
    .X(net5279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4756 (.A(_00852_),
    .X(net5280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4757 (.A(net974),
    .X(net5281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4758 (.A(\rbzero.spi_registers.buf_mapdxw[1] ),
    .X(net5282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4759 (.A(net865),
    .X(net5283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(net5405),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4760 (.A(_00850_),
    .X(net5284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4761 (.A(net866),
    .X(net5285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4762 (.A(\rbzero.spi_registers.texadd3[19] ),
    .X(net5286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4763 (.A(net1002),
    .X(net5287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4764 (.A(_00797_),
    .X(net5288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4765 (.A(net1003),
    .X(net5289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4766 (.A(\rbzero.spi_registers.texadd3[22] ),
    .X(net5290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4767 (.A(net983),
    .X(net5291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4768 (.A(_00800_),
    .X(net5292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4769 (.A(net984),
    .X(net5293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(net5407),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4770 (.A(\rbzero.spi_registers.texadd0[22] ),
    .X(net5294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4771 (.A(net919),
    .X(net5295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4772 (.A(_00728_),
    .X(net5296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4773 (.A(\rbzero.spi_registers.texadd1[0] ),
    .X(net5297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4774 (.A(net956),
    .X(net5298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4775 (.A(_00730_),
    .X(net5299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4776 (.A(net957),
    .X(net5300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4777 (.A(\rbzero.spi_registers.buf_vshift[4] ),
    .X(net5301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4778 (.A(net991),
    .X(net5302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4779 (.A(_00834_),
    .X(net5303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(net5286),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4780 (.A(net992),
    .X(net5304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4781 (.A(\rbzero.spi_registers.texadd1[1] ),
    .X(net5305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4782 (.A(net1038),
    .X(net5306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4783 (.A(_00731_),
    .X(net5307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4784 (.A(net1039),
    .X(net5308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4785 (.A(\rbzero.traced_texa[-5] ),
    .X(net5309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4786 (.A(net884),
    .X(net5310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4787 (.A(_00505_),
    .X(net5311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4788 (.A(net885),
    .X(net5312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4789 (.A(\rbzero.spi_registers.texadd1[17] ),
    .X(net5313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(net5288),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4790 (.A(net964),
    .X(net5314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4791 (.A(_00747_),
    .X(net5315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4792 (.A(net965),
    .X(net5316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4793 (.A(\rbzero.spi_registers.buf_texadd0[5] ),
    .X(net5317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4794 (.A(net939),
    .X(net5318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4795 (.A(_00858_),
    .X(net5319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4796 (.A(net940),
    .X(net5320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4797 (.A(\rbzero.spi_registers.buf_mapdxw[0] ),
    .X(net5321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4798 (.A(net904),
    .X(net5322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4799 (.A(_00849_),
    .X(net5323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(net5352),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4800 (.A(net905),
    .X(net5324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4801 (.A(\rbzero.color_floor[2] ),
    .X(net5325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4802 (.A(net1027),
    .X(net5326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4803 (.A(_00696_),
    .X(net5327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4804 (.A(net1028),
    .X(net5328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4805 (.A(\rbzero.color_floor[0] ),
    .X(net5329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4806 (.A(net915),
    .X(net5330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4807 (.A(_00694_),
    .X(net5331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4808 (.A(net916),
    .X(net5332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4809 (.A(\rbzero.texV[-8] ),
    .X(net5333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(net5354),
    .X(net1005));
 sky130_fd_sc_hd__buf_1 hold4810 (.A(net872),
    .X(net5334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4811 (.A(_01592_),
    .X(net5335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4812 (.A(net873),
    .X(net5336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4813 (.A(\rbzero.spi_registers.texadd3[4] ),
    .X(net5337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4814 (.A(net1025),
    .X(net5338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4815 (.A(_00782_),
    .X(net5339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4816 (.A(net1026),
    .X(net5340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4817 (.A(\rbzero.spi_registers.texadd1[4] ),
    .X(net5341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4818 (.A(net966),
    .X(net5342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4819 (.A(_00734_),
    .X(net5343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(net5427),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4820 (.A(net967),
    .X(net5344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4821 (.A(\rbzero.spi_registers.texadd3[5] ),
    .X(net5345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4822 (.A(net975),
    .X(net5346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4823 (.A(_00783_),
    .X(net5347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4824 (.A(net976),
    .X(net5348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4825 (.A(\rbzero.spi_registers.buf_texadd0[14] ),
    .X(net5349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4826 (.A(net606),
    .X(net5350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4827 (.A(_00867_),
    .X(net5351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4828 (.A(\rbzero.spi_registers.texadd0[8] ),
    .X(net5352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4829 (.A(net1004),
    .X(net5353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(net5429),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4830 (.A(_00714_),
    .X(net5354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4831 (.A(\rbzero.color_sky[5] ),
    .X(net5355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4832 (.A(net947),
    .X(net5356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4833 (.A(_00693_),
    .X(net5357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4834 (.A(net948),
    .X(net5358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4835 (.A(\rbzero.spi_registers.buf_vshift[5] ),
    .X(net5359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4836 (.A(net962),
    .X(net5360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4837 (.A(_00835_),
    .X(net5361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4838 (.A(net963),
    .X(net5362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4839 (.A(\rbzero.spi_registers.texadd0[23] ),
    .X(net5363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(net5446),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4840 (.A(net1052),
    .X(net5364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4841 (.A(_00729_),
    .X(net5365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4842 (.A(\rbzero.spi_registers.buf_otherx[1] ),
    .X(net5366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4843 (.A(net981),
    .X(net5367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4844 (.A(_00821_),
    .X(net5368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4845 (.A(net982),
    .X(net5369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4846 (.A(\rbzero.spi_registers.buf_mapdy[1] ),
    .X(net5370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4847 (.A(net993),
    .X(net5371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4848 (.A(_00844_),
    .X(net5372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4849 (.A(net994),
    .X(net5373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net5448),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4850 (.A(\rbzero.spi_registers.buf_othery[4] ),
    .X(net5374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4851 (.A(net960),
    .X(net5375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4852 (.A(_00829_),
    .X(net5376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4853 (.A(net961),
    .X(net5377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4854 (.A(\rbzero.traced_texa[-7] ),
    .X(net5378));
 sky130_fd_sc_hd__buf_1 hold4855 (.A(net945),
    .X(net5379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4856 (.A(_00503_),
    .X(net5380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4857 (.A(net946),
    .X(net5381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4858 (.A(\rbzero.pov.spi_buffer[42] ),
    .X(net5382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4859 (.A(net1284),
    .X(net5383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(net7498),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4860 (.A(_01078_),
    .X(net5384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4861 (.A(net1285),
    .X(net5385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4862 (.A(\rbzero.pov.spi_buffer[41] ),
    .X(net5386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4863 (.A(net1318),
    .X(net5387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4864 (.A(_01077_),
    .X(net5388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4865 (.A(net1319),
    .X(net5389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4866 (.A(\rbzero.spi_registers.buf_texadd0[9] ),
    .X(net5390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4867 (.A(net1045),
    .X(net5391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4868 (.A(_00862_),
    .X(net5392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4869 (.A(net1046),
    .X(net5393));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold487 (.A(\rbzero.traced_texa[-9] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4870 (.A(\rbzero.spi_registers.texadd0[15] ),
    .X(net5394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4871 (.A(net1066),
    .X(net5395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4872 (.A(_00721_),
    .X(net5396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4873 (.A(\rbzero.spi_registers.texadd3[2] ),
    .X(net5397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4874 (.A(net1056),
    .X(net5398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4875 (.A(_00780_),
    .X(net5399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4876 (.A(net1057),
    .X(net5400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4877 (.A(\rbzero.spi_registers.buf_otherx[4] ),
    .X(net5401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4878 (.A(net1021),
    .X(net5402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4879 (.A(_00824_),
    .X(net5403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(net7520),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4880 (.A(net1022),
    .X(net5404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4881 (.A(\rbzero.spi_registers.buf_othery[1] ),
    .X(net5405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4882 (.A(net1000),
    .X(net5406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4883 (.A(_00826_),
    .X(net5407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4884 (.A(net1001),
    .X(net5408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4885 (.A(\rbzero.pov.spi_buffer[7] ),
    .X(net5409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4886 (.A(net1222),
    .X(net5410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4887 (.A(_01043_),
    .X(net5411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4888 (.A(\rbzero.spi_registers.texadd3[18] ),
    .X(net5412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4889 (.A(net1029),
    .X(net5413));
 sky130_fd_sc_hd__buf_1 hold489 (.A(\rbzero.pov.ready_buffer[67] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4890 (.A(_00796_),
    .X(net5414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4891 (.A(net1030),
    .X(net5415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4892 (.A(\rbzero.spi_registers.texadd0[16] ),
    .X(net5416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4893 (.A(net1050),
    .X(net5417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4894 (.A(_00722_),
    .X(net5418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4895 (.A(\rbzero.wall_tracer.mapX[10] ),
    .X(net5419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4896 (.A(net977),
    .X(net5420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4897 (.A(_00527_),
    .X(net5421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4898 (.A(net978),
    .X(net5422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4899 (.A(\rbzero.texV[-6] ),
    .X(net5423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_03501_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4900 (.A(net998),
    .X(net5424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4901 (.A(_01594_),
    .X(net5425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4902 (.A(net999),
    .X(net5426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4903 (.A(\rbzero.spi_registers.buf_vshift[1] ),
    .X(net5427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4904 (.A(net1006),
    .X(net5428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4905 (.A(_00831_),
    .X(net5429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4906 (.A(net1007),
    .X(net5430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4907 (.A(net5444),
    .X(net5431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4908 (.A(net1493),
    .X(net5432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4909 (.A(_01086_),
    .X(net5433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(net4220),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4910 (.A(\rbzero.spi_registers.texadd3[3] ),
    .X(net5434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4911 (.A(net1043),
    .X(net5435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4912 (.A(_00781_),
    .X(net5436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4913 (.A(net1044),
    .X(net5437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4914 (.A(\rbzero.pov.spi_buffer[40] ),
    .X(net5438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4915 (.A(net1491),
    .X(net5439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4916 (.A(_01076_),
    .X(net5440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4917 (.A(\rbzero.mapdyw[0] ),
    .X(net5441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4918 (.A(net1054),
    .X(net5442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4919 (.A(_00680_),
    .X(net5443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(net5454),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4920 (.A(\rbzero.pov.spi_buffer[49] ),
    .X(net5444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4921 (.A(_01085_),
    .X(net5445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4922 (.A(\rbzero.mapdxw[1] ),
    .X(net5446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4923 (.A(net1008),
    .X(net5447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4924 (.A(_00679_),
    .X(net5448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4925 (.A(\rbzero.pov.spi_buffer[48] ),
    .X(net5449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4926 (.A(_01084_),
    .X(net5450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4927 (.A(\rbzero.spi_registers.texadd0[18] ),
    .X(net5451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4928 (.A(net1086),
    .X(net5452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4929 (.A(_00724_),
    .X(net5453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(net5456),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4930 (.A(\rbzero.texV[-5] ),
    .X(net5454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4931 (.A(net1016),
    .X(net5455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4932 (.A(_01595_),
    .X(net5456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4933 (.A(net1017),
    .X(net5457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4934 (.A(\rbzero.spi_registers.buf_othery[0] ),
    .X(net5458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4935 (.A(net1058),
    .X(net5459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4936 (.A(_00825_),
    .X(net5460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4937 (.A(net1059),
    .X(net5461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4938 (.A(net8009),
    .X(net5462));
 sky130_fd_sc_hd__buf_1 hold4939 (.A(net2933),
    .X(net5463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\rbzero.pov.ready_buffer[52] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4940 (.A(_00957_),
    .X(net5464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4941 (.A(net2934),
    .X(net5465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4942 (.A(\rbzero.pov.ready ),
    .X(net5466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4943 (.A(net1070),
    .X(net5467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4944 (.A(_01174_),
    .X(net5468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4945 (.A(net1071),
    .X(net5469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4946 (.A(\rbzero.traced_texa[-6] ),
    .X(net5470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4947 (.A(net985),
    .X(net5471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4948 (.A(_00504_),
    .X(net5472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4949 (.A(net986),
    .X(net5473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_03552_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4950 (.A(\rbzero.pov.spi_buffer[8] ),
    .X(net5474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4951 (.A(_01044_),
    .X(net5475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4952 (.A(\rbzero.spi_registers.texadd1[3] ),
    .X(net5476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4953 (.A(net1078),
    .X(net5477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4954 (.A(_00733_),
    .X(net5478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4955 (.A(net1079),
    .X(net5479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4956 (.A(net5484),
    .X(net5480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4957 (.A(net1335),
    .X(net5481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4958 (.A(_03714_),
    .X(net5482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4959 (.A(_01063_),
    .X(net5483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net4289),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4960 (.A(\rbzero.pov.spi_buffer[26] ),
    .X(net5484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4961 (.A(_01062_),
    .X(net5485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4962 (.A(\rbzero.spi_registers.texadd2[21] ),
    .X(net5486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4963 (.A(net1096),
    .X(net5487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4964 (.A(_00775_),
    .X(net5488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4965 (.A(net1097),
    .X(net5489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4966 (.A(\rbzero.wall_tracer.mapY[9] ),
    .X(net5490));
 sky130_fd_sc_hd__buf_1 hold4967 (.A(net2907),
    .X(net5491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4968 (.A(_00389_),
    .X(net5492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4969 (.A(net2908),
    .X(net5493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(net5401),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4970 (.A(\rbzero.pov.spi_buffer[29] ),
    .X(net5494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4971 (.A(_01065_),
    .X(net5495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4972 (.A(\rbzero.mapdxw[0] ),
    .X(net5496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4973 (.A(net1068),
    .X(net5497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4974 (.A(_00678_),
    .X(net5498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4975 (.A(\rbzero.pov.spi_buffer[16] ),
    .X(net5499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4976 (.A(net1105),
    .X(net5500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4977 (.A(_01052_),
    .X(net5501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4978 (.A(net1106),
    .X(net5502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4979 (.A(\rbzero.spi_registers.texadd2[17] ),
    .X(net5503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net5403),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4980 (.A(net1164),
    .X(net5504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4981 (.A(_00771_),
    .X(net5505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4982 (.A(net1165),
    .X(net5506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4983 (.A(\rbzero.pov.spi_buffer[4] ),
    .X(net5507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4984 (.A(_01040_),
    .X(net5508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4985 (.A(\rbzero.wall_tracer.mapY[10] ),
    .X(net5509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4986 (.A(net1064),
    .X(net5510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4987 (.A(_00390_),
    .X(net5511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4988 (.A(\rbzero.floor_leak[0] ),
    .X(net5512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4989 (.A(net1113),
    .X(net5513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net4247),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4990 (.A(_00682_),
    .X(net5514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4991 (.A(net1114),
    .X(net5515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4992 (.A(\rbzero.pov.spi_buffer[22] ),
    .X(net5516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4993 (.A(net1288),
    .X(net5517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4994 (.A(_01058_),
    .X(net5518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4995 (.A(\rbzero.pov.spi_buffer[23] ),
    .X(net5519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4996 (.A(net1263),
    .X(net5520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4997 (.A(_01059_),
    .X(net5521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4998 (.A(\rbzero.spi_registers.texadd2[20] ),
    .X(net5522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4999 (.A(net1118),
    .X(net5523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net4249),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5000 (.A(_00774_),
    .X(net5524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5001 (.A(net1119),
    .X(net5525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5002 (.A(\rbzero.spi_registers.texadd2[18] ),
    .X(net5526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5003 (.A(net1151),
    .X(net5527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5004 (.A(_00772_),
    .X(net5528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5005 (.A(net1152),
    .X(net5529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5006 (.A(\rbzero.pov.spi_buffer[10] ),
    .X(net5530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5007 (.A(_01046_),
    .X(net5531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5008 (.A(\rbzero.pov.spi_buffer[34] ),
    .X(net5532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5009 (.A(net1510),
    .X(net5533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(net5337),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5010 (.A(_01070_),
    .X(net5534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5011 (.A(\rbzero.spi_registers.texadd3[6] ),
    .X(net5535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5012 (.A(net1194),
    .X(net5536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5013 (.A(_00784_),
    .X(net5537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5014 (.A(net1195),
    .X(net5538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5015 (.A(\rbzero.pov.spi_buffer[18] ),
    .X(net5539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5016 (.A(net1294),
    .X(net5540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5017 (.A(_01054_),
    .X(net5541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5018 (.A(net1295),
    .X(net5542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5019 (.A(\rbzero.pov.spi_buffer[24] ),
    .X(net5543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(net5339),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5020 (.A(net1292),
    .X(net5544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5021 (.A(_01060_),
    .X(net5545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5022 (.A(\rbzero.spi_registers.buf_vshift[2] ),
    .X(net5546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5023 (.A(net1146),
    .X(net5547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5024 (.A(_00832_),
    .X(net5548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5025 (.A(net1147),
    .X(net5549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5026 (.A(\rbzero.pov.spi_buffer[5] ),
    .X(net5550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5027 (.A(net1204),
    .X(net5551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5028 (.A(_01041_),
    .X(net5552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5029 (.A(\rbzero.pov.spi_buffer[11] ),
    .X(net5553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(net5325),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5030 (.A(net1286),
    .X(net5554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5031 (.A(_01047_),
    .X(net5555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5032 (.A(\rbzero.pov.spi_buffer[3] ),
    .X(net5556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5033 (.A(_01039_),
    .X(net5557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5034 (.A(\rbzero.map_overlay.i_mapdx[5] ),
    .X(net5558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5035 (.A(net1185),
    .X(net5559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5036 (.A(_00671_),
    .X(net5560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5037 (.A(\rbzero.spi_registers.buf_otherx[2] ),
    .X(net5561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5038 (.A(net1123),
    .X(net5562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5039 (.A(_00822_),
    .X(net5563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(net5327),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5040 (.A(net1124),
    .X(net5564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5041 (.A(\rbzero.pov.spi_buffer[14] ),
    .X(net5565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5042 (.A(net1168),
    .X(net5566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5043 (.A(_01050_),
    .X(net5567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5044 (.A(\rbzero.pov.spi_buffer[25] ),
    .X(net5568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5045 (.A(_01061_),
    .X(net5569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5046 (.A(\rbzero.pov.spi_buffer[0] ),
    .X(net5570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5047 (.A(net3268),
    .X(net5571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5048 (.A(_03681_),
    .X(net5572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5049 (.A(_01037_),
    .X(net5573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net5412),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5050 (.A(\rbzero.pov.spi_buffer[19] ),
    .X(net5574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5051 (.A(net1389),
    .X(net5575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5052 (.A(_01055_),
    .X(net5576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5053 (.A(\rbzero.spi_registers.texadd3[13] ),
    .X(net5577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5054 (.A(net1261),
    .X(net5578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5055 (.A(_00791_),
    .X(net5579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5056 (.A(net1262),
    .X(net5580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5057 (.A(\rbzero.pov.spi_buffer[17] ),
    .X(net5581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5058 (.A(net1276),
    .X(net5582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5059 (.A(_01053_),
    .X(net5583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(net5414),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5060 (.A(\rbzero.pov.spi_buffer[15] ),
    .X(net5584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5061 (.A(net1162),
    .X(net5585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5062 (.A(_01051_),
    .X(net5586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5063 (.A(\rbzero.pov.spi_buffer[58] ),
    .X(net5587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5064 (.A(net1265),
    .X(net5588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5065 (.A(_01094_),
    .X(net5589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5066 (.A(\rbzero.pov.spi_buffer[20] ),
    .X(net5590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5067 (.A(net1280),
    .X(net5591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5068 (.A(_01056_),
    .X(net5592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5069 (.A(\rbzero.spi_registers.texadd2[1] ),
    .X(net5593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(net6350),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5070 (.A(net1308),
    .X(net5594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5071 (.A(_00755_),
    .X(net5595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5072 (.A(net1309),
    .X(net5596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5073 (.A(\rbzero.pov.mosi ),
    .X(net5597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5074 (.A(net953),
    .X(net5598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5075 (.A(_01036_),
    .X(net5599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5076 (.A(\rbzero.pov.spi_buffer[12] ),
    .X(net5600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5077 (.A(_01048_),
    .X(net5601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5078 (.A(\rbzero.pov.spi_buffer[21] ),
    .X(net5602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5079 (.A(_01057_),
    .X(net5603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(net6352),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5080 (.A(\rbzero.spi_registers.texadd3[7] ),
    .X(net5604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5081 (.A(net1255),
    .X(net5605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5082 (.A(_00785_),
    .X(net5606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5083 (.A(net1256),
    .X(net5607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5084 (.A(\rbzero.spi_registers.texadd0[4] ),
    .X(net5608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5085 (.A(net1310),
    .X(net5609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5086 (.A(_00710_),
    .X(net5610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5087 (.A(\rbzero.pov.spi_buffer[2] ),
    .X(net5611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5088 (.A(_01038_),
    .X(net5612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5089 (.A(\rbzero.spi_registers.texadd1[13] ),
    .X(net5613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_01129_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5090 (.A(net1377),
    .X(net5614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5091 (.A(_00743_),
    .X(net5615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5092 (.A(net1378),
    .X(net5616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5093 (.A(\rbzero.pov.spi_buffer[28] ),
    .X(net5617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5094 (.A(\rbzero.spi_registers.spi_counter[6] ),
    .X(net5618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5095 (.A(net1296),
    .X(net5619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5096 (.A(_00627_),
    .X(net5620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5097 (.A(net1297),
    .X(net5621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5098 (.A(\rbzero.pov.spi_buffer[53] ),
    .X(net5622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5099 (.A(net1337),
    .X(net5623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(net3309),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5100 (.A(_01089_),
    .X(net5624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5101 (.A(\rbzero.pov.spi_buffer[37] ),
    .X(net5625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5102 (.A(net1341),
    .X(net5626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5103 (.A(_01073_),
    .X(net5627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5104 (.A(\rbzero.spi_registers.texadd2[22] ),
    .X(net5628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5105 (.A(net1300),
    .X(net5629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5106 (.A(_00776_),
    .X(net5630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5107 (.A(net1301),
    .X(net5631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5108 (.A(\rbzero.spi_registers.texadd2[4] ),
    .X(net5632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5109 (.A(net1368),
    .X(net5633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_03522_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5110 (.A(_00758_),
    .X(net5634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5111 (.A(net1369),
    .X(net5635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5112 (.A(\rbzero.pov.spi_buffer[52] ),
    .X(net5636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5113 (.A(_01088_),
    .X(net5637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5114 (.A(\rbzero.spi_registers.texadd0[5] ),
    .X(net5638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5115 (.A(net1420),
    .X(net5639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5116 (.A(_00711_),
    .X(net5640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5117 (.A(\rbzero.spi_registers.texadd2[2] ),
    .X(net5641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5118 (.A(net1345),
    .X(net5642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5119 (.A(_00756_),
    .X(net5643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_03524_),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5120 (.A(net1346),
    .X(net5644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5121 (.A(\rbzero.pov.spi_buffer[38] ),
    .X(net5645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5122 (.A(net1475),
    .X(net5646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5123 (.A(_01074_),
    .X(net5647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5124 (.A(\rbzero.spi_registers.texadd0[9] ),
    .X(net5648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5125 (.A(net1320),
    .X(net5649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5126 (.A(_00715_),
    .X(net5650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5127 (.A(\rbzero.spi_registers.texadd2[3] ),
    .X(net5651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5128 (.A(net1330),
    .X(net5652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5129 (.A(_00757_),
    .X(net5653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_00968_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5130 (.A(net1331),
    .X(net5654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5131 (.A(\rbzero.floor_leak[3] ),
    .X(net5655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5132 (.A(net1326),
    .X(net5656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5133 (.A(_00685_),
    .X(net5657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5134 (.A(net1327),
    .X(net5658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5135 (.A(\rbzero.spi_registers.texadd1[21] ),
    .X(net5659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5136 (.A(net1391),
    .X(net5660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5137 (.A(_00751_),
    .X(net5661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5138 (.A(net1392),
    .X(net5662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5139 (.A(\rbzero.pov.spi_buffer[13] ),
    .X(net5663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(net5305),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5140 (.A(\rbzero.pov.spi_buffer[54] ),
    .X(net5664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5141 (.A(net1400),
    .X(net5665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5142 (.A(_01090_),
    .X(net5666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5143 (.A(\rbzero.pov.spi_buffer[39] ),
    .X(net5667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5144 (.A(\rbzero.spi_registers.texadd0[2] ),
    .X(net5668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5145 (.A(net1350),
    .X(net5669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5146 (.A(_00708_),
    .X(net5670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5147 (.A(\rbzero.pov.spi_buffer[36] ),
    .X(net5671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5148 (.A(_01072_),
    .X(net5672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5149 (.A(\rbzero.spi_registers.texadd2[5] ),
    .X(net5673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(net5307),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5150 (.A(net1404),
    .X(net5674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5151 (.A(_00759_),
    .X(net5675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5152 (.A(net1405),
    .X(net5676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5153 (.A(\rbzero.mapdyw[1] ),
    .X(net5677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5154 (.A(net1312),
    .X(net5678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5155 (.A(_00681_),
    .X(net5679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5156 (.A(\rbzero.spi_registers.texadd0[19] ),
    .X(net5680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5157 (.A(net1379),
    .X(net5681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5158 (.A(_00725_),
    .X(net5682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5159 (.A(net7833),
    .X(net5683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net6370),
    .X(net1040));
 sky130_fd_sc_hd__buf_1 hold5160 (.A(net3063),
    .X(net5684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5161 (.A(_08162_),
    .X(net5685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5162 (.A(_08169_),
    .X(net5686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5163 (.A(\rbzero.pov.spi_buffer[35] ),
    .X(net5687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5164 (.A(_01071_),
    .X(net5688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5165 (.A(\rbzero.spi_registers.texadd3[8] ),
    .X(net5689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5166 (.A(net1415),
    .X(net5690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5167 (.A(_00786_),
    .X(net5691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5168 (.A(net1416),
    .X(net5692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5169 (.A(\rbzero.pov.spi_buffer[51] ),
    .X(net5693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net6372),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5170 (.A(_01087_),
    .X(net5694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5171 (.A(\rbzero.pov.ready_buffer[21] ),
    .X(net5695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5172 (.A(net1440),
    .X(net5696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5173 (.A(_01017_),
    .X(net5697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5174 (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .X(net5698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5175 (.A(net3619),
    .X(net5699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5176 (.A(_00670_),
    .X(net5700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5177 (.A(\rbzero.floor_leak[4] ),
    .X(net5701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5178 (.A(net1402),
    .X(net5702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5179 (.A(_00686_),
    .X(net5703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_01572_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5180 (.A(net1403),
    .X(net5704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5181 (.A(\rbzero.wall_tracer.mapY[7] ),
    .X(net5705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5182 (.A(net2768),
    .X(net5706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5183 (.A(_00387_),
    .X(net5707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5184 (.A(net2769),
    .X(net5708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5185 (.A(\rbzero.floor_leak[2] ),
    .X(net5709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5186 (.A(net1524),
    .X(net5710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5187 (.A(_00684_),
    .X(net5711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5188 (.A(net1525),
    .X(net5712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5189 (.A(\rbzero.spi_registers.texadd1[22] ),
    .X(net5713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net5434),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5190 (.A(net1585),
    .X(net5714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5191 (.A(_00752_),
    .X(net5715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5192 (.A(net1586),
    .X(net5716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5193 (.A(\rbzero.spi_registers.buf_texadd2[15] ),
    .X(net5717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5194 (.A(net1214),
    .X(net5718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5195 (.A(_03415_),
    .X(net5719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5196 (.A(\rbzero.spi_registers.vshift[1] ),
    .X(net5720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5197 (.A(net1529),
    .X(net5721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5198 (.A(_00701_),
    .X(net5722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5199 (.A(\rbzero.spi_registers.texadd1[23] ),
    .X(net5723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net5436),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5200 (.A(net1557),
    .X(net5724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5201 (.A(_00753_),
    .X(net5725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5202 (.A(net1558),
    .X(net5726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5203 (.A(\rbzero.spi_registers.buf_texadd2[0] ),
    .X(net5727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5204 (.A(net1083),
    .X(net5728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5205 (.A(_03396_),
    .X(net5729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5206 (.A(_00901_),
    .X(net5730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5207 (.A(net1573),
    .X(net5731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5208 (.A(\rbzero.map_overlay.i_mapdy[5] ),
    .X(net5732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5209 (.A(net1506),
    .X(net5733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(net5390),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5210 (.A(_00677_),
    .X(net5734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5211 (.A(\rbzero.spi_registers.texadd2[7] ),
    .X(net5735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5212 (.A(net1589),
    .X(net5736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5213 (.A(_00761_),
    .X(net5737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5214 (.A(net1590),
    .X(net5738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5215 (.A(\rbzero.spi_registers.texadd0[0] ),
    .X(net5739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5216 (.A(net1827),
    .X(net5740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5217 (.A(_00706_),
    .X(net5741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5218 (.A(\rbzero.spi_registers.texadd0[3] ),
    .X(net5742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5219 (.A(net1593),
    .X(net5743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net5392),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5220 (.A(_00709_),
    .X(net5744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5221 (.A(\rbzero.wall_tracer.mapX[9] ),
    .X(net5745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5222 (.A(net2787),
    .X(net5746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5223 (.A(_00526_),
    .X(net5747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5224 (.A(net2788),
    .X(net5748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5225 (.A(\rbzero.spi_registers.texadd2[9] ),
    .X(net5749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5226 (.A(net1618),
    .X(net5750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5227 (.A(_00763_),
    .X(net5751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5228 (.A(net1619),
    .X(net5752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5229 (.A(\rbzero.spi_registers.buf_leak[1] ),
    .X(net5753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(net6340),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5230 (.A(net1141),
    .X(net5754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5231 (.A(_03268_),
    .X(net5755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5232 (.A(_00815_),
    .X(net5756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5233 (.A(\rbzero.spi_registers.texadd2[8] ),
    .X(net5757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5234 (.A(net1695),
    .X(net5758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5235 (.A(_00762_),
    .X(net5759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5236 (.A(net1696),
    .X(net5760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5237 (.A(\rbzero.spi_registers.buf_texadd2[23] ),
    .X(net5761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5238 (.A(net1115),
    .X(net5762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5239 (.A(_03423_),
    .X(net5763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_04158_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5240 (.A(_00924_),
    .X(net5764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5241 (.A(net1614),
    .X(net5765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5242 (.A(\rbzero.pov.spi_buffer[55] ),
    .X(net5766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5243 (.A(\rbzero.tex_b0[1] ),
    .X(net5767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5244 (.A(_04596_),
    .X(net5768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5245 (.A(net1522),
    .X(net5769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5246 (.A(\rbzero.pov.spi_buffer[59] ),
    .X(net5770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5247 (.A(_01095_),
    .X(net5771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5248 (.A(\rbzero.spi_registers.vshift[0] ),
    .X(net5772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5249 (.A(net1650),
    .X(net5773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_01651_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5250 (.A(_00700_),
    .X(net5774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5251 (.A(\rbzero.tex_r0[1] ),
    .X(net5775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5252 (.A(_04314_),
    .X(net5776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5253 (.A(net1489),
    .X(net5777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5254 (.A(\rbzero.pov.spi_buffer[56] ),
    .X(net5778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5255 (.A(\rbzero.spi_registers.vshift[2] ),
    .X(net5779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5256 (.A(net1569),
    .X(net5780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5257 (.A(_00702_),
    .X(net5781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5258 (.A(\rbzero.spi_registers.buf_leak[5] ),
    .X(net5782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5259 (.A(net1634),
    .X(net5783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net5416),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5260 (.A(_03272_),
    .X(net5784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5261 (.A(_00819_),
    .X(net5785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5262 (.A(net1728),
    .X(net5786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5263 (.A(\rbzero.spi_registers.texadd0[1] ),
    .X(net5787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5264 (.A(net1721),
    .X(net5788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5265 (.A(_00707_),
    .X(net5789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5266 (.A(\rbzero.pov.spi_buffer[57] ),
    .X(net5790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5267 (.A(\rbzero.spi_registers.buf_texadd2[6] ),
    .X(net5791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5268 (.A(net1217),
    .X(net5792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5269 (.A(_03403_),
    .X(net5793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(net5418),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5270 (.A(\rbzero.spi_registers.buf_texadd2[12] ),
    .X(net5794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5271 (.A(net1655),
    .X(net5795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5272 (.A(_03411_),
    .X(net5796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5273 (.A(_00913_),
    .X(net5797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5274 (.A(\rbzero.tex_r1[38] ),
    .X(net5798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5275 (.A(_04198_),
    .X(net5799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5276 (.A(net1763),
    .X(net5800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5277 (.A(\rbzero.spi_registers.vshift[5] ),
    .X(net5801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5278 (.A(net1915),
    .X(net5802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5279 (.A(_00705_),
    .X(net5803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net5363),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5280 (.A(net5941),
    .X(net5804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5281 (.A(_04247_),
    .X(net5805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5282 (.A(net1933),
    .X(net5806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5283 (.A(\rbzero.map_overlay.i_otherx[3] ),
    .X(net5807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5284 (.A(net2043),
    .X(net5808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5285 (.A(_00658_),
    .X(net5809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5286 (.A(\rbzero.tex_r1[37] ),
    .X(net5810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5287 (.A(net1992),
    .X(net5811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5288 (.A(_04199_),
    .X(net5812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5289 (.A(net1993),
    .X(net5813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net5365),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5290 (.A(\rbzero.tex_b1[60] ),
    .X(net5814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5291 (.A(_04462_),
    .X(net5815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5292 (.A(net2141),
    .X(net5816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5293 (.A(\rbzero.tex_b0[58] ),
    .X(net5817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5294 (.A(_04534_),
    .X(net5818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5295 (.A(net1968),
    .X(net5819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5296 (.A(\rbzero.tex_r1[40] ),
    .X(net5820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5297 (.A(net588),
    .X(net5821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5298 (.A(_04197_),
    .X(net5822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5299 (.A(net589),
    .X(net5823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(net5441),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5300 (.A(\rbzero.tex_r1[58] ),
    .X(net5824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5301 (.A(_04176_),
    .X(net5825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5302 (.A(net2428),
    .X(net5826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5303 (.A(\rbzero.tex_r1[57] ),
    .X(net5827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5304 (.A(net2472),
    .X(net5828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5305 (.A(_04177_),
    .X(net5829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5306 (.A(net2473),
    .X(net5830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5307 (.A(\rbzero.tex_g1[2] ),
    .X(net5831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5308 (.A(_04384_),
    .X(net5832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5309 (.A(net2443),
    .X(net5833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net5443),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5310 (.A(\rbzero.tex_g0[34] ),
    .X(net5834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5311 (.A(_04420_),
    .X(net5835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5312 (.A(net1957),
    .X(net5836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5313 (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .X(net5837));
 sky130_fd_sc_hd__clkbuf_2 hold5314 (.A(net614),
    .X(net5838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5315 (.A(_00935_),
    .X(net5839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5316 (.A(net649),
    .X(net5840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5317 (.A(\rbzero.tex_b1[2] ),
    .X(net5841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5318 (.A(_04525_),
    .X(net5842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5319 (.A(net2038),
    .X(net5843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(net5397),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5320 (.A(\rbzero.tex_g1[46] ),
    .X(net5844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5321 (.A(_04336_),
    .X(net5845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5322 (.A(net2397),
    .X(net5846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5323 (.A(\rbzero.tex_b1[61] ),
    .X(net5847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5324 (.A(net1832),
    .X(net5848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5325 (.A(_04461_),
    .X(net5849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5326 (.A(net1833),
    .X(net5850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5327 (.A(\rbzero.spi_registers.vshift[3] ),
    .X(net5851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5328 (.A(net2194),
    .X(net5852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5329 (.A(_00703_),
    .X(net5853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(net5399),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5330 (.A(\rbzero.tex_g1[32] ),
    .X(net5854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5331 (.A(_04351_),
    .X(net5855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5332 (.A(net2002),
    .X(net5856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5333 (.A(\rbzero.tex_r1[4] ),
    .X(net5857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5334 (.A(_04235_),
    .X(net5858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5335 (.A(net1459),
    .X(net5859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5336 (.A(\rbzero.spi_registers.buf_texadd3[14] ),
    .X(net5860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5337 (.A(net2155),
    .X(net5861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5338 (.A(_03227_),
    .X(net5862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5339 (.A(_00792_),
    .X(net5863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net5458),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5340 (.A(net2353),
    .X(net5864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5341 (.A(\rbzero.tex_b1[28] ),
    .X(net5865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5342 (.A(_04497_),
    .X(net5866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5343 (.A(net2120),
    .X(net5867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5344 (.A(\rbzero.tex_b1[42] ),
    .X(net5868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5345 (.A(_04482_),
    .X(net5869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5346 (.A(net1857),
    .X(net5870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5347 (.A(\rbzero.tex_b1[29] ),
    .X(net5871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5348 (.A(net2464),
    .X(net5872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5349 (.A(_04496_),
    .X(net5873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(net5460),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5350 (.A(net2465),
    .X(net5874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5351 (.A(\rbzero.map_overlay.i_othery[3] ),
    .X(net5875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5352 (.A(net2536),
    .X(net5876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5353 (.A(_00663_),
    .X(net5877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5354 (.A(\rbzero.tex_g1[3] ),
    .X(net5878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5355 (.A(net2097),
    .X(net5879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5356 (.A(_04383_),
    .X(net5880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5357 (.A(net2098),
    .X(net5881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5358 (.A(\rbzero.spi_registers.vshift[4] ),
    .X(net5882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5359 (.A(net2467),
    .X(net5883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(net7449),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5360 (.A(_00704_),
    .X(net5884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5361 (.A(\rbzero.tex_r1[3] ),
    .X(net5885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5362 (.A(net2393),
    .X(net5886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5363 (.A(_04237_),
    .X(net5887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5364 (.A(net2394),
    .X(net5888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5365 (.A(\rbzero.tex_b1[3] ),
    .X(net5889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5366 (.A(net1874),
    .X(net5890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5367 (.A(_04524_),
    .X(net5891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5368 (.A(net1875),
    .X(net5892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5369 (.A(\rbzero.tex_g1[52] ),
    .X(net5893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net6366),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5370 (.A(_04328_),
    .X(net5894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5371 (.A(net2633),
    .X(net5895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5372 (.A(\rbzero.tex_g1[33] ),
    .X(net5896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5373 (.A(net1780),
    .X(net5897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5374 (.A(_04350_),
    .X(net5898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5375 (.A(net1781),
    .X(net5899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5376 (.A(\rbzero.tex_b1[24] ),
    .X(net5900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5377 (.A(_04501_),
    .X(net5901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5378 (.A(net2180),
    .X(net5902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5379 (.A(\rbzero.tex_b1[43] ),
    .X(net5903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(net6368),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5380 (.A(net2176),
    .X(net5904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5381 (.A(_04480_),
    .X(net5905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5382 (.A(net2177),
    .X(net5906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5383 (.A(\rbzero.map_overlay.i_otherx[0] ),
    .X(net5907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5384 (.A(net2677),
    .X(net5908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5385 (.A(_00655_),
    .X(net5909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5386 (.A(\rbzero.tex_r0[2] ),
    .X(net5910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5387 (.A(net2562),
    .X(net5911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5388 (.A(_04313_),
    .X(net5912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5389 (.A(net2563),
    .X(net5913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_01432_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5390 (.A(\rbzero.tex_r1[28] ),
    .X(net5914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5391 (.A(_04210_),
    .X(net5915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5392 (.A(net2557),
    .X(net5916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5393 (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .X(net5917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5394 (.A(net2802),
    .X(net5918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5395 (.A(_00672_),
    .X(net5919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5396 (.A(\rbzero.tex_g0[1] ),
    .X(net5920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5397 (.A(_04455_),
    .X(net5921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5398 (.A(net751),
    .X(net5922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5399 (.A(\rbzero.tex_b0[2] ),
    .X(net5923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(net5509),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5400 (.A(net2650),
    .X(net5924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5401 (.A(_04595_),
    .X(net5925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5402 (.A(net2651),
    .X(net5926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5403 (.A(net5975),
    .X(net5927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5404 (.A(_04227_),
    .X(net5928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5405 (.A(net1684),
    .X(net5929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5406 (.A(\rbzero.tex_g1[47] ),
    .X(net5930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5407 (.A(net1941),
    .X(net5931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5408 (.A(_04335_),
    .X(net5932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5409 (.A(net1942),
    .X(net5933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(net5511),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5410 (.A(\rbzero.tex_g0[0] ),
    .X(net5934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5411 (.A(net2191),
    .X(net5935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5412 (.A(_04456_),
    .X(net5936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5413 (.A(net2192),
    .X(net5937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5414 (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .X(net5938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5415 (.A(net2726),
    .X(net5939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5416 (.A(_00676_),
    .X(net5940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5417 (.A(\rbzero.tex_r0[62] ),
    .X(net5941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5418 (.A(net5804),
    .X(net5942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5419 (.A(\rbzero.map_overlay.i_otherx[1] ),
    .X(net5943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(net5394),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5420 (.A(net2705),
    .X(net5944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5421 (.A(_00656_),
    .X(net5945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5422 (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .X(net5946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5423 (.A(net2791),
    .X(net5947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5424 (.A(_00675_),
    .X(net5948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5425 (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .X(net5949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5426 (.A(net2825),
    .X(net5950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5427 (.A(_00668_),
    .X(net5951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5428 (.A(\rbzero.tex_b0[59] ),
    .X(net5952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5429 (.A(net1970),
    .X(net5953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(net5396),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5430 (.A(_04533_),
    .X(net5954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5431 (.A(net1971),
    .X(net5955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5432 (.A(\gpout0.vpos[7] ),
    .X(net5956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5433 (.A(net4001),
    .X(net5957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5434 (.A(\rbzero.map_overlay.i_othery[2] ),
    .X(net5958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5435 (.A(net2864),
    .X(net5959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5436 (.A(_00662_),
    .X(net5960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5437 (.A(\rbzero.tex_b1[25] ),
    .X(net5961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5438 (.A(net2182),
    .X(net5962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5439 (.A(_04500_),
    .X(net5963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(net5496),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5440 (.A(net2183),
    .X(net5964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5441 (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .X(net5965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5442 (.A(net2774),
    .X(net5966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5443 (.A(_00666_),
    .X(net5967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5444 (.A(\rbzero.wall_tracer.mapX[7] ),
    .X(net5968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5445 (.A(net2611),
    .X(net5969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5446 (.A(_00524_),
    .X(net5970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5447 (.A(net2612),
    .X(net5971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5448 (.A(\rbzero.map_overlay.i_otherx[4] ),
    .X(net5972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5449 (.A(net2839),
    .X(net5973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(net5498),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5450 (.A(_00659_),
    .X(net5974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5451 (.A(\rbzero.tex_r1[12] ),
    .X(net5975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5452 (.A(net5927),
    .X(net5976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5453 (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .X(net5977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5454 (.A(net2789),
    .X(net5978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5455 (.A(_00674_),
    .X(net5979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5456 (.A(\rbzero.tex_r1[29] ),
    .X(net5980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5457 (.A(net2493),
    .X(net5981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5458 (.A(_04209_),
    .X(net5982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5459 (.A(net2494),
    .X(net5983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(net5466),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5460 (.A(\rbzero.tex_g0[35] ),
    .X(net5984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5461 (.A(net1938),
    .X(net5985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5462 (.A(_04419_),
    .X(net5986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5463 (.A(net1939),
    .X(net5987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5464 (.A(\rbzero.tex_g1[53] ),
    .X(net5988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5465 (.A(net1554),
    .X(net5989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5466 (.A(_04327_),
    .X(net5990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5467 (.A(net1555),
    .X(net5991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5468 (.A(\rbzero.map_overlay.i_othery[4] ),
    .X(net5992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5469 (.A(net2823),
    .X(net5993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(net5468),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5470 (.A(_00664_),
    .X(net5994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5471 (.A(\rbzero.floor_leak[5] ),
    .X(net5995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5472 (.A(net4076),
    .X(net5996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5473 (.A(_00687_),
    .X(net5997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5474 (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .X(net5998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5475 (.A(net2895),
    .X(net5999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5476 (.A(_00667_),
    .X(net6000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5477 (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .X(net6001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5478 (.A(net2879),
    .X(net6002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5479 (.A(_00673_),
    .X(net6003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(net7712),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5480 (.A(\rbzero.map_overlay.i_othery[1] ),
    .X(net6004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5481 (.A(net2905),
    .X(net6005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5482 (.A(_00661_),
    .X(net6006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5483 (.A(\rbzero.pov.ready_buffer[63] ),
    .X(net6007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5484 (.A(net3732),
    .X(net6008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5485 (.A(_03492_),
    .X(net6009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5486 (.A(_03493_),
    .X(net6010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5487 (.A(_00959_),
    .X(net6011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5488 (.A(net2936),
    .X(net6012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5489 (.A(\rbzero.map_overlay.i_otherx[2] ),
    .X(net6013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(net6390),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5490 (.A(net2917),
    .X(net6014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5491 (.A(_00657_),
    .X(net6015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5492 (.A(\rbzero.map_overlay.i_othery[0] ),
    .X(net6016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5493 (.A(net2925),
    .X(net6017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5494 (.A(_00660_),
    .X(net6018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5495 (.A(\rbzero.pov.ready_buffer[10] ),
    .X(net6019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5496 (.A(net2900),
    .X(net6020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5497 (.A(_01028_),
    .X(net6021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5498 (.A(\rbzero.row_render.size[4] ),
    .X(net6022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5499 (.A(net2993),
    .X(net6023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net6392),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5500 (.A(\gpout0.hpos[3] ),
    .X(net6024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5501 (.A(net3908),
    .X(net6025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5502 (.A(_01253_),
    .X(net6026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5503 (.A(net2989),
    .X(net6027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5504 (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .X(net6028));
 sky130_fd_sc_hd__clkbuf_2 hold5505 (.A(net3072),
    .X(net6029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5506 (.A(_00894_),
    .X(net6030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5507 (.A(net1861),
    .X(net6031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5508 (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .X(net6032));
 sky130_fd_sc_hd__buf_1 hold5509 (.A(net1613),
    .X(net6033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_01342_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5510 (.A(_00948_),
    .X(net6034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5511 (.A(net2875),
    .X(net6035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5512 (.A(\rbzero.spi_registers.buf_texadd3[21] ),
    .X(net6036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5513 (.A(net2230),
    .X(net6037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5514 (.A(_03456_),
    .X(net6038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5515 (.A(_00946_),
    .X(net6039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5516 (.A(\gpout0.vpos[8] ),
    .X(net6040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5517 (.A(net3929),
    .X(net6041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5518 (.A(\rbzero.spi_registers.buf_texadd1[23] ),
    .X(net6042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5519 (.A(net1548),
    .X(net6043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(net7639),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5520 (.A(_03390_),
    .X(net6044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5521 (.A(_00900_),
    .X(net6045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5522 (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .X(net6046));
 sky130_fd_sc_hd__clkbuf_2 hold5523 (.A(net2948),
    .X(net6047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5524 (.A(\gpout0.hpos[2] ),
    .X(net6048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5525 (.A(net3987),
    .X(net6049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5526 (.A(\rbzero.spi_registers.buf_texadd3[22] ),
    .X(net6050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5527 (.A(net2282),
    .X(net6051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5528 (.A(_03457_),
    .X(net6052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5529 (.A(_00947_),
    .X(net6053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(net4480),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5530 (.A(\rbzero.spi_registers.buf_texadd2[21] ),
    .X(net6054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5531 (.A(net1574),
    .X(net6055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5532 (.A(_03421_),
    .X(net6056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5533 (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .X(net6057));
 sky130_fd_sc_hd__clkbuf_2 hold5534 (.A(net1591),
    .X(net6058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5535 (.A(\rbzero.spi_registers.buf_texadd3[17] ),
    .X(net6059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5536 (.A(net1844),
    .X(net6060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5537 (.A(\rbzero.spi_registers.buf_texadd1[21] ),
    .X(net6061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5538 (.A(net1712),
    .X(net6062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5539 (.A(_03388_),
    .X(net6063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(net5476),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5540 (.A(_00898_),
    .X(net6064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5541 (.A(\rbzero.spi_registers.buf_texadd2[17] ),
    .X(net6065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5542 (.A(net1644),
    .X(net6066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5544 (.A(_02842_),
    .X(net6068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5545 (.A(net3164),
    .X(net6069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5546 (.A(\rbzero.spi_registers.buf_texadd1[22] ),
    .X(net6070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5547 (.A(net1670),
    .X(net6071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5548 (.A(_03389_),
    .X(net6072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5549 (.A(_00899_),
    .X(net6073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(net5478),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5550 (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .X(net6074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5551 (.A(\rbzero.spi_registers.buf_texadd2[22] ),
    .X(net6075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5552 (.A(net2354),
    .X(net6076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5553 (.A(_03422_),
    .X(net6077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5555 (.A(_02568_),
    .X(net6079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5556 (.A(net3204),
    .X(net6080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5557 (.A(\rbzero.debug_overlay.playerY[-8] ),
    .X(net6081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5558 (.A(net3024),
    .X(net6082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5559 (.A(_00971_),
    .X(net6083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(net6346),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5561 (.A(_02578_),
    .X(net6085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5562 (.A(net3238),
    .X(net6086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5564 (.A(_02786_),
    .X(net6088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5565 (.A(net3247),
    .X(net6089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5567 (.A(_08204_),
    .X(net6091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5568 (.A(net3334),
    .X(net6092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_04013_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5570 (.A(_02659_),
    .X(net6094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5571 (.A(net3371),
    .X(net6095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5572 (.A(\rbzero.debug_overlay.playerY[-6] ),
    .X(net6096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5573 (.A(net2942),
    .X(net6097));
 sky130_fd_sc_hd__clkbuf_4 hold5574 (.A(net3222),
    .X(net6098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5575 (.A(_08232_),
    .X(net6099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5577 (.A(_02876_),
    .X(net6101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5578 (.A(net3409),
    .X(net6102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5579 (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .X(net6103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_01588_),
    .X(net1082));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5580 (.A(net642),
    .X(net6104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5581 (.A(_00896_),
    .X(net6105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5582 (.A(net1770),
    .X(net6106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5584 (.A(_02796_),
    .X(net6108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5585 (.A(net3458),
    .X(net6109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5586 (.A(\rbzero.spi_registers.buf_texadd3[19] ),
    .X(net6110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5587 (.A(net1631),
    .X(net6111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5588 (.A(\rbzero.map_rom.i_row[4] ),
    .X(net6112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5589 (.A(\rbzero.spi_registers.buf_texadd3[16] ),
    .X(net6113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net5727),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5590 (.A(net1566),
    .X(net6114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5592 (.A(_02600_),
    .X(net6116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5593 (.A(net3595),
    .X(net6117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5595 (.A(_02817_),
    .X(net6119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5596 (.A(net3726),
    .X(net6120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5598 (.A(_08197_),
    .X(net6122));
 sky130_fd_sc_hd__clkbuf_4 hold5599 (.A(net4524),
    .X(net6123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_03177_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5601 (.A(_08210_),
    .X(net6125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5602 (.A(\rbzero.debug_overlay.playerY[-4] ),
    .X(net6126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5603 (.A(net3003),
    .X(net6127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5604 (.A(_00975_),
    .X(net6128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5605 (.A(\rbzero.debug_overlay.playerX[-3] ),
    .X(net6129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5606 (.A(net3008),
    .X(net6130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5607 (.A(_00961_),
    .X(net6131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5609 (.A(_08193_),
    .X(net6133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(net4192),
    .X(net1085));
 sky130_fd_sc_hd__buf_1 hold5610 (.A(net3633),
    .X(net6134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5611 (.A(_08241_),
    .X(net6135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5612 (.A(net3634),
    .X(net6136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5614 (.A(_08202_),
    .X(net6138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5615 (.A(net3791),
    .X(net6139));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5616 (.A(\rbzero.debug_overlay.playerX[5] ),
    .X(net6140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5617 (.A(_02964_),
    .X(net6141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5618 (.A(_02965_),
    .X(net6142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(net5451),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5620 (.A(_08208_),
    .X(net6144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5621 (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .X(net6145));
 sky130_fd_sc_hd__clkbuf_4 hold5622 (.A(net3772),
    .X(net6146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5623 (.A(_08238_),
    .X(net6147));
 sky130_fd_sc_hd__clkbuf_4 hold5624 (.A(net3627),
    .X(net6148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5625 (.A(_08234_),
    .X(net6149));
 sky130_fd_sc_hd__clkbuf_4 hold5626 (.A(net3718),
    .X(net6150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5627 (.A(_08236_),
    .X(net6151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5629 (.A(_08206_),
    .X(net6153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(net5453),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5630 (.A(\rbzero.debug_overlay.playerX[0] ),
    .X(net6154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5631 (.A(net3821),
    .X(net6155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5632 (.A(_00964_),
    .X(net6156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5633 (.A(net746),
    .X(net6157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5634 (.A(\rbzero.map_rom.i_col[4] ),
    .X(net6158));
 sky130_fd_sc_hd__clkbuf_4 hold5638 (.A(net7886),
    .X(net6162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5639 (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .X(net6163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(net6374),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_2 hold5640 (.A(net3050),
    .X(net6164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5641 (.A(_00932_),
    .X(net6165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5642 (.A(net2072),
    .X(net6166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5643 (.A(\rbzero.trace_state[2] ),
    .X(net6167));
 sky130_fd_sc_hd__clkbuf_2 hold5644 (.A(net2982),
    .X(net6168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5645 (.A(\rbzero.spi_registers.buf_texadd1[7] ),
    .X(net6169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5646 (.A(net2090),
    .X(net6170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5647 (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .X(net6171));
 sky130_fd_sc_hd__buf_2 hold5648 (.A(net3093),
    .X(net6172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5649 (.A(_00933_),
    .X(net6173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(net6376),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5650 (.A(net1691),
    .X(net6174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5651 (.A(\rbzero.pov.spi_done ),
    .X(net6175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5652 (.A(net3249),
    .X(net6176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5653 (.A(_01249_),
    .X(net6177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5654 (.A(net2939),
    .X(net6178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5655 (.A(\rbzero.spi_registers.buf_texadd1[8] ),
    .X(net6179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5656 (.A(net2256),
    .X(net6180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5657 (.A(\rbzero.debug_overlay.playerX[2] ),
    .X(net6181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5658 (.A(net4090),
    .X(net6182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5659 (.A(_00966_),
    .X(net6183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_01282_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5660 (.A(net677),
    .X(net6184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5661 (.A(net6208),
    .X(net6185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5662 (.A(_06184_),
    .X(net6186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5663 (.A(_02735_),
    .X(net6187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5664 (.A(_02737_),
    .X(net6188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5665 (.A(_02738_),
    .X(net6189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5666 (.A(\rbzero.debug_overlay.playerY[-3] ),
    .X(net6190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5667 (.A(net4063),
    .X(net6191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5668 (.A(_00976_),
    .X(net6192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5669 (.A(net2958),
    .X(net6193));
 sky130_fd_sc_hd__buf_1 hold567 (.A(net7640),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5670 (.A(\rbzero.spi_registers.buf_texadd2[7] ),
    .X(net6194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5671 (.A(net2455),
    .X(net6195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5672 (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .X(net6196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5673 (.A(net3095),
    .X(net6197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5674 (.A(\rbzero.debug_overlay.playerX[-2] ),
    .X(net6198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5675 (.A(net3028),
    .X(net6199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5676 (.A(_00962_),
    .X(net6200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5677 (.A(\rbzero.spi_registers.buf_texadd2[8] ),
    .X(net6201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5678 (.A(net2533),
    .X(net6202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(net4553),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5680 (.A(_08212_),
    .X(net6204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5681 (.A(_00420_),
    .X(net6205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5682 (.A(\rbzero.debug_overlay.playerY[0] ),
    .X(net6206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5683 (.A(net3917),
    .X(net6207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5684 (.A(\rbzero.map_rom.c6 ),
    .X(net6208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5685 (.A(\rbzero.debug_overlay.playerX[3] ),
    .X(net6209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5686 (.A(net3921),
    .X(net6210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5687 (.A(_00967_),
    .X(net6211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5688 (.A(\rbzero.debug_overlay.playerY[3] ),
    .X(net6212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5689 (.A(net3893),
    .X(net6213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(net6378),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5690 (.A(_00982_),
    .X(net6214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5691 (.A(net749),
    .X(net6215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5692 (.A(\rbzero.map_rom.f1 ),
    .X(net6216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5693 (.A(_06222_),
    .X(net6217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5694 (.A(_02958_),
    .X(net6218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5695 (.A(\gpout0.vpos[9] ),
    .X(net6219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5696 (.A(net3936),
    .X(net6220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5697 (.A(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(net6221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5698 (.A(net2884),
    .X(net6222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5699 (.A(_02776_),
    .X(net6223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(net6380),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5700 (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(net6224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5701 (.A(net1726),
    .X(net6225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5702 (.A(_00807_),
    .X(net6226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5703 (.A(net1792),
    .X(net6227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5704 (.A(\rbzero.spi_registers.buf_sky[3] ),
    .X(net6228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5705 (.A(net1531),
    .X(net6229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5706 (.A(_03247_),
    .X(net6230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5707 (.A(_00805_),
    .X(net6231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5708 (.A(\rbzero.spi_registers.buf_texadd3[5] ),
    .X(net6232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5709 (.A(net1661),
    .X(net6233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(_01352_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5710 (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .X(net6234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5711 (.A(\rbzero.spi_registers.buf_texadd2[5] ),
    .X(net6235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5712 (.A(net1883),
    .X(net6236));
 sky130_fd_sc_hd__buf_2 hold5713 (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(net6237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5714 (.A(_02551_),
    .X(net6238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5715 (.A(_02552_),
    .X(net6239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5716 (.A(_02553_),
    .X(net6240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5717 (.A(_02555_),
    .X(net6241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5718 (.A(_02558_),
    .X(net6242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5719 (.A(net2920),
    .X(net6243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(net5486),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5720 (.A(\rbzero.spi_registers.buf_sky[1] ),
    .X(net6244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5721 (.A(net1595),
    .X(net6245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5722 (.A(_03244_),
    .X(net6246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5723 (.A(_00803_),
    .X(net6247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5724 (.A(net6311),
    .X(net6248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5725 (.A(_06216_),
    .X(net6249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5726 (.A(_02950_),
    .X(net6250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5727 (.A(net6268),
    .X(net6251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5728 (.A(_01613_),
    .X(net6252));
 sky130_fd_sc_hd__buf_2 hold5729 (.A(net692),
    .X(net6253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(net5488),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5730 (.A(_08214_),
    .X(net6254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5731 (.A(\rbzero.spi_registers.buf_texadd2[9] ),
    .X(net6255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5732 (.A(net1806),
    .X(net6256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5733 (.A(\rbzero.spi_registers.buf_texadd1[5] ),
    .X(net6257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5734 (.A(net1604),
    .X(net6258));
 sky130_fd_sc_hd__buf_2 hold5735 (.A(net673),
    .X(net6259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5736 (.A(_08224_),
    .X(net6260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5737 (.A(_00424_),
    .X(net6261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5738 (.A(\rbzero.spi_registers.buf_texadd3[9] ),
    .X(net6262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5739 (.A(net1744),
    .X(net6263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net7645),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5740 (.A(\gpout0.vpos[1] ),
    .X(net6264));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5741 (.A(net3897),
    .X(net6265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5742 (.A(_03949_),
    .X(net6266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5743 (.A(_01252_),
    .X(net6267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5744 (.A(\rbzero.map_rom.f4 ),
    .X(net6268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5745 (.A(\rbzero.map_rom.a6 ),
    .X(net6269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5746 (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(net6270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5747 (.A(net1571),
    .X(net6271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5748 (.A(_00814_),
    .X(net6272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5749 (.A(net2543),
    .X(net6273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(net4414),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5750 (.A(\rbzero.spi_registers.buf_leak[2] ),
    .X(net6274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5751 (.A(net2553),
    .X(net6275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5752 (.A(_03269_),
    .X(net6276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5753 (.A(_00816_),
    .X(net6277));
 sky130_fd_sc_hd__clkbuf_2 hold5754 (.A(net695),
    .X(net6278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5755 (.A(_08217_),
    .X(net6279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5756 (.A(_00422_),
    .X(net6280));
 sky130_fd_sc_hd__clkbuf_2 hold5757 (.A(net656),
    .X(net6281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5758 (.A(_08221_),
    .X(net6282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5759 (.A(_00423_),
    .X(net6283));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold576 (.A(net7569),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5760 (.A(\rbzero.spi_registers.buf_texadd1[9] ),
    .X(net6284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5761 (.A(net1912),
    .X(net6285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5762 (.A(\gpout0.vpos[0] ),
    .X(net6286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5763 (.A(net3964),
    .X(net6287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5764 (.A(\rbzero.map_rom.d6 ),
    .X(net6288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5765 (.A(\rbzero.spi_registers.buf_leak[3] ),
    .X(net6289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5766 (.A(net1735),
    .X(net6290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5767 (.A(_03270_),
    .X(net6291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5768 (.A(_00817_),
    .X(net6292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5769 (.A(\rbzero.spi_registers.buf_leak[4] ),
    .X(net6293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(net4286),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5770 (.A(net2590),
    .X(net6294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5771 (.A(_03271_),
    .X(net6295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5772 (.A(_00818_),
    .X(net6296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5773 (.A(\rbzero.spi_registers.buf_texadd3[0] ),
    .X(net6297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5774 (.A(net1559),
    .X(net6298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5775 (.A(\rbzero.spi_registers.buf_texadd1[0] ),
    .X(net6299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5776 (.A(net1703),
    .X(net6300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5777 (.A(\rbzero.spi_registers.buf_floor[0] ),
    .X(net6301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5778 (.A(net1534),
    .X(net6302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5779 (.A(_03253_),
    .X(net6303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(net6398),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_2 hold5780 (.A(net3197),
    .X(net6304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5781 (.A(_02728_),
    .X(net6305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5782 (.A(\rbzero.spi_registers.mosi ),
    .X(net6306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5783 (.A(net1467),
    .X(net6307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5784 (.A(\rbzero.wall_tracer.mapY[5] ),
    .X(net6308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5785 (.A(net3034),
    .X(net6309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5786 (.A(_02749_),
    .X(net6310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5787 (.A(\rbzero.map_rom.f3 ),
    .X(net6311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5788 (.A(\gpout0.hpos[9] ),
    .X(net6312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5789 (.A(net3991),
    .X(net6313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(net6400),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5790 (.A(_00481_),
    .X(net6314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5791 (.A(\rbzero.tex_g0[32] ),
    .X(net6315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5792 (.A(net633),
    .X(net6316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5793 (.A(_04422_),
    .X(net6317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5794 (.A(net634),
    .X(net6318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5796 (.A(_02944_),
    .X(net6320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5797 (.A(\rbzero.pov.ss_buffer[0] ),
    .X(net6321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5798 (.A(net624),
    .X(net6322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5799 (.A(\rbzero.pov.sclk_buffer[0] ),
    .X(net6323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_01159_),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5800 (.A(net621),
    .X(net6324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5802 (.A(_02625_),
    .X(net6326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5803 (.A(\rbzero.spi_registers.mosi_buffer[0] ),
    .X(net6327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5804 (.A(net627),
    .X(net6328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5805 (.A(\gpout0.vpos[3] ),
    .X(net6329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5806 (.A(net4013),
    .X(net6330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5807 (.A(_01257_),
    .X(net6331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5808 (.A(\rbzero.tex_b0[10] ),
    .X(net6332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5809 (.A(net728),
    .X(net6333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(net5499),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5810 (.A(_04587_),
    .X(net6334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5811 (.A(net729),
    .X(net6335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5812 (.A(\rbzero.tex_b1[6] ),
    .X(net6336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5813 (.A(net760),
    .X(net6337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5814 (.A(_04521_),
    .X(net6338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5815 (.A(net761),
    .X(net6339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5816 (.A(\gpout4.clk_div[1] ),
    .X(net6340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5817 (.A(net1047),
    .X(net6341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5818 (.A(\rbzero.tex_g1[8] ),
    .X(net6342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5819 (.A(net828),
    .X(net6343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(net5501),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5820 (.A(_04378_),
    .X(net6344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5821 (.A(net829),
    .X(net6345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5822 (.A(\gpout5.clk_div[1] ),
    .X(net6346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5823 (.A(net1080),
    .X(net6347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5824 (.A(\gpout0.clk_div[1] ),
    .X(net6348));
 sky130_fd_sc_hd__buf_1 hold5825 (.A(net1127),
    .X(net6349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5826 (.A(\rbzero.tex_b0[20] ),
    .X(net6350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5827 (.A(net1031),
    .X(net6351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5828 (.A(_04576_),
    .X(net6352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5829 (.A(net1032),
    .X(net6353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net6364),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5830 (.A(\gpout2.clk_div[1] ),
    .X(net6354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5831 (.A(net1182),
    .X(net6355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5832 (.A(\gpout3.clk_div[1] ),
    .X(net6356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5833 (.A(net1135),
    .X(net6357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5834 (.A(\rbzero.tex_r1[20] ),
    .X(net6358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5835 (.A(net995),
    .X(net6359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5836 (.A(_04219_),
    .X(net6360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5837 (.A(net996),
    .X(net6361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5838 (.A(\rbzero.spi_registers.sclk_buffer[0] ),
    .X(net6362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5839 (.A(net1172),
    .X(net6363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_03946_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5840 (.A(\rbzero.pov.mosi_buffer[0] ),
    .X(net6364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5841 (.A(net1107),
    .X(net6365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5842 (.A(\rbzero.tex_g1[38] ),
    .X(net6366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5843 (.A(net1061),
    .X(net6367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5844 (.A(_04345_),
    .X(net6368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5845 (.A(net1062),
    .X(net6369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5846 (.A(\rbzero.tex_r1[50] ),
    .X(net6370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5847 (.A(net1040),
    .X(net6371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5848 (.A(_04186_),
    .X(net6372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5849 (.A(net1041),
    .X(net6373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_01251_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5850 (.A(\rbzero.tex_b1[16] ),
    .X(net6374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5851 (.A(net1088),
    .X(net6375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5852 (.A(_04510_),
    .X(net6376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5853 (.A(net1089),
    .X(net6377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5854 (.A(\rbzero.tex_g0[22] ),
    .X(net6378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5855 (.A(net1093),
    .X(net6379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5856 (.A(_04433_),
    .X(net6380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5857 (.A(net1094),
    .X(net6381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5858 (.A(\rbzero.tex_g0[52] ),
    .X(net6382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5859 (.A(net1110),
    .X(net6383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(net6382),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5860 (.A(_04399_),
    .X(net6384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5861 (.A(net1111),
    .X(net6385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5862 (.A(\rbzero.tex_b1[46] ),
    .X(net6386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5863 (.A(net1138),
    .X(net6387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5864 (.A(_04477_),
    .X(net6388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5865 (.A(net1139),
    .X(net6389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5866 (.A(\rbzero.tex_g0[12] ),
    .X(net6390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5867 (.A(net1073),
    .X(net6391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5868 (.A(_04444_),
    .X(net6392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5869 (.A(net1074),
    .X(net6393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(net6384),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5870 (.A(\rbzero.tex_r0[54] ),
    .X(net6394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5871 (.A(net1148),
    .X(net6395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5872 (.A(_04256_),
    .X(net6396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5873 (.A(net1149),
    .X(net6397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5874 (.A(\rbzero.tex_b0[50] ),
    .X(net6398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5875 (.A(net1102),
    .X(net6399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5876 (.A(_04543_),
    .X(net6400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5877 (.A(net1103),
    .X(net6401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5878 (.A(\rbzero.tex_r0[24] ),
    .X(net6402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5879 (.A(net1159),
    .X(net6403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_01382_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5880 (.A(_04289_),
    .X(net6404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5881 (.A(net1160),
    .X(net6405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5882 (.A(\rbzero.tex_r0[34] ),
    .X(net6406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5883 (.A(net1153),
    .X(net6407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5884 (.A(_04278_),
    .X(net6408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5885 (.A(net1154),
    .X(net6409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5886 (.A(\rbzero.tex_g1[58] ),
    .X(net6410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5887 (.A(net1120),
    .X(net6411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5888 (.A(_04322_),
    .X(net6412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5889 (.A(net1121),
    .X(net6413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(net5512),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5890 (.A(\rbzero.tex_g1[18] ),
    .X(net6414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5891 (.A(net1201),
    .X(net6415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5892 (.A(_04367_),
    .X(net6416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5893 (.A(net1202),
    .X(net6417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5894 (.A(\rbzero.tex_r1[30] ),
    .X(net6418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5895 (.A(net1179),
    .X(net6419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5896 (.A(\rbzero.tex_b1[36] ),
    .X(net6420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5897 (.A(net1234),
    .X(net6421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5898 (.A(_04488_),
    .X(net6422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5899 (.A(net1235),
    .X(net6423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(net5514),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5900 (.A(\rbzero.tex_b1[45] ),
    .X(net6424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5901 (.A(net1372),
    .X(net6425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5902 (.A(_04478_),
    .X(net6426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5903 (.A(net1373),
    .X(net6427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5904 (.A(\rbzero.tex_b0[40] ),
    .X(net6428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5905 (.A(net1196),
    .X(net6429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5906 (.A(_04554_),
    .X(net6430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5907 (.A(net1197),
    .X(net6431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5908 (.A(\rbzero.tex_g1[28] ),
    .X(net6432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5909 (.A(net1206),
    .X(net6433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net5761),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5910 (.A(_04356_),
    .X(net6434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5911 (.A(net1207),
    .X(net6435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5912 (.A(\rbzero.tex_r0[14] ),
    .X(net6436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5913 (.A(net1258),
    .X(net6437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5914 (.A(_04300_),
    .X(net6438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5915 (.A(net1259),
    .X(net6439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5916 (.A(\rbzero.tex_b1[56] ),
    .X(net6440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5917 (.A(net1267),
    .X(net6441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5918 (.A(_04466_),
    .X(net6442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5919 (.A(net1268),
    .X(net6443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_03206_),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5920 (.A(\rbzero.tex_r1[10] ),
    .X(net6444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5921 (.A(net1347),
    .X(net6445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5922 (.A(_04230_),
    .X(net6446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5923 (.A(net1348),
    .X(net6447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5924 (.A(\rbzero.tex_g0[42] ),
    .X(net6448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5925 (.A(net1191),
    .X(net6449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5926 (.A(_04411_),
    .X(net6450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5927 (.A(net1192),
    .X(net6451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5928 (.A(\rbzero.tex_r1[0] ),
    .X(net6452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5929 (.A(net1453),
    .X(net6453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(net4195),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5930 (.A(_04240_),
    .X(net6454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5931 (.A(net1454),
    .X(net6455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5932 (.A(\rbzero.tex_g0[28] ),
    .X(net6456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5933 (.A(net1332),
    .X(net6457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5934 (.A(_04427_),
    .X(net6458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5935 (.A(net1333),
    .X(net6459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5936 (.A(\rbzero.tex_b0[6] ),
    .X(net6460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5937 (.A(net1357),
    .X(net6461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5938 (.A(_04591_),
    .X(net6462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5939 (.A(net1358),
    .X(net6463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(net5522),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5940 (.A(\rbzero.tex_r0[44] ),
    .X(net6464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5941 (.A(net1352),
    .X(net6465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5942 (.A(_04267_),
    .X(net6466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5943 (.A(net1353),
    .X(net6467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5944 (.A(\rbzero.tex_b0[46] ),
    .X(net6468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5945 (.A(net1386),
    .X(net6469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5946 (.A(_04547_),
    .X(net6470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5947 (.A(net1387),
    .X(net6471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5948 (.A(\rbzero.tex_b1[0] ),
    .X(net6472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5949 (.A(net1480),
    .X(net6473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(net5524),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5950 (.A(_04526_),
    .X(net6474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5951 (.A(net1481),
    .X(net6475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5952 (.A(\rbzero.tex_b0[30] ),
    .X(net6476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5953 (.A(net1417),
    .X(net6477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5954 (.A(_04565_),
    .X(net6478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5955 (.A(net1418),
    .X(net6479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5956 (.A(\rbzero.tex_g1[0] ),
    .X(net6480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5957 (.A(net1501),
    .X(net6481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5958 (.A(_04385_),
    .X(net6482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5959 (.A(net1502),
    .X(net6483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(net6410),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5960 (.A(\rbzero.tex_g0[62] ),
    .X(net6484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5961 (.A(net1445),
    .X(net6485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5962 (.A(_04388_),
    .X(net6486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5963 (.A(net1446),
    .X(net6487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5964 (.A(\rbzero.tex_r0[49] ),
    .X(net6488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5965 (.A(net1424),
    .X(net6489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5966 (.A(_04261_),
    .X(net6490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5967 (.A(net1425),
    .X(net6491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5968 (.A(\rbzero.tex_b1[32] ),
    .X(net6492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5969 (.A(net1397),
    .X(net6493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net6412),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5970 (.A(_04493_),
    .X(net6494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5971 (.A(net1398),
    .X(net6495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5972 (.A(\rbzero.wall_hot[0] ),
    .X(net6496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5973 (.A(_04639_),
    .X(net6497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5974 (.A(_09944_),
    .X(net6498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5975 (.A(\rbzero.tex_r0[19] ),
    .X(net6499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5976 (.A(net1477),
    .X(net6500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5977 (.A(_04294_),
    .X(net6501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5978 (.A(net1478),
    .X(net6502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5979 (.A(\rbzero.tex_b1[26] ),
    .X(net6503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_01452_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5980 (.A(net1383),
    .X(net6504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5981 (.A(\rbzero.tex_b0[60] ),
    .X(net6505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5982 (.A(net1461),
    .X(net6506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5983 (.A(\rbzero.tex_b0[26] ),
    .X(net6507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5984 (.A(net1442),
    .X(net6508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5985 (.A(_04569_),
    .X(net6509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5986 (.A(net1443),
    .X(net6510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5987 (.A(\rbzero.tex_g1[24] ),
    .X(net6511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5988 (.A(net1427),
    .X(net6512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5989 (.A(_04360_),
    .X(net6513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(net5561),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5990 (.A(net1428),
    .X(net6514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5991 (.A(\rbzero.tex_r1[60] ),
    .X(net6515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5992 (.A(net1464),
    .X(net6516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5993 (.A(_04175_),
    .X(net6517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5994 (.A(net1465),
    .X(net6518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5995 (.A(\rbzero.tex_r1[16] ),
    .X(net6519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5996 (.A(net1448),
    .X(net6520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5997 (.A(_04223_),
    .X(net6521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5998 (.A(net1449),
    .X(net6522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5999 (.A(\rbzero.spi_registers.buf_floor[4] ),
    .X(net6523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(net5563),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6000 (.A(net1540),
    .X(net6524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6001 (.A(_03259_),
    .X(net6525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6002 (.A(\rbzero.tex_g1[12] ),
    .X(net6526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6003 (.A(net1515),
    .X(net6527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6004 (.A(_04373_),
    .X(net6528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6005 (.A(net1516),
    .X(net6529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6006 (.A(\rbzero.tex_r0[10] ),
    .X(net6530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6007 (.A(net1430),
    .X(net6531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6008 (.A(_04304_),
    .X(net6532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6009 (.A(net1431),
    .X(net6533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(net3584),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6010 (.A(\rbzero.tex_b0[35] ),
    .X(net6534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6011 (.A(net1497),
    .X(net6535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6012 (.A(_04559_),
    .X(net6536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6013 (.A(net1498),
    .X(net6537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6014 (.A(\rbzero.tex_b1[22] ),
    .X(net6538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6015 (.A(net1435),
    .X(net6539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6016 (.A(_04504_),
    .X(net6540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6017 (.A(net1436),
    .X(net6541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6018 (.A(\rbzero.tex_g0[57] ),
    .X(net6542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6019 (.A(net1526),
    .X(net6543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(net5475),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6020 (.A(_04394_),
    .X(net6544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6021 (.A(net1527),
    .X(net6545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6022 (.A(\rbzero.tex_b1[62] ),
    .X(net6546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6023 (.A(net1518),
    .X(net6547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6024 (.A(\rbzero.spi_registers.buf_texadd3[15] ),
    .X(net6548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6025 (.A(net1543),
    .X(net6549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6026 (.A(\rbzero.tex_g1[35] ),
    .X(net6550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6027 (.A(net1512),
    .X(net6551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6028 (.A(_04348_),
    .X(net6552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6029 (.A(net1513),
    .X(net6553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(net6348),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6030 (.A(\gpout1.clk_div[1] ),
    .X(net6554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6031 (.A(net1920),
    .X(net6555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6032 (.A(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(net6556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6033 (.A(net1577),
    .X(net6557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6034 (.A(\rbzero.spi_registers.buf_floor[2] ),
    .X(net6558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6035 (.A(net1615),
    .X(net6559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6036 (.A(_03256_),
    .X(net6560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6037 (.A(\rbzero.spi_registers.buf_texadd1[12] ),
    .X(net6561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6038 (.A(net1625),
    .X(net6562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6039 (.A(\rbzero.tex_r1[45] ),
    .X(net6563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_04142_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6040 (.A(net1628),
    .X(net6564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6041 (.A(_04191_),
    .X(net6565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6042 (.A(net1629),
    .X(net6566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6043 (.A(\rbzero.spi_registers.buf_texadd2[1] ),
    .X(net6567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6044 (.A(net1909),
    .X(net6568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6045 (.A(\rbzero.tex_g0[3] ),
    .X(net6569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6046 (.A(net1610),
    .X(net6570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6047 (.A(_04454_),
    .X(net6571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6048 (.A(net1611),
    .X(net6572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6049 (.A(\rbzero.tex_g0[47] ),
    .X(net6573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_01635_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6050 (.A(net1641),
    .X(net6574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6051 (.A(_04406_),
    .X(net6575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6052 (.A(net1642),
    .X(net6576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6053 (.A(\rbzero.tex_r0[39] ),
    .X(net6577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6054 (.A(net1551),
    .X(net6578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6055 (.A(_04272_),
    .X(net6579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6056 (.A(net1552),
    .X(net6580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6057 (.A(\rbzero.tex_g1[30] ),
    .X(net6581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6058 (.A(net1680),
    .X(net6582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6059 (.A(_04353_),
    .X(net6583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net4886),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6060 (.A(net1681),
    .X(net6584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6061 (.A(\rbzero.spi_registers.buf_texadd1[11] ),
    .X(net6585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6062 (.A(net1647),
    .X(net6586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6063 (.A(\rbzero.spi_registers.buf_texadd1[13] ),
    .X(net6587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6064 (.A(net1692),
    .X(net6588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6065 (.A(\rbzero.spi_registers.buf_texadd3[3] ),
    .X(net6589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6066 (.A(net1686),
    .X(net6590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6067 (.A(\rbzero.tex_b0[41] ),
    .X(net6591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6068 (.A(net1824),
    .X(net6592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6069 (.A(\rbzero.tex_b1[55] ),
    .X(net6593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(net4888),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6070 (.A(net1485),
    .X(net6594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6071 (.A(_04467_),
    .X(net6595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6072 (.A(net1486),
    .X(net6596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6073 (.A(\rbzero.tex_b0[9] ),
    .X(net6597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6074 (.A(net1620),
    .X(net6598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6075 (.A(_04588_),
    .X(net6599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6076 (.A(net1621),
    .X(net6600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6077 (.A(\rbzero.spi_registers.buf_texadd1[1] ),
    .X(net6601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6078 (.A(net1652),
    .X(net6602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6079 (.A(\rbzero.tex_r0[28] ),
    .X(net6603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(net1637),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6080 (.A(net1664),
    .X(net6604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6081 (.A(_04284_),
    .X(net6605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6082 (.A(net1665),
    .X(net6606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6083 (.A(\rbzero.spi_registers.buf_texadd1[3] ),
    .X(net6607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6084 (.A(net1667),
    .X(net6608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6085 (.A(\rbzero.tex_g0[37] ),
    .X(net6609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6086 (.A(net1877),
    .X(net6610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6087 (.A(_04417_),
    .X(net6611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6088 (.A(net1878),
    .X(net6612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6089 (.A(\rbzero.tex_b0[53] ),
    .X(net6613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_03202_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6090 (.A(net1738),
    .X(net6614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6091 (.A(_04539_),
    .X(net6615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6092 (.A(net1739),
    .X(net6616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6093 (.A(\rbzero.tex_g0[49] ),
    .X(net6617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6094 (.A(net1658),
    .X(net6618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6095 (.A(_04402_),
    .X(net6619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6096 (.A(net1659),
    .X(net6620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6097 (.A(\rbzero.spi_registers.buf_texadd1[18] ),
    .X(net6621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6098 (.A(net1729),
    .X(net6622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6099 (.A(\rbzero.spi_registers.buf_texadd3[1] ),
    .X(net6623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(net4171),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6100 (.A(net1903),
    .X(net6624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6101 (.A(\rbzero.tex_r1[35] ),
    .X(net6625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6102 (.A(net1891),
    .X(net6626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6103 (.A(_04202_),
    .X(net6627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6104 (.A(net1892),
    .X(net6628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6105 (.A(\rbzero.spi_registers.buf_texadd1[4] ),
    .X(net6629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6106 (.A(net1829),
    .X(net6630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6107 (.A(\rbzero.tex_r0[23] ),
    .X(net6631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6108 (.A(net1777),
    .X(net6632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6109 (.A(_04290_),
    .X(net6633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(net6356),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6110 (.A(net1778),
    .X(net6634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6111 (.A(\rbzero.tex_g1[15] ),
    .X(net6635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6112 (.A(net1706),
    .X(net6636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6113 (.A(_04370_),
    .X(net6637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6114 (.A(net1707),
    .X(net6638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6115 (.A(\rbzero.tex_g0[13] ),
    .X(net6639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6116 (.A(net1888),
    .X(net6640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6117 (.A(\rbzero.tex_r1[23] ),
    .X(net6641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6118 (.A(net1747),
    .X(net6642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6119 (.A(_04216_),
    .X(net6643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_04157_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6120 (.A(net1748),
    .X(net6644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6121 (.A(\rbzero.tex_g1[17] ),
    .X(net6645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6122 (.A(net1771),
    .X(net6646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6123 (.A(_04368_),
    .X(net6647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6124 (.A(net1772),
    .X(net6648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6125 (.A(\rbzero.spi_registers.buf_texadd3[13] ),
    .X(net6649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6126 (.A(net1718),
    .X(net6650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6127 (.A(\rbzero.tex_r0[53] ),
    .X(net6651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6128 (.A(net1723),
    .X(net6652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6129 (.A(_04257_),
    .X(net6653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_01649_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6130 (.A(net1724),
    .X(net6654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6131 (.A(\rbzero.tex_g0[9] ),
    .X(net6655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6132 (.A(net1715),
    .X(net6656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6133 (.A(_04447_),
    .X(net6657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6134 (.A(net1716),
    .X(net6658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6135 (.A(\rbzero.spi_registers.buf_texadd3[6] ),
    .X(net6659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6136 (.A(net1964),
    .X(net6660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6137 (.A(\rbzero.spi_registers.buf_texadd2[4] ),
    .X(net6661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6138 (.A(net2113),
    .X(net6662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6139 (.A(\rbzero.tex_g0[23] ),
    .X(net6663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(net6386),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6140 (.A(net1674),
    .X(net6664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6141 (.A(\rbzero.tex_g0[26] ),
    .X(net6665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6142 (.A(net1944),
    .X(net6666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6143 (.A(_04429_),
    .X(net6667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6144 (.A(net1945),
    .X(net6668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6145 (.A(\rbzero.tex_g0[17] ),
    .X(net6669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6146 (.A(net1850),
    .X(net6670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6147 (.A(_04439_),
    .X(net6671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6148 (.A(net1851),
    .X(net6672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6149 (.A(\rbzero.tex_r0[21] ),
    .X(net6673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(net6388),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6150 (.A(net1841),
    .X(net6674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6151 (.A(_04292_),
    .X(net6675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6152 (.A(net1842),
    .X(net6676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6153 (.A(\rbzero.tex_g0[41] ),
    .X(net6677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6154 (.A(net1765),
    .X(net6678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6155 (.A(_04412_),
    .X(net6679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6156 (.A(net1766),
    .X(net6680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6157 (.A(\rbzero.spi_registers.buf_texadd2[2] ),
    .X(net6681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6158 (.A(net1787),
    .X(net6682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6159 (.A(\rbzero.tex_g0[55] ),
    .X(net6683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_01312_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6160 (.A(net1797),
    .X(net6684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6161 (.A(_04396_),
    .X(net6685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6162 (.A(net1798),
    .X(net6686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6163 (.A(\rbzero.tex_r1[43] ),
    .X(net6687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6164 (.A(net1853),
    .X(net6688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6165 (.A(_04194_),
    .X(net6689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6166 (.A(net1854),
    .X(net6690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6167 (.A(\rbzero.tex_b0[61] ),
    .X(net6691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6168 (.A(net1906),
    .X(net6692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6169 (.A(\rbzero.spi_registers.buf_texadd3[2] ),
    .X(net6693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(net5753),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6170 (.A(net1709),
    .X(net6694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6171 (.A(\rbzero.tex_b1[17] ),
    .X(net6695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6172 (.A(net1800),
    .X(net6696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6173 (.A(\rbzero.tex_r0[13] ),
    .X(net6697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6174 (.A(net2063),
    .X(net6698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6175 (.A(_04301_),
    .X(net6699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6176 (.A(net2064),
    .X(net6700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6177 (.A(\rbzero.tex_r0[15] ),
    .X(net6701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6178 (.A(net1973),
    .X(net6702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6179 (.A(\rbzero.tex_r0[41] ),
    .X(net6703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_03076_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6180 (.A(net1677),
    .X(net6704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6181 (.A(_04270_),
    .X(net6705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6182 (.A(net1678),
    .X(net6706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6183 (.A(\rbzero.tex_b1[19] ),
    .X(net6707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6184 (.A(net1838),
    .X(net6708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6185 (.A(_04507_),
    .X(net6709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6186 (.A(net1839),
    .X(net6710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6187 (.A(\rbzero.tex_r0[25] ),
    .X(net6711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6188 (.A(net2054),
    .X(net6712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6189 (.A(\rbzero.tex_r0[45] ),
    .X(net6713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(net4198),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6190 (.A(net1732),
    .X(net6714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6191 (.A(\rbzero.tex_g0[20] ),
    .X(net6715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6192 (.A(net1917),
    .X(net6716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6193 (.A(_04435_),
    .X(net6717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6194 (.A(net1918),
    .X(net6718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6195 (.A(\rbzero.spi_registers.buf_texadd3[4] ),
    .X(net6719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6196 (.A(net1871),
    .X(net6720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6197 (.A(\rbzero.spi_registers.buf_texadd3[18] ),
    .X(net6721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6198 (.A(net1847),
    .X(net6722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6199 (.A(\rbzero.tex_b0[45] ),
    .X(net6723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(net4935),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6200 (.A(net1753),
    .X(net6724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6201 (.A(_04548_),
    .X(net6725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6202 (.A(net1754),
    .X(net6726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6203 (.A(\rbzero.tex_b0[42] ),
    .X(net6727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6204 (.A(net2390),
    .X(net6728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6205 (.A(\rbzero.spi_registers.buf_texadd1[6] ),
    .X(net6729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6206 (.A(net2274),
    .X(net6730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6207 (.A(\rbzero.tex_b0[14] ),
    .X(net6731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6208 (.A(net1947),
    .X(net6732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6209 (.A(_04582_),
    .X(net6733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(net4525),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6210 (.A(net1948),
    .X(net6734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6211 (.A(\rbzero.tex_b1[41] ),
    .X(net6735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6212 (.A(net1856),
    .X(net6736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6213 (.A(_04483_),
    .X(net6737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6214 (.A(net1924),
    .X(net6738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6215 (.A(\rbzero.spi_registers.buf_texadd2[3] ),
    .X(net6739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6216 (.A(net1868),
    .X(net6740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6217 (.A(\rbzero.tex_b0[51] ),
    .X(net6741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6218 (.A(net1815),
    .X(net6742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6219 (.A(\rbzero.tex_r0[29] ),
    .X(net6743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(net5546),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6220 (.A(net1759),
    .X(net6744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6221 (.A(\rbzero.tex_b0[37] ),
    .X(net6745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6222 (.A(net2073),
    .X(net6746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6223 (.A(_04557_),
    .X(net6747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6224 (.A(net2074),
    .X(net6748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6225 (.A(\rbzero.tex_b1[44] ),
    .X(net6749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6226 (.A(net2188),
    .X(net6750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6227 (.A(\rbzero.tex_g1[42] ),
    .X(net6751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6228 (.A(net2017),
    .X(net6752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6229 (.A(_04340_),
    .X(net6753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(net5548),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6230 (.A(net2018),
    .X(net6754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6231 (.A(\rbzero.tex_g0[4] ),
    .X(net6755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6232 (.A(net2349),
    .X(net6756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6233 (.A(\rbzero.tex_b1[18] ),
    .X(net6757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6234 (.A(net1880),
    .X(net6758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6235 (.A(\rbzero.tex_r1[32] ),
    .X(net6759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6236 (.A(net1774),
    .X(net6760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6237 (.A(_04206_),
    .X(net6761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6238 (.A(net1775),
    .X(net6762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6239 (.A(\rbzero.tex_b1[54] ),
    .X(net6763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(net6394),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6240 (.A(net2149),
    .X(net6764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6241 (.A(_04468_),
    .X(net6765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6242 (.A(net2150),
    .X(net6766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6243 (.A(\rbzero.tex_g1[13] ),
    .X(net6767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6244 (.A(net1741),
    .X(net6768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6245 (.A(\rbzero.tex_g0[29] ),
    .X(net6769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6246 (.A(net2048),
    .X(net6770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6247 (.A(\rbzero.tex_r0[43] ),
    .X(net6771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6248 (.A(net2304),
    .X(net6772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6249 (.A(_04268_),
    .X(net6773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(net6396),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6250 (.A(net2305),
    .X(net6774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6251 (.A(\rbzero.tex_b1[33] ),
    .X(net6775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6252 (.A(net1809),
    .X(net6776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6253 (.A(\rbzero.tex_g1[4] ),
    .X(net6777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6254 (.A(net1979),
    .X(net6778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6255 (.A(\rbzero.tex_b1[4] ),
    .X(net6779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6256 (.A(net2104),
    .X(net6780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6257 (.A(\rbzero.tex_r1[44] ),
    .X(net6781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6258 (.A(net2224),
    .X(net6782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6259 (.A(\rbzero.spi_registers.buf_texadd2[18] ),
    .X(net6783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_01512_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6260 (.A(net2020),
    .X(net6784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6261 (.A(\rbzero.tex_r1[22] ),
    .X(net6785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6262 (.A(net2328),
    .X(net6786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6263 (.A(_04217_),
    .X(net6787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6264 (.A(net2329),
    .X(net6788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6265 (.A(\rbzero.tex_b1[34] ),
    .X(net6789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6266 (.A(net2206),
    .X(net6790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6267 (.A(\rbzero.tex_g0[7] ),
    .X(net6791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6268 (.A(net1794),
    .X(net6792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6269 (.A(_04450_),
    .X(net6793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(net5526),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6270 (.A(net1795),
    .X(net6794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6271 (.A(\rbzero.tex_r0[30] ),
    .X(net6795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6272 (.A(net2060),
    .X(net6796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6273 (.A(\rbzero.tex_b0[4] ),
    .X(net6797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6274 (.A(net1803),
    .X(net6798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6275 (.A(_04593_),
    .X(net6799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6276 (.A(net1804),
    .X(net6800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6277 (.A(\rbzero.tex_g0[53] ),
    .X(net6801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6278 (.A(net1897),
    .X(net6802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6279 (.A(\rbzero.tex_b0[27] ),
    .X(net6803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(net5528),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6280 (.A(net2277),
    .X(net6804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6281 (.A(\rbzero.tex_b0[24] ),
    .X(net6805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6282 (.A(net2481),
    .X(net6806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6283 (.A(_04571_),
    .X(net6807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6284 (.A(net2482),
    .X(net6808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6285 (.A(\rbzero.tex_b1[8] ),
    .X(net6809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6286 (.A(net2605),
    .X(net6810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6287 (.A(_04519_),
    .X(net6811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6288 (.A(net2606),
    .X(net6812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6289 (.A(\rbzero.tex_b1[52] ),
    .X(net6813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(net6406),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6290 (.A(net2433),
    .X(net6814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6291 (.A(_04471_),
    .X(net6815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6292 (.A(net2434),
    .X(net6816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6293 (.A(\rbzero.tex_r1[49] ),
    .X(net6817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6294 (.A(net2066),
    .X(net6818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6295 (.A(_04187_),
    .X(net6819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6296 (.A(net2067),
    .X(net6820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6297 (.A(\rbzero.tex_b0[31] ),
    .X(net6821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6298 (.A(net1894),
    .X(net6822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6299 (.A(\rbzero.tex_r0[9] ),
    .X(net6823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(net6408),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6300 (.A(net2107),
    .X(net6824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6301 (.A(_04305_),
    .X(net6825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6302 (.A(net2108),
    .X(net6826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6303 (.A(\rbzero.tex_r0[37] ),
    .X(net6827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6304 (.A(net1818),
    .X(net6828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6305 (.A(_04274_),
    .X(net6829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6306 (.A(net1819),
    .X(net6830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6307 (.A(\rbzero.tex_b0[29] ),
    .X(net6831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6308 (.A(net2295),
    .X(net6832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6309 (.A(_04566_),
    .X(net6833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_01492_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6310 (.A(net2296),
    .X(net6834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6311 (.A(\rbzero.tex_g1[25] ),
    .X(net6835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6312 (.A(net1821),
    .X(net6836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6313 (.A(\rbzero.tex_b0[34] ),
    .X(net6837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6314 (.A(net2331),
    .X(net6838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6315 (.A(_04560_),
    .X(net6839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6316 (.A(net2332),
    .X(net6840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6317 (.A(\rbzero.tex_b1[47] ),
    .X(net6841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6318 (.A(net2200),
    .X(net6842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6319 (.A(\rbzero.tex_g0[24] ),
    .X(net6843));
 sky130_fd_sc_hd__buf_1 hold632 (.A(\rbzero.pov.ready_buffer[60] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6320 (.A(net2360),
    .X(net6844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6321 (.A(\rbzero.tex_b0[54] ),
    .X(net6845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6322 (.A(net2146),
    .X(net6846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6323 (.A(\rbzero.tex_r1[41] ),
    .X(net6847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6324 (.A(net2082),
    .X(net6848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6325 (.A(\rbzero.tex_g1[29] ),
    .X(net6849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6326 (.A(net1697),
    .X(net6850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6327 (.A(\rbzero.tex_r1[21] ),
    .X(net6851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6328 (.A(net2007),
    .X(net6852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6329 (.A(\rbzero.spi_registers.buf_texadd1[2] ),
    .X(net6853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_03487_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6330 (.A(net2076),
    .X(net6854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6331 (.A(\rbzero.tex_g1[20] ),
    .X(net6855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6332 (.A(net2240),
    .X(net6856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6333 (.A(_04364_),
    .X(net6857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6334 (.A(net2241),
    .X(net6858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6335 (.A(\rbzero.tex_b1[9] ),
    .X(net6859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6336 (.A(net2319),
    .X(net6860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6337 (.A(\rbzero.tex_b1[13] ),
    .X(net6861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6338 (.A(net2340),
    .X(net6862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6339 (.A(_04513_),
    .X(net6863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(net4307),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6340 (.A(net2341),
    .X(net6864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6341 (.A(\rbzero.tex_r0[20] ),
    .X(net6865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6342 (.A(net2376),
    .X(net6866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6343 (.A(\rbzero.tex_r1[9] ),
    .X(net6867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6344 (.A(net1900),
    .X(net6868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6345 (.A(_04231_),
    .X(net6869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6346 (.A(net1901),
    .X(net6870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6347 (.A(\rbzero.tex_b0[33] ),
    .X(net6871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6348 (.A(net2027),
    .X(net6872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6349 (.A(_04561_),
    .X(net6873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(net6402),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6350 (.A(net2028),
    .X(net6874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6351 (.A(\rbzero.tex_g1[16] ),
    .X(net6875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6352 (.A(net2134),
    .X(net6876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6353 (.A(\rbzero.tex_g0[50] ),
    .X(net6877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6354 (.A(net1995),
    .X(net6878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6355 (.A(\rbzero.tex_r1[13] ),
    .X(net6879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6356 (.A(net1683),
    .X(net6880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6357 (.A(_04226_),
    .X(net6881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6358 (.A(net2086),
    .X(net6882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6359 (.A(\rbzero.tex_b1[59] ),
    .X(net6883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net6404),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6360 (.A(net2140),
    .X(net6884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6361 (.A(_04463_),
    .X(net6885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6362 (.A(net2213),
    .X(net6886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6363 (.A(\rbzero.tex_b0[38] ),
    .X(net6887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6364 (.A(net2581),
    .X(net6888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6365 (.A(\rbzero.tex_g1[34] ),
    .X(net6889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6366 (.A(net2125),
    .X(net6890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6367 (.A(\rbzero.tex_g0[14] ),
    .X(net6891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6368 (.A(net1985),
    .X(net6892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6369 (.A(\rbzero.tex_g1[22] ),
    .X(net6893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_01482_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6370 (.A(net2524),
    .X(net6894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6371 (.A(_04362_),
    .X(net6895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6372 (.A(net2525),
    .X(net6896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6373 (.A(\rbzero.tex_r1[7] ),
    .X(net6897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6374 (.A(net2079),
    .X(net6898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6375 (.A(_04233_),
    .X(net6899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6376 (.A(net2080),
    .X(net6900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6377 (.A(\rbzero.tex_r1[61] ),
    .X(net6901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6378 (.A(net1835),
    .X(net6902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6379 (.A(\rbzero.tex_g1[54] ),
    .X(net6903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(net5584),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6380 (.A(net2334),
    .X(net6904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6381 (.A(\rbzero.tex_r1[48] ),
    .X(net6905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6382 (.A(net2469),
    .X(net6906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6383 (.A(_04188_),
    .X(net6907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6384 (.A(net2470),
    .X(net6908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6385 (.A(\rbzero.tex_r1[51] ),
    .X(net6909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6386 (.A(net2137),
    .X(net6910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6387 (.A(\rbzero.tex_b1[35] ),
    .X(net6911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6388 (.A(net2227),
    .X(net6912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6389 (.A(\rbzero.tex_g0[30] ),
    .X(net6913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(net5586),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6390 (.A(net2402),
    .X(net6914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6391 (.A(\rbzero.tex_g1[62] ),
    .X(net6915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6392 (.A(net2110),
    .X(net6916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6393 (.A(_04317_),
    .X(net6917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6394 (.A(net2111),
    .X(net6918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6395 (.A(\rbzero.tex_b0[3] ),
    .X(net6919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6396 (.A(net2370),
    .X(net6920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6397 (.A(\rbzero.tex_r0[3] ),
    .X(net6921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6398 (.A(net2163),
    .X(net6922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6399 (.A(\rbzero.tex_g0[31] ),
    .X(net6923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net5820),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(net5503),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6400 (.A(net2313),
    .X(net6924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6401 (.A(\rbzero.tex_b1[20] ),
    .X(net6925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6402 (.A(net2166),
    .X(net6926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6403 (.A(\rbzero.spi_registers.buf_texadd1[14] ),
    .X(net6927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6404 (.A(net2593),
    .X(net6928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6405 (.A(\rbzero.tex_g1[43] ),
    .X(net6929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6406 (.A(net2209),
    .X(net6930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6407 (.A(\rbzero.tex_g0[51] ),
    .X(net6931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6408 (.A(net1950),
    .X(net6932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6409 (.A(\rbzero.tex_b0[28] ),
    .X(net6933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(net5505),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6410 (.A(net2430),
    .X(net6934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6411 (.A(\rbzero.tex_r0[42] ),
    .X(net6935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6412 (.A(net2421),
    .X(net6936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6413 (.A(\rbzero.tex_b1[14] ),
    .X(net6937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6414 (.A(net2584),
    .X(net6938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6415 (.A(\rbzero.tex_g0[43] ),
    .X(net6939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6416 (.A(net2218),
    .X(net6940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6417 (.A(\rbzero.tex_r1[24] ),
    .X(net6941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6418 (.A(net2373),
    .X(net6942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6419 (.A(\rbzero.tex_r0[33] ),
    .X(net6943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(net4502),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6420 (.A(net2445),
    .X(net6944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6421 (.A(_04279_),
    .X(net6945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6422 (.A(net2446),
    .X(net6946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6423 (.A(\rbzero.tex_b0[23] ),
    .X(net6947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6424 (.A(net2030),
    .X(net6948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6425 (.A(_04572_),
    .X(net6949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6426 (.A(net2031),
    .X(net6950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6427 (.A(\rbzero.tex_b0[17] ),
    .X(net6951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6428 (.A(net2268),
    .X(net6952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6429 (.A(_04579_),
    .X(net6953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(net4504),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6430 (.A(net2269),
    .X(net6954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6431 (.A(\rbzero.tex_b0[36] ),
    .X(net6955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6432 (.A(net2051),
    .X(net6956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6433 (.A(\rbzero.tex_g1[7] ),
    .X(net6957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6434 (.A(net2514),
    .X(net6958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6435 (.A(_04379_),
    .X(net6959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6436 (.A(net2515),
    .X(net6960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6437 (.A(\rbzero.tex_g0[39] ),
    .X(net6961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6438 (.A(net1812),
    .X(net6962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6439 (.A(_04414_),
    .X(net6963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(net5565),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6440 (.A(net1813),
    .X(net6964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6441 (.A(\rbzero.tex_g0[16] ),
    .X(net6965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6442 (.A(net1935),
    .X(net6966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6443 (.A(_04440_),
    .X(net6967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6444 (.A(net1936),
    .X(net6968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6445 (.A(\rbzero.tex_b0[18] ),
    .X(net6969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6446 (.A(net2511),
    .X(net6970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6447 (.A(\rbzero.tex_b1[49] ),
    .X(net6971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6448 (.A(net2285),
    .X(net6972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6449 (.A(_04474_),
    .X(net6973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(net5567),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6450 (.A(net2286),
    .X(net6974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6451 (.A(\rbzero.tex_b0[47] ),
    .X(net6975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6452 (.A(net1961),
    .X(net6976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6453 (.A(\rbzero.tex_b0[15] ),
    .X(net6977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6454 (.A(net2608),
    .X(net6978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6455 (.A(\rbzero.tex_g0[10] ),
    .X(net6979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6456 (.A(net2116),
    .X(net6980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6457 (.A(\rbzero.tex_g1[26] ),
    .X(net6981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6458 (.A(net1865),
    .X(net6982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6459 (.A(\rbzero.tex_b0[7] ),
    .X(net6983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(net3589),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6460 (.A(net2408),
    .X(net6984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6461 (.A(\rbzero.tex_g1[14] ),
    .X(net6985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6462 (.A(net2004),
    .X(net6986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6463 (.A(\rbzero.tex_g1[61] ),
    .X(net6987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6464 (.A(net2057),
    .X(net6988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6465 (.A(_04318_),
    .X(net6989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6466 (.A(net2058),
    .X(net6990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6467 (.A(\rbzero.tex_r0[11] ),
    .X(net6991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6468 (.A(net2143),
    .X(net6992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6469 (.A(\rbzero.tex_g0[46] ),
    .X(net6993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(net5612),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6470 (.A(net2550),
    .X(net6994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6471 (.A(_04407_),
    .X(net6995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6472 (.A(net2551),
    .X(net6996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6473 (.A(\rbzero.tex_g0[59] ),
    .X(net6997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6474 (.A(net2301),
    .X(net6998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6475 (.A(_04391_),
    .X(net6999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6476 (.A(net2302),
    .X(net7000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6477 (.A(\rbzero.tex_b1[7] ),
    .X(net7001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6478 (.A(net2653),
    .X(net7002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6479 (.A(\rbzero.tex_r0[60] ),
    .X(net7003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(net6362),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6480 (.A(net1953),
    .X(net7004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6481 (.A(\rbzero.tex_r1[46] ),
    .X(net7005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6482 (.A(net2379),
    .X(net7006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6483 (.A(_04189_),
    .X(net7007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6484 (.A(net2406),
    .X(net7008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6485 (.A(\rbzero.tex_b0[8] ),
    .X(net7009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6486 (.A(net2215),
    .X(net7010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6487 (.A(\rbzero.tex_g0[60] ),
    .X(net7011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6488 (.A(net2131),
    .X(net7012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6489 (.A(\rbzero.tex_b0[43] ),
    .X(net7013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(_03978_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6490 (.A(net2530),
    .X(net7014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6491 (.A(\rbzero.tex_g0[11] ),
    .X(net7015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6492 (.A(net1750),
    .X(net7016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6493 (.A(\rbzero.tex_r0[61] ),
    .X(net7017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6494 (.A(net1932),
    .X(net7018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6495 (.A(\rbzero.tex_b1[5] ),
    .X(net7019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6496 (.A(net2436),
    .X(net7020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6497 (.A(\rbzero.tex_g1[10] ),
    .X(net7021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6498 (.A(net2547),
    .X(net7022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6499 (.A(_04375_),
    .X(net7023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net5822),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_01265_),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6500 (.A(net2548),
    .X(net7024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6501 (.A(\rbzero.tex_r1[62] ),
    .X(net7025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6502 (.A(net2262),
    .X(net7026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6503 (.A(\rbzero.tex_g0[36] ),
    .X(net7027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6504 (.A(net2237),
    .X(net7028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6505 (.A(\rbzero.tex_b0[39] ),
    .X(net7029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6506 (.A(net2399),
    .X(net7030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6507 (.A(\rbzero.tex_g0[27] ),
    .X(net7031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6508 (.A(net2527),
    .X(net7032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6509 (.A(\rbzero.tex_g1[36] ),
    .X(net7033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(net3475),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6510 (.A(net2045),
    .X(net7034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6511 (.A(\rbzero.tex_r0[22] ),
    .X(net7035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6512 (.A(net2475),
    .X(net7036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6513 (.A(\rbzero.tex_b0[56] ),
    .X(net7037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6514 (.A(net2160),
    .X(net7038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6515 (.A(_04536_),
    .X(net7039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6516 (.A(net2161),
    .X(net7040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6517 (.A(\rbzero.tex_b1[50] ),
    .X(net7041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6518 (.A(net2322),
    .X(net7042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6519 (.A(\rbzero.tex_r1[42] ),
    .X(net7043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(net4854),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6520 (.A(net2298),
    .X(net7044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6521 (.A(\rbzero.tex_b1[51] ),
    .X(net7045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6522 (.A(net2249),
    .X(net7046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6523 (.A(\rbzero.tex_b0[21] ),
    .X(net7047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6524 (.A(net2203),
    .X(net7048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6525 (.A(\rbzero.tex_g0[15] ),
    .X(net7049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6526 (.A(net2271),
    .X(net7050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6527 (.A(\rbzero.tex_g1[19] ),
    .X(net7051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6528 (.A(net2357),
    .X(net7052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6529 (.A(\rbzero.tex_b1[30] ),
    .X(net7053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(net3465),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6530 (.A(net2185),
    .X(net7054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6531 (.A(\rbzero.tex_r1[33] ),
    .X(net7055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6532 (.A(net2343),
    .X(net7056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6533 (.A(\rbzero.tex_r0[16] ),
    .X(net7057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6534 (.A(net2010),
    .X(net7058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6535 (.A(\rbzero.tex_r0[57] ),
    .X(net7059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6536 (.A(net2505),
    .X(net7060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6537 (.A(_04252_),
    .X(net7061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6538 (.A(net2506),
    .X(net7062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6539 (.A(\rbzero.tex_g0[58] ),
    .X(net7063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_01049_),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6540 (.A(net2439),
    .X(net7064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6541 (.A(\rbzero.tex_r0[5] ),
    .X(net7065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6542 (.A(net2385),
    .X(net7066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6543 (.A(_04309_),
    .X(net7067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6544 (.A(\rbzero.tex_r0[17] ),
    .X(net7068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6545 (.A(net2040),
    .X(net7069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6546 (.A(\rbzero.tex_g0[5] ),
    .X(net7070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6547 (.A(net1926),
    .X(net7071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6548 (.A(\rbzero.tex_r1[8] ),
    .X(net7072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6549 (.A(net2221),
    .X(net7073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(net6418),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6550 (.A(\rbzero.tex_g1[49] ),
    .X(net7074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6551 (.A(net2246),
    .X(net7075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6552 (.A(_04330_),
    .X(net7076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6553 (.A(net2247),
    .X(net7077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6554 (.A(\rbzero.tex_r0[52] ),
    .X(net7078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6555 (.A(net1976),
    .X(net7079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6556 (.A(_04258_),
    .X(net7080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6557 (.A(net1977),
    .X(net7081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6558 (.A(\rbzero.tex_g0[25] ),
    .X(net7082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6559 (.A(net2128),
    .X(net7083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_04208_),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6560 (.A(\rbzero.tex_r0[12] ),
    .X(net7084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6561 (.A(net2458),
    .X(net7085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6562 (.A(\rbzero.tex_b0[62] ),
    .X(net7086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6563 (.A(net2415),
    .X(net7087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6564 (.A(\rbzero.tex_r1[5] ),
    .X(net7088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6565 (.A(net1458),
    .X(net7089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6566 (.A(_04234_),
    .X(net7090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6567 (.A(net2383),
    .X(net7091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6568 (.A(\rbzero.tex_g0[6] ),
    .X(net7092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6569 (.A(net2616),
    .X(net7093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_01552_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6570 (.A(\rbzero.tex_g0[44] ),
    .X(net7094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6571 (.A(net2265),
    .X(net7095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6572 (.A(\rbzero.tex_b1[38] ),
    .X(net7096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6573 (.A(net2596),
    .X(net7097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6574 (.A(\rbzero.tex_g0[56] ),
    .X(net7098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6575 (.A(net2659),
    .X(net7099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6576 (.A(\rbzero.tex_g1[40] ),
    .X(net7100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6577 (.A(net2310),
    .X(net7101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6578 (.A(_04342_),
    .X(net7102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6579 (.A(net2311),
    .X(net7103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(net6354),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6580 (.A(\rbzero.tex_g1[9] ),
    .X(net7104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6581 (.A(net2478),
    .X(net7105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6582 (.A(\rbzero.tex_b1[37] ),
    .X(net7106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6583 (.A(net2587),
    .X(net7107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6584 (.A(\rbzero.tex_g1[21] ),
    .X(net7108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6585 (.A(net2638),
    .X(net7109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6586 (.A(\rbzero.tex_g0[8] ),
    .X(net7110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6587 (.A(net2521),
    .X(net7111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6588 (.A(\rbzero.tex_g0[40] ),
    .X(net7112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6589 (.A(net2424),
    .X(net7113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_04156_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6590 (.A(\rbzero.tex_r0[8] ),
    .X(net7114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6591 (.A(net2292),
    .X(net7115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6592 (.A(_04306_),
    .X(net7116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6593 (.A(net2293),
    .X(net7117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6594 (.A(\rbzero.tex_b1[58] ),
    .X(net7118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6595 (.A(net2212),
    .X(net7119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6596 (.A(\rbzero.tex_r0[58] ),
    .X(net7120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6597 (.A(net2679),
    .X(net7121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6598 (.A(\rbzero.tex_b0[48] ),
    .X(net7122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6599 (.A(net2502),
    .X(net7123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_01562_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_01647_),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6600 (.A(\rbzero.tex_b0[22] ),
    .X(net7124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6601 (.A(net2711),
    .X(net7125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6602 (.A(\rbzero.tex_g1[44] ),
    .X(net7126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6603 (.A(net2461),
    .X(net7127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6604 (.A(\rbzero.tex_g1[6] ),
    .X(net7128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6605 (.A(net2599),
    .X(net7129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6606 (.A(_04380_),
    .X(net7130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6607 (.A(net2600),
    .X(net7131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6608 (.A(\rbzero.tex_g1[23] ),
    .X(net7132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6609 (.A(net2765),
    .X(net7133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net5558),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6610 (.A(\rbzero.tex_b0[49] ),
    .X(net7134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6611 (.A(net2346),
    .X(net7135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6612 (.A(\rbzero.tex_b0[13] ),
    .X(net7136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6613 (.A(net2734),
    .X(net7137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6614 (.A(_04583_),
    .X(net7138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6615 (.A(net2735),
    .X(net7139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6616 (.A(\rbzero.tex_r1[34] ),
    .X(net7140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6617 (.A(net2568),
    .X(net7141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6618 (.A(\rbzero.tex_g0[45] ),
    .X(net7142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6619 (.A(net2538),
    .X(net7143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(net5560),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6620 (.A(\rbzero.tex_g1[5] ),
    .X(net7144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6621 (.A(net2325),
    .X(net7145));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold6622 (.A(net3194),
    .X(net7146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6623 (.A(_02715_),
    .X(net7147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6624 (.A(\rbzero.tex_r0[32] ),
    .X(net7148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6625 (.A(net2641),
    .X(net7149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6626 (.A(_04280_),
    .X(net7150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6627 (.A(net2642),
    .X(net7151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6628 (.A(\rbzero.tex_r1[53] ),
    .X(net7152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6629 (.A(net2363),
    .X(net7153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(net4860),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6630 (.A(_04183_),
    .X(net7154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6631 (.A(net2364),
    .X(net7155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6632 (.A(\rbzero.tex_g1[55] ),
    .X(net7156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6633 (.A(net2452),
    .X(net7157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6634 (.A(_04324_),
    .X(net7158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6635 (.A(net2497),
    .X(net7159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6636 (.A(\rbzero.tex_r1[54] ),
    .X(net7160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6637 (.A(net2571),
    .X(net7161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6638 (.A(\rbzero.tex_r0[36] ),
    .X(net7162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6639 (.A(net2644),
    .X(net7163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net4862),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6640 (.A(_04275_),
    .X(net7164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6641 (.A(net2645),
    .X(net7165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6642 (.A(\rbzero.tex_g1[59] ),
    .X(net7166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6643 (.A(net2625),
    .X(net7167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6644 (.A(\rbzero.tex_r1[15] ),
    .X(net7168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6645 (.A(net2728),
    .X(net7169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6646 (.A(_04224_),
    .X(net7170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6647 (.A(net2729),
    .X(net7171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6648 (.A(\rbzero.tex_r0[38] ),
    .X(net7172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6649 (.A(net2307),
    .X(net7173));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold665 (.A(net7881),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6650 (.A(\rbzero.tex_r1[31] ),
    .X(net7174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6651 (.A(net2635),
    .X(net7175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6652 (.A(\rbzero.tex_g1[60] ),
    .X(net7176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6653 (.A(net2781),
    .X(net7177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6654 (.A(\rbzero.tex_b0[44] ),
    .X(net7178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6655 (.A(net2316),
    .X(net7179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6656 (.A(\rbzero.tex_r1[52] ),
    .X(net7180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6657 (.A(net2602),
    .X(net7181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6658 (.A(\rbzero.tex_g1[27] ),
    .X(net7182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6659 (.A(net2490),
    .X(net7183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(net4272),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6660 (.A(\rbzero.tex_b0[16] ),
    .X(net7184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6661 (.A(net2816),
    .X(net7185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6662 (.A(\rbzero.tex_b1[11] ),
    .X(net7186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6663 (.A(net2784),
    .X(net7187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6664 (.A(_04516_),
    .X(net7188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6665 (.A(net2785),
    .X(net7189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6666 (.A(\rbzero.tex_r0[46] ),
    .X(net7190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6667 (.A(net2622),
    .X(net7191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6668 (.A(\rbzero.tex_r0[50] ),
    .X(net7192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6669 (.A(net2689),
    .X(net7193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net6448),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6670 (.A(\rbzero.spi_registers.buf_texadd1[15] ),
    .X(net7194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6671 (.A(net2487),
    .X(net7195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6672 (.A(\rbzero.tex_r1[18] ),
    .X(net7196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6673 (.A(net2731),
    .X(net7197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6674 (.A(_04221_),
    .X(net7198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6675 (.A(net2732),
    .X(net7199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6676 (.A(\rbzero.tex_b1[31] ),
    .X(net7200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6677 (.A(net2508),
    .X(net7201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6678 (.A(\rbzero.tex_r0[47] ),
    .X(net7202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6679 (.A(net2169),
    .X(net7203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(net6450),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6680 (.A(\rbzero.spi_registers.ss_buffer[0] ),
    .X(net7204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6681 (.A(net1211),
    .X(net7205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6682 (.A(\rbzero.tex_r0[40] ),
    .X(net7206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6683 (.A(net2759),
    .X(net7207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6684 (.A(\rbzero.tex_r1[25] ),
    .X(net7208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6685 (.A(net2484),
    .X(net7209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6686 (.A(\rbzero.tex_b0[19] ),
    .X(net7210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6687 (.A(net2656),
    .X(net7211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6688 (.A(\rbzero.tex_g1[37] ),
    .X(net7212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6689 (.A(net2737),
    .X(net7213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_01372_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6690 (.A(\rbzero.tex_b1[48] ),
    .X(net7214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6691 (.A(net2544),
    .X(net7215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6692 (.A(\rbzero.tex_g0[18] ),
    .X(net7216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6693 (.A(net2665),
    .X(net7217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6694 (.A(\rbzero.tex_b0[11] ),
    .X(net7218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6695 (.A(net2692),
    .X(net7219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6696 (.A(\rbzero.tex_r0[18] ),
    .X(net7220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6697 (.A(net2559),
    .X(net7221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6698 (.A(\rbzero.tex_b0[32] ),
    .X(net7222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6699 (.A(net2619),
    .X(net7223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net2093),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(net5535),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6700 (.A(\rbzero.tex_b1[40] ),
    .X(net7224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6701 (.A(net1923),
    .X(net7225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6702 (.A(\rbzero.tex_g1[39] ),
    .X(net7226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6703 (.A(net2674),
    .X(net7227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6704 (.A(\rbzero.tex_g1[51] ),
    .X(net7228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6705 (.A(net2632),
    .X(net7229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6706 (.A(_04329_),
    .X(net7230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6707 (.A(net2763),
    .X(net7231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6708 (.A(\rbzero.tex_r0[48] ),
    .X(net7232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6709 (.A(net2499),
    .X(net7233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(net5537),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6710 (.A(\rbzero.tex_r0[7] ),
    .X(net7234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6711 (.A(net2695),
    .X(net7235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6712 (.A(_04307_),
    .X(net7236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6713 (.A(net2696),
    .X(net7237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6714 (.A(\rbzero.tex_b1[53] ),
    .X(net7238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6715 (.A(net2743),
    .X(net7239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6716 (.A(\rbzero.tex_r1[27] ),
    .X(net7240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6717 (.A(net2556),
    .X(net7241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6718 (.A(\rbzero.tex_r0[55] ),
    .X(net7242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6719 (.A(net2418),
    .X(net7243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(net6428),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6720 (.A(\rbzero.tex_g0[48] ),
    .X(net7244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6721 (.A(net2662),
    .X(net7245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6722 (.A(\rbzero.tex_r0[6] ),
    .X(net7246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6723 (.A(net2682),
    .X(net7247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6724 (.A(\rbzero.tex_r1[2] ),
    .X(net7248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6725 (.A(net2723),
    .X(net7249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6726 (.A(\rbzero.tex_b1[21] ),
    .X(net7250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6727 (.A(net2796),
    .X(net7251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6728 (.A(\rbzero.tex_b1[15] ),
    .X(net7252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6729 (.A(net2866),
    .X(net7253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(net6430),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6730 (.A(\rbzero.tex_g0[19] ),
    .X(net7254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6731 (.A(net2717),
    .X(net7255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6732 (.A(\rbzero.debug_overlay.playerY[4] ),
    .X(net7256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6733 (.A(\rbzero.tex_b0[25] ),
    .X(net7257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6734 (.A(net2804),
    .X(net7258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6735 (.A(\rbzero.tex_g0[61] ),
    .X(net7259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6736 (.A(net2671),
    .X(net7260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6737 (.A(\rbzero.tex_r0[26] ),
    .X(net7261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6738 (.A(net2851),
    .X(net7262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6739 (.A(\rbzero.tex_b0[5] ),
    .X(net7263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_01149_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6740 (.A(net2793),
    .X(net7264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6741 (.A(\rbzero.tex_r1[17] ),
    .X(net7265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6742 (.A(net2702),
    .X(net7266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6743 (.A(\rbzero.tex_b1[10] ),
    .X(net7267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6744 (.A(net2858),
    .X(net7268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6745 (.A(\rbzero.tex_b0[52] ),
    .X(net7269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6746 (.A(net2799),
    .X(net7270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6747 (.A(\rbzero.tex_r1[55] ),
    .X(net7271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6748 (.A(net2750),
    .X(net7272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6749 (.A(\rbzero.tex_g0[21] ),
    .X(net7273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(net3678),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6750 (.A(net2740),
    .X(net7274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6751 (.A(\rbzero.tex_b0[12] ),
    .X(net7275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6752 (.A(net2809),
    .X(net7276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6753 (.A(\rbzero.tex_r1[1] ),
    .X(net7277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6754 (.A(net2753),
    .X(net7278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6755 (.A(\rbzero.tex_r1[19] ),
    .X(net7279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6756 (.A(net2827),
    .X(net7280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6757 (.A(\rbzero.tex_r0[56] ),
    .X(net7281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6758 (.A(net2756),
    .X(net7282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6759 (.A(\rbzero.tex_r0[31] ),
    .X(net7283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(net4857),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6760 (.A(net2668),
    .X(net7284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6761 (.A(\rbzero.tex_g1[11] ),
    .X(net7285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6762 (.A(net2876),
    .X(net7286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6763 (.A(\rbzero.tex_g1[41] ),
    .X(net7287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6764 (.A(net2830),
    .X(net7288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6765 (.A(\rbzero.tex_r0[35] ),
    .X(net7289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6766 (.A(net2845),
    .X(net7290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6767 (.A(\rbzero.tex_r0[51] ),
    .X(net7291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6768 (.A(net2848),
    .X(net7292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6769 (.A(\rbzero.tex_b0[55] ),
    .X(net7293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(net6414),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6770 (.A(net2613),
    .X(net7294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6771 (.A(\rbzero.tex_g0[54] ),
    .X(net7295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6772 (.A(net2897),
    .X(net7296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6773 (.A(\rbzero.tex_b1[12] ),
    .X(net7297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6774 (.A(net2881),
    .X(net7298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6775 (.A(\rbzero.tex_r0[4] ),
    .X(net7299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6776 (.A(net2714),
    .X(net7300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6777 (.A(\rbzero.tex_g0[38] ),
    .X(net7301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6778 (.A(net2870),
    .X(net7302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6779 (.A(\rbzero.tex_g1[57] ),
    .X(net7303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(net6416),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6780 (.A(net2861),
    .X(net7304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6781 (.A(_04323_),
    .X(net7305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6782 (.A(net2862),
    .X(net7306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6783 (.A(\gpout0.vpos[2] ),
    .X(net7307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6784 (.A(\rbzero.tex_r0[27] ),
    .X(net7308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6785 (.A(net2902),
    .X(net7309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6786 (.A(\rbzero.pov.ready_buffer[69] ),
    .X(net7310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6787 (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .X(net7311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6788 (.A(_03304_),
    .X(net7312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6789 (.A(_00840_),
    .X(net7313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_01412_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6790 (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .X(net7314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6791 (.A(_02496_),
    .X(net7315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6792 (.A(_00841_),
    .X(net7316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6793 (.A(\rbzero.wall_hot[1] ),
    .X(net7317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6794 (.A(_04638_),
    .X(net7318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6795 (.A(_09945_),
    .X(net7319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6797 (.A(_02931_),
    .X(net7321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6798 (.A(net7363),
    .X(net7322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6799 (.A(_03089_),
    .X(net7323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_03193_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(net5550),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6800 (.A(\rbzero.pov.spi_counter[3] ),
    .X(net7324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6801 (.A(\rbzero.color_floor[1] ),
    .X(net7325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6802 (.A(_03097_),
    .X(net7326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6803 (.A(net7365),
    .X(net7327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6804 (.A(_03100_),
    .X(net7328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6805 (.A(\rbzero.pov.spi_counter[5] ),
    .X(net7329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6806 (.A(_03671_),
    .X(net7330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6807 (.A(_03672_),
    .X(net7331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6809 (.A(_03607_),
    .X(net7333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(net5552),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6811 (.A(_03611_),
    .X(net7335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6813 (.A(_03603_),
    .X(net7337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6814 (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .X(net7338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6815 (.A(_00865_),
    .X(net7339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6817 (.A(_03605_),
    .X(net7341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6819 (.A(_03599_),
    .X(net7343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(net6432),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6821 (.A(_03589_),
    .X(net7345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6822 (.A(\rbzero.debug_overlay.playerX[4] ),
    .X(net7346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6823 (.A(\rbzero.pov.spi_counter[4] ),
    .X(net7347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6825 (.A(_03587_),
    .X(net7349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6827 (.A(_03591_),
    .X(net7351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6828 (.A(\gpout0.hpos[4] ),
    .X(net7352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6829 (.A(\rbzero.trace_state[3] ),
    .X(net7353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(net6434),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6830 (.A(\rbzero.spi_registers.spi_counter[1] ),
    .X(net7354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6831 (.A(_02970_),
    .X(net7355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6832 (.A(\rbzero.spi_registers.spi_counter[3] ),
    .X(net7356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6833 (.A(_02976_),
    .X(net7357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6834 (.A(\rbzero.spi_registers.spi_counter[4] ),
    .X(net7358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6835 (.A(\rbzero.spi_registers.spi_counter[0] ),
    .X(net7359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6836 (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .X(net7360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6837 (.A(\gpout0.hpos[8] ),
    .X(net7361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6838 (.A(_04815_),
    .X(net7362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6839 (.A(\rbzero.color_sky[2] ),
    .X(net7363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_01422_),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6840 (.A(\gpout0.hpos[5] ),
    .X(net7364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6841 (.A(\rbzero.color_floor[3] ),
    .X(net7365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6842 (.A(\rbzero.spi_registers.buf_sky[4] ),
    .X(net7366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6843 (.A(net7725),
    .X(net7367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6844 (.A(net2985),
    .X(net7368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6845 (.A(\rbzero.debug_overlay.playerX[-9] ),
    .X(net7369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6846 (.A(net4335),
    .X(net7370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6847 (.A(_09287_),
    .X(net7371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6848 (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .X(net7372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6849 (.A(net3272),
    .X(net7373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(net4832),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6850 (.A(_10574_),
    .X(net7374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6851 (.A(_10576_),
    .X(net7375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6852 (.A(_10578_),
    .X(net7376));
 sky130_fd_sc_hd__clkbuf_1 hold6853 (.A(net4827),
    .X(net7377));
 sky130_fd_sc_hd__clkbuf_4 hold6854 (.A(_09790_),
    .X(net7378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6855 (.A(\rbzero.debug_overlay.playerY[-5] ),
    .X(net7379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6856 (.A(net4294),
    .X(net7380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6857 (.A(_09404_),
    .X(net7381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(net4834),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net7204),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6877 (.A(_08337_),
    .X(net7401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6878 (.A(_08338_),
    .X(net7402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6879 (.A(_08339_),
    .X(net7403));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold688 (.A(_02490_),
    .X(net1212));
 sky130_fd_sc_hd__buf_1 hold6880 (.A(_08341_),
    .X(net7404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6881 (.A(_08381_),
    .X(net7405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6882 (.A(_09296_),
    .X(net7406));
 sky130_fd_sc_hd__buf_2 hold6883 (.A(_09297_),
    .X(net7407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6884 (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .X(net7408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_00573_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net4262),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(net5717),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6903 (.A(\rbzero.debug_overlay.playerX[-4] ),
    .X(net7427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6904 (.A(net4300),
    .X(net7428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6906 (.A(_08170_),
    .X(net7430));
 sky130_fd_sc_hd__clkbuf_2 hold6907 (.A(_06712_),
    .X(net7431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6908 (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .X(net7432));
 sky130_fd_sc_hd__buf_2 hold6909 (.A(_06733_),
    .X(net7433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_03196_),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_2 hold6910 (.A(net7912),
    .X(net7434));
 sky130_fd_sc_hd__buf_1 hold6912 (.A(_06765_),
    .X(net7436));
 sky130_fd_sc_hd__buf_1 hold6913 (.A(_08130_),
    .X(net7437));
 sky130_fd_sc_hd__buf_2 hold6914 (.A(_07311_),
    .X(net7438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6915 (.A(_08119_),
    .X(net7439));
 sky130_fd_sc_hd__clkbuf_4 hold6916 (.A(net4779),
    .X(net7440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6917 (.A(_09665_),
    .X(net7441));
 sky130_fd_sc_hd__clkbuf_4 hold6918 (.A(net6134),
    .X(net7442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(net4209),
    .X(net1216));
 sky130_fd_sc_hd__clkbuf_4 hold6920 (.A(net7945),
    .X(net7444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6921 (.A(\rbzero.debug_overlay.playerY[-2] ),
    .X(net7445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6922 (.A(net4358),
    .X(net7446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6923 (.A(_09770_),
    .X(net7447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6924 (.A(\rbzero.traced_texVinit[8] ),
    .X(net7448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6925 (.A(net4184),
    .X(net7449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6926 (.A(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(net7450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6927 (.A(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(net7451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6929 (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .X(net7453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(net5791),
    .X(net1217));
 sky130_fd_sc_hd__clkbuf_2 hold6933 (.A(net7568),
    .X(net7457));
 sky130_fd_sc_hd__clkbuf_2 hold6934 (.A(_06800_),
    .X(net7458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6935 (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .X(net7459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6936 (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .X(net7460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_03184_),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6940 (.A(net7923),
    .X(net7464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6943 (.A(\rbzero.wall_tracer.stepDistY[-3] ),
    .X(net7467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6944 (.A(net3504),
    .X(net7468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6947 (.A(\rbzero.traced_texVinit[7] ),
    .X(net7471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6948 (.A(net4141),
    .X(net7472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(net4212),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6951 (.A(\rbzero.wall_tracer.stepDistX[-3] ),
    .X(net7475));
 sky130_fd_sc_hd__clkbuf_4 hold6952 (.A(net4581),
    .X(net7476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6953 (.A(_08329_),
    .X(net7477));
 sky130_fd_sc_hd__buf_1 hold6954 (.A(_06721_),
    .X(net7478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6955 (.A(\rbzero.wall_tracer.stepDistX[2] ),
    .X(net7479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6956 (.A(net4348),
    .X(net7480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6957 (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .X(net7481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6958 (.A(\rbzero.traced_texVinit[0] ),
    .X(net7482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6959 (.A(net4110),
    .X(net7483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(net3382),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6962 (.A(\rbzero.traced_texVinit[2] ),
    .X(net7486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6963 (.A(net4158),
    .X(net7487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6964 (.A(\rbzero.wall_tracer.stepDistY[1] ),
    .X(net7488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6965 (.A(net4371),
    .X(net7489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6966 (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .X(net7490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6967 (.A(\rbzero.traced_texVinit[6] ),
    .X(net7491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6968 (.A(net4139),
    .X(net7492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6969 (.A(\rbzero.wall_tracer.stepDistX[1] ),
    .X(net7493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(net4885),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6970 (.A(net4410),
    .X(net7494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6973 (.A(\rbzero.traced_texVinit[3] ),
    .X(net7497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6974 (.A(net4182),
    .X(net7498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6975 (.A(\rbzero.traced_texVinit[5] ),
    .X(net7499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6976 (.A(net4165),
    .X(net7500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6977 (.A(\rbzero.traced_texVinit[4] ),
    .X(net7501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6978 (.A(net4163),
    .X(net7502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(net5409),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6982 (.A(_00502_),
    .X(net7506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6983 (.A(net4203),
    .X(net7507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6986 (.A(_08348_),
    .X(net7510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6987 (.A(_08349_),
    .X(net7511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6989 (.A(_00500_),
    .X(net7513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(net5411),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6990 (.A(net4233),
    .X(net7514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6992 (.A(_00499_),
    .X(net7516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6993 (.A(net4252),
    .X(net7517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6995 (.A(_00501_),
    .X(net7519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6996 (.A(net4298),
    .X(net7520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6997 (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .X(net7521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6998 (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .X(net7522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6999 (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(net7523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net1562),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(net3683),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7000 (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .X(net7524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7001 (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .X(net7525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7002 (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .X(net7526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7003 (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .X(net7527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7004 (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .X(net7528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7005 (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(net7529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7006 (.A(net4488),
    .X(net7530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7007 (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .X(net7531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7008 (.A(net4486),
    .X(net7532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7009 (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .X(net7533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(net5531),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7010 (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .X(net7534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7011 (.A(net4484),
    .X(net7535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7012 (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .X(net7536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7013 (.A(\rbzero.traced_texa[9] ),
    .X(net7537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7014 (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .X(net7538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7015 (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(net7539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7016 (.A(net4510),
    .X(net7540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7017 (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .X(net7541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7018 (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .X(net7542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7019 (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .X(net7543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(net3351),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7020 (.A(net4490),
    .X(net7544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7021 (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .X(net7545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7022 (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .X(net7546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7023 (.A(net4594),
    .X(net7547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7024 (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .X(net7548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7025 (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .X(net7549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7026 (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .X(net7550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7027 (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .X(net7551));
 sky130_fd_sc_hd__clkbuf_4 hold7028 (.A(net4783),
    .X(net7552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7029 (.A(_00511_),
    .X(net7553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(net4589),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_2 hold7030 (.A(net7377),
    .X(net7554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7031 (.A(_00520_),
    .X(net7555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7033 (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .X(net7557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7034 (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .X(net7558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7036 (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .X(net7560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7037 (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(net7561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7038 (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .X(net7562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(net5211),
    .X(net1228));
 sky130_fd_sc_hd__clkbuf_4 hold7042 (.A(_06660_),
    .X(net7566));
 sky130_fd_sc_hd__buf_1 hold7044 (.A(_06788_),
    .X(net7568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7045 (.A(\rbzero.traced_texa[2] ),
    .X(net7569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7047 (.A(_02673_),
    .X(net7571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7048 (.A(_02675_),
    .X(net7572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7049 (.A(\rbzero.traced_texa[8] ),
    .X(net7573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(net5213),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7051 (.A(_02798_),
    .X(net7575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7052 (.A(_02800_),
    .X(net7576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7053 (.A(_00603_),
    .X(net7577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7056 (.A(_02890_),
    .X(net7580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7057 (.A(_02891_),
    .X(net7581));
 sky130_fd_sc_hd__buf_4 hold7058 (.A(net4732),
    .X(net7582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7059 (.A(_00001_),
    .X(net7583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(net3659),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7061 (.A(_02581_),
    .X(net7585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7062 (.A(_02583_),
    .X(net7586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7065 (.A(_08321_),
    .X(net7589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7066 (.A(_08322_),
    .X(net7590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(net5601),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7070 (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .X(net7594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7071 (.A(net4398),
    .X(net7595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7072 (.A(_10054_),
    .X(net7596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7074 (.A(_02878_),
    .X(net7598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7075 (.A(_02883_),
    .X(net7599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7077 (.A(_02602_),
    .X(net7601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7078 (.A(_02605_),
    .X(net7602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(net5250),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7082 (.A(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(net7606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7084 (.A(_02661_),
    .X(net7608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7085 (.A(_02666_),
    .X(net7609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7087 (.A(_02819_),
    .X(net7611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7088 (.A(_02822_),
    .X(net7612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7089 (.A(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(net7613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(net5252),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7090 (.A(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(net7614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7091 (.A(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(net7615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7092 (.A(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(net7616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7093 (.A(\rbzero.spi_registers.texadd1[16] ),
    .X(net7617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7095 (.A(_00506_),
    .X(net7619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7096 (.A(\rbzero.spi_registers.buf_texadd0[13] ),
    .X(net7620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7097 (.A(\rbzero.pov.ready_buffer[36] ),
    .X(net7621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7098 (.A(\rbzero.spi_registers.texadd3[11] ),
    .X(net7622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7099 (.A(\rbzero.spi_registers.texadd0[11] ),
    .X(net7623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_03195_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(net6420),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7100 (.A(\rbzero.spi_registers.texadd3[12] ),
    .X(net7624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7101 (.A(\rbzero.spi_registers.texadd0[14] ),
    .X(net7625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7103 (.A(_02843_),
    .X(net7627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7104 (.A(\rbzero.spi_registers.texadd1[10] ),
    .X(net7628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7105 (.A(\rbzero.wall_tracer.rayAddendY[-6] ),
    .X(net7629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7107 (.A(_02626_),
    .X(net7631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7108 (.A(\rbzero.pov.ready_buffer[2] ),
    .X(net7632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7109 (.A(\rbzero.traced_texa[-2] ),
    .X(net7633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(net6422),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7110 (.A(\rbzero.spi_registers.texadd0[12] ),
    .X(net7634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7111 (.A(\rbzero.traced_texa[-3] ),
    .X(net7635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7112 (.A(\rbzero.spi_registers.texadd2[19] ),
    .X(net7636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7113 (.A(\rbzero.traced_texa[5] ),
    .X(net7637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7114 (.A(\rbzero.pov.ready_buffer[28] ),
    .X(net7638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7115 (.A(\rbzero.wall_tracer.rayAddendX[-5] ),
    .X(net7639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7116 (.A(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(net7640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7117 (.A(\rbzero.traced_texa[-1] ),
    .X(net7641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7118 (.A(\rbzero.traced_texa[7] ),
    .X(net7642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7119 (.A(\rbzero.traced_texa[6] ),
    .X(net7643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_01302_),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7120 (.A(\rbzero.traced_texa[0] ),
    .X(net7644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7121 (.A(\rbzero.pov.ready_buffer[27] ),
    .X(net7645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7122 (.A(\rbzero.spi_registers.texadd2[0] ),
    .X(net7646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7123 (.A(\rbzero.pov.ready_buffer[35] ),
    .X(net7647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7124 (.A(\rbzero.traced_texa[4] ),
    .X(net7648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7125 (.A(\rbzero.spi_registers.texadd2[23] ),
    .X(net7649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7126 (.A(\rbzero.wall_tracer.mapY[6] ),
    .X(net7650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7127 (.A(\rbzero.floor_leak[1] ),
    .X(net7651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7128 (.A(\rbzero.pov.ready_buffer[13] ),
    .X(net7652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7129 (.A(\rbzero.wall_tracer.mapX[6] ),
    .X(net7653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(net3640),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7130 (.A(\rbzero.spi_registers.texadd2[16] ),
    .X(net7654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7131 (.A(\rbzero.texV[3] ),
    .X(net7655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7132 (.A(\rbzero.spi_registers.texadd2[15] ),
    .X(net7656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7133 (.A(\rbzero.spi_registers.texadd2[6] ),
    .X(net7657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7134 (.A(\rbzero.spi_registers.buf_texadd2[20] ),
    .X(net7658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7135 (.A(\rbzero.spi_registers.buf_texadd3[10] ),
    .X(net7659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7136 (.A(\rbzero.spi_registers.texadd2[12] ),
    .X(net7660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7137 (.A(\rbzero.spi_registers.buf_texadd3[7] ),
    .X(net7661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7138 (.A(\rbzero.row_render.texu[4] ),
    .X(net7662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7139 (.A(\rbzero.spi_registers.texadd2[11] ),
    .X(net7663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(net5573),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7140 (.A(\rbzero.spi_registers.buf_texadd1[17] ),
    .X(net7664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7141 (.A(\rbzero.spi_registers.buf_texadd3[8] ),
    .X(net7665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7142 (.A(\rbzero.spi_registers.buf_texadd3[23] ),
    .X(net7666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7143 (.A(\rbzero.spi_registers.buf_texadd1[19] ),
    .X(net7667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7144 (.A(\rbzero.spi_registers.texadd2[13] ),
    .X(net7668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7145 (.A(\rbzero.spi_registers.buf_texadd2[10] ),
    .X(net7669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7146 (.A(\rbzero.row_render.texu[3] ),
    .X(net7670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7147 (.A(\rbzero.row_render.texu[1] ),
    .X(net7671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7148 (.A(\rbzero.spi_registers.buf_leak[0] ),
    .X(net7672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7149 (.A(\rbzero.spi_registers.texadd3[14] ),
    .X(net7673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(net3274),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7150 (.A(\rbzero.spi_registers.buf_sky[5] ),
    .X(net7674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7151 (.A(\rbzero.spi_registers.texadd2[14] ),
    .X(net7675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7152 (.A(\rbzero.traced_texa[-11] ),
    .X(net7676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7153 (.A(\rbzero.row_render.texu[2] ),
    .X(net7677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7154 (.A(\rbzero.pov.ready_buffer[30] ),
    .X(net7678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7155 (.A(\rbzero.row_render.texu[0] ),
    .X(net7679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(net5450),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(net3669),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net4846),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7187 (.A(\rbzero.traced_texVinit[1] ),
    .X(net7711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7188 (.A(net4189),
    .X(net7712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(net3736),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7193 (.A(\rbzero.traced_texVinit[9] ),
    .X(net7717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7194 (.A(net4200),
    .X(net7718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7197 (.A(\rbzero.traced_texVinit[10] ),
    .X(net7721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7198 (.A(net4230),
    .X(net7722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7199 (.A(\rbzero.row_render.size[5] ),
    .X(net7723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net4292),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(net5508),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7200 (.A(net4283),
    .X(net7724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7201 (.A(\rbzero.texu_hot[5] ),
    .X(net7725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7202 (.A(net7367),
    .X(net7726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7207 (.A(\rbzero.debug_overlay.playerX[-6] ),
    .X(net7731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7208 (.A(net4338),
    .X(net7732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7209 (.A(_09277_),
    .X(net7733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(net5208),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7211 (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .X(net7735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7212 (.A(net4341),
    .X(net7736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7213 (.A(\rbzero.texu_hot[3] ),
    .X(net7737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7214 (.A(net4383),
    .X(net7738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7215 (.A(\rbzero.texu_hot[2] ),
    .X(net7739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7216 (.A(net4312),
    .X(net7740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7217 (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .X(net7741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7218 (.A(net4432),
    .X(net7742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7219 (.A(\rbzero.wall_tracer.stepDistY[2] ),
    .X(net7743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(net5210),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7220 (.A(net4422),
    .X(net7744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7223 (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .X(net7747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7224 (.A(\rbzero.row_render.size[6] ),
    .X(net7748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7226 (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .X(net7750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7227 (.A(net4576),
    .X(net7751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7228 (.A(\rbzero.debug_overlay.playerX[-8] ),
    .X(net7752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7229 (.A(\rbzero.texu_hot[4] ),
    .X(net7753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(net3487),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7230 (.A(net4518),
    .X(net7754));
 sky130_fd_sc_hd__buf_4 hold7233 (.A(_06611_),
    .X(net7757));
 sky130_fd_sc_hd__clkbuf_2 hold7235 (.A(_06725_),
    .X(net7759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7237 (.A(_08335_),
    .X(net7761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7238 (.A(\rbzero.wall_tracer.stepDistX[-11] ),
    .X(net7762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(net5771),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7240 (.A(_08487_),
    .X(net7764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7242 (.A(_08427_),
    .X(net7766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7243 (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .X(net7767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7245 (.A(_08600_),
    .X(net7769));
 sky130_fd_sc_hd__buf_2 hold7246 (.A(net7554),
    .X(net7770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7247 (.A(_06717_),
    .X(net7771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7249 (.A(_08451_),
    .X(net7773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net4921),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7251 (.A(_08406_),
    .X(net7775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7253 (.A(_08389_),
    .X(net7777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7255 (.A(_08360_),
    .X(net7779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7256 (.A(\rbzero.wall_tracer.stepDistY[-7] ),
    .X(net7780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7257 (.A(net4381),
    .X(net7781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7258 (.A(_02364_),
    .X(net7782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(net4923),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7263 (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .X(net7787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7264 (.A(net4385),
    .X(net7788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7265 (.A(_02463_),
    .X(net7789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7266 (.A(_02464_),
    .X(net7790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7267 (.A(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(net7791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7268 (.A(net4314),
    .X(net7792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7269 (.A(_02343_),
    .X(net7793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(net3322),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7270 (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .X(net7794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7271 (.A(net4369),
    .X(net7795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7272 (.A(_10027_),
    .X(net7796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7273 (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .X(net7797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7274 (.A(_01977_),
    .X(net7798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7275 (.A(_01978_),
    .X(net7799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7276 (.A(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(net7800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7277 (.A(_02390_),
    .X(net7801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(net4465),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7280 (.A(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(net7804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7281 (.A(_02350_),
    .X(net7805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7282 (.A(\rbzero.wall_tracer.stepDistY[0] ),
    .X(net7806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7283 (.A(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(net7807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7285 (.A(_08368_),
    .X(net7809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7286 (.A(_08369_),
    .X(net7810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7287 (.A(\rbzero.wall_tracer.stepDistX[3] ),
    .X(net7811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7288 (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .X(net7812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7289 (.A(net4377),
    .X(net7813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(net3704),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7290 (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .X(net7814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7291 (.A(_02077_),
    .X(net7815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7292 (.A(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(net7816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7293 (.A(net4373),
    .X(net7817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7294 (.A(_02379_),
    .X(net7818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7295 (.A(\rbzero.wall_tracer.stepDistY[-5] ),
    .X(net7819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7296 (.A(net4472),
    .X(net7820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7298 (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .X(net7822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7299 (.A(net4333),
    .X(net7823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net2013),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(net4852),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7300 (.A(_10086_),
    .X(net7824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7301 (.A(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(net7825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7302 (.A(net4434),
    .X(net7826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7303 (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(net7827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7304 (.A(net4361),
    .X(net7828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7309 (.A(\rbzero.wall_tracer.stepDistY[4] ),
    .X(net7833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(net5604),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7310 (.A(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(net7834));
 sky130_fd_sc_hd__clkbuf_2 hold7312 (.A(_06716_),
    .X(net7836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7314 (.A(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(net7838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7315 (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(net7839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7316 (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(net7840));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7319 (.A(_06663_),
    .X(net7843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(net5606),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7320 (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(net7844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7321 (.A(\rbzero.row_render.size[3] ),
    .X(net7845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7322 (.A(\rbzero.row_render.size[0] ),
    .X(net7846));
 sky130_fd_sc_hd__buf_1 hold733 (.A(net7718),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(net6436),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(net6438),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7356 (.A(\rbzero.texu_hot[1] ),
    .X(net7880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7357 (.A(net4350),
    .X(net7881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_01472_),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7362 (.A(_08046_),
    .X(net7886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7363 (.A(\rbzero.row_render.size[9] ),
    .X(net7887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7364 (.A(net4508),
    .X(net7888));
 sky130_fd_sc_hd__clkbuf_2 hold7367 (.A(_06838_),
    .X(net7891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7368 (.A(\rbzero.wall_tracer.stepDistY[8] ),
    .X(net7892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(net5577),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7375 (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .X(net7899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7376 (.A(\rbzero.texu_hot[0] ),
    .X(net7900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7377 (.A(net4375),
    .X(net7901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7378 (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .X(net7902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(net5579),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7380 (.A(\rbzero.debug_overlay.playerX[-5] ),
    .X(net7904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7382 (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .X(net7906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7383 (.A(net4331),
    .X(net7907));
 sky130_fd_sc_hd__buf_2 hold7384 (.A(_06689_),
    .X(net7908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7388 (.A(_06722_),
    .X(net7912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(net5519),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7390 (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .X(net7914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7391 (.A(\rbzero.wall_tracer.stepDistY[5] ),
    .X(net7915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7392 (.A(net4367),
    .X(net7916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7394 (.A(\rbzero.wall_tracer.stepDistY[7] ),
    .X(net7918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7399 (.A(_08301_),
    .X(net7923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_03222_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(net5521),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7400 (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .X(net7924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(net5587),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7415 (.A(net656),
    .X(net7939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7418 (.A(\rbzero.row_render.size[2] ),
    .X(net7942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(net5589),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7421 (.A(_08623_),
    .X(net7945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7427 (.A(net6146),
    .X(net7951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(net6440),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(net6442),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(_01322_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(net5239),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(net5241),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7475 (.A(\rbzero.debug_overlay.playerY[-9] ),
    .X(net7999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(net3290),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7485 (.A(\rbzero.debug_overlay.playerX[-7] ),
    .X(net8009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7486 (.A(_09282_),
    .X(net8010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(net5603),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7492 (.A(_06158_),
    .X(net8016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7493 (.A(net7440),
    .X(net8017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net4119),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(net5048),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(net5050),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(net5581),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(net5583),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(net5113),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(net5115),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(net5590),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(net5592),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(net4849),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_01097_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net1988),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(net5382),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7602 (.A(_06146_),
    .X(net8126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(net5384),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(net5553),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(net5555),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(net5516),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(net5518),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(net5192),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(net5194),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net5543),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(net5545),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_03223_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(net5539),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(net5541),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(net5618),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(net5620),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(net7652),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(net4448),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(net5628),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(net5630),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(net4880),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(net4882),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net4113),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(net7740),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(net4304),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(net3799),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(net5637),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(net5593),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(net5595),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(net5608),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(net5610),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(net5677),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(net5679),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net5120),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(net3411),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(net5688),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(net3567),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(_01093_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(net5386),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(net5388),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(net5648),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(net5650),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(net3645),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(_01092_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_03127_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(net5218),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(net5220),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(net5655),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(net5657),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(net3816),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(net5557),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(net5651),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(net5653),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(net6456),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(net6458),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net4122),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_01358_),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(net5480),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(net5485),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(net5622),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(net5624),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(net3842),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(net5569),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(net5625),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(net5627),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(net3341),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net5349),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(net5433),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(net5641),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(net5643),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(net6444),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(net6446),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(_01532_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(net5668),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(net5670),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(net6464),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(net6466),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_03131_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_01502_),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(net3751),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(net4841),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(net6460),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(net6462),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(_01115_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(net3513),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_01104_),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(net3597),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_01091_),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net4128),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(net4700),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(net4702),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(net3448),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(net4774),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(net5632),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(net5634),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(net3664),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(net5672),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(net6424),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(net6426),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net968),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_01311_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(net5204),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(net5206),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(net5613),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(net5615),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(net5680),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(net5682),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(net3781),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(net5176),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(net6503),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_03129_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_04499_),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_01292_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(net6468),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(net6470),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_01155_),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(net5574),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(net5576),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(net5659),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(net5661),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(net7738),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net4150),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(net4281),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(net3434),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(net5694),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(net6492),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(net6494),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(_01298_),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(net5664),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(net5666),
    .X(net1401));
 sky130_fd_sc_hd__buf_1 hold878 (.A(net5701),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(net5703),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net3021),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(net5673),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(net5675),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(net1783),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(_03197_),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(net4206),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(net3556),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(net5483),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(net3495),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_01105_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(net3529),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net4237),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_01075_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(net5689),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(net5691),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(net6476),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(net6478),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(_01139_),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(net5638),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(net5640),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(net7901),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(net4240),
    .X(net1423));
 sky130_fd_sc_hd__buf_2 hold90 (.A(net5837),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(net6488),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(net6490),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_01507_),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(net6511),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(net6513),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(_01418_),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net6530),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(net6532),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_01468_),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(net5232),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net4259),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(net5234),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(net6538),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(net6540),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(_01288_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(net3650),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(_01064_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(net5695),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(net5697),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(net6507),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(net6509),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net3037),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_01135_),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(net6484),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(net6486),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(_01392_),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(net6519),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(net6521),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_01538_),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(net4102),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(net6267),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(net6452),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net5797),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(net6454),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(_01523_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(net4541),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(net4543),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(net7088),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(net5858),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_01527_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(net6505),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_04532_),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(_01169_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net3010),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(net6515),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(net6517),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_01582_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(net6306),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_02991_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(_00628_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(net5174),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(net5495),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(net2100),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(_04250_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_03158_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_01517_),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(net5645),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(net5647),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(net6499),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(net6501),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(_01477_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(net6472),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(net6474),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_01267_),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(net3811),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net4125),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(net4848),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(net6593),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(net6595),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(_01321_),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\rbzero.tex_r0[0] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(net5776),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_01459_),
    .X(net1490));
 sky130_fd_sc_hd__buf_1 hold967 (.A(net5438),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(net5440),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(net5431),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net6323),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(net5445),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(net7754),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(net4255),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(net6534),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(net6536),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(_01144_),
    .X(net1499));
 sky130_fd_sc_hd__buf_1 hold976 (.A(net7722),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(net6480),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(net6482),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(_01395_),
    .X(net1503));
 sky130_fd_sc_hd__buf_1 hold98 (.A(_03028_),
    .X(net622));
 sky130_fd_sc_hd__buf_1 hold980 (.A(net4652),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(net4654),
    .X(net1505));
 sky130_fd_sc_hd__buf_1 hold982 (.A(net5732),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(net5734),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(net4867),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(net4869),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(net5532),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(net5534),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(net6550),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(net6552),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_00653_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_01429_),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(net6526),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(net6528),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(_01406_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(net6546),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(_04460_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_01328_),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\rbzero.tex_b0[0] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(net5768),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(_01110_),
    .X(net1523));
 sky130_fd_sc_hd__buf_2 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(i_gpout1_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(i_gpout1_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(i_gpout1_sel[2]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(i_gpout1_sel[3]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(i_gpout1_sel[4]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(i_gpout1_sel[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(i_gpout2_sel[0]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(i_gpout2_sel[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(i_gpout2_sel[2]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(i_gpout2_sel[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(i_debug_trace_overlay),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(i_gpout2_sel[4]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(i_gpout2_sel[5]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(i_gpout3_sel[0]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(i_gpout3_sel[1]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(i_gpout3_sel[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(i_gpout3_sel[3]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(i_gpout3_sel[4]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(i_gpout3_sel[5]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(i_gpout4_sel[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(i_gpout4_sel[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(i_debug_vec_overlay),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(i_gpout4_sel[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(i_gpout4_sel[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(i_gpout4_sel[4]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(i_gpout4_sel[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(i_gpout5_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(i_gpout5_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(i_gpout5_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(i_gpout5_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(i_gpout5_sel[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(i_gpout5_sel[5]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(i_gpout0_sel[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_8 input40 (.A(i_mode[0]),
    .X(net40));
 sky130_fd_sc_hd__buf_6 input41 (.A(i_mode[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(i_mode[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_4 input43 (.A(i_reg_csb),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(i_reg_mosi),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(i_reg_outs_enb),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(i_reg_sclk),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(i_reset_lock_a),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_reset_lock_b),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(i_test_uc2),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(i_gpout0_sel[1]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(i_test_wci),
    .X(net50));
 sky130_fd_sc_hd__buf_8 input51 (.A(i_tex_in[0]),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(i_tex_in[1]),
    .X(net52));
 sky130_fd_sc_hd__buf_8 input53 (.A(i_tex_in[2]),
    .X(net53));
 sky130_fd_sc_hd__buf_8 input54 (.A(i_tex_in[3]),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(i_vec_csb),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(i_vec_mosi),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input57 (.A(i_vec_sclk),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input6 (.A(i_gpout0_sel[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(i_gpout0_sel[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(i_gpout0_sel[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(i_gpout0_sel[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 max_cap77 (.A(_09366_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 max_cap78 (.A(_07878_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 max_cap82 (.A(_06481_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 max_cap83 (.A(_04816_),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap84 (.A(_06429_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 max_cap87 (.A(_02609_),
    .X(net87));
 sky130_fd_sc_hd__buf_4 max_cap89 (.A(_04167_),
    .X(net89));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_1_1__leaf__04800_),
    .Y(net141));
 sky130_fd_sc_hd__buf_1 output58 (.A(net58),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__buf_1 output59 (.A(net59),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__buf_1 output60 (.A(net60),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__buf_1 output61 (.A(net61),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__buf_1 output62 (.A(net62),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__buf_1 output63 (.A(net63),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(o_hsync));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(o_reset));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(o_tex_csb));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(o_tex_out0));
 sky130_fd_sc_hd__buf_1 output75 (.A(net140),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(o_vsync));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(net526),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(net533),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 rebuffer11 (.A(_07103_),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_2 rebuffer12 (.A(net3203),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(_07141_),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_1 rebuffer14 (.A(_06530_),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(net538),
    .X(net539));
 sky130_fd_sc_hd__buf_6 rebuffer16 (.A(net3132),
    .X(net540));
 sky130_fd_sc_hd__buf_1 rebuffer17 (.A(_06896_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net541),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 rebuffer19 (.A(net542),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(_07110_),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_1 rebuffer20 (.A(net543),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(net542),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(_06896_),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(net546),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 rebuffer25 (.A(_07112_),
    .X(net549));
 sky130_fd_sc_hd__buf_1 rebuffer26 (.A(_07109_),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_1 rebuffer27 (.A(_07137_),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(_06819_),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_1 rebuffer29 (.A(net562),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 rebuffer3 (.A(_07963_),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(net553),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_1 rebuffer31 (.A(_07104_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(_06827_),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 rebuffer33 (.A(net556),
    .X(net557));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer34 (.A(_07058_),
    .X(net1998));
 sky130_fd_sc_hd__clkbuf_2 rebuffer35 (.A(_07231_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_2 rebuffer36 (.A(_07249_),
    .X(net560));
 sky130_fd_sc_hd__buf_1 rebuffer37 (.A(_06781_),
    .X(net561));
 sky130_fd_sc_hd__buf_6 rebuffer38 (.A(_06819_),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 rebuffer39 (.A(net562),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(_07156_),
    .X(net528));
 sky130_fd_sc_hd__buf_1 rebuffer40 (.A(_06973_),
    .X(net564));
 sky130_fd_sc_hd__buf_1 rebuffer41 (.A(_06942_),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_1 rebuffer42 (.A(_07062_),
    .X(net566));
 sky130_fd_sc_hd__buf_1 rebuffer43 (.A(_06857_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd2_1 rebuffer44 (.A(net567),
    .X(net568));
 sky130_fd_sc_hd__buf_1 rebuffer45 (.A(net568),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_1 rebuffer46 (.A(_07035_),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_1 rebuffer47 (.A(_07076_),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_1 rebuffer48 (.A(_06893_),
    .X(net572));
 sky130_fd_sc_hd__buf_1 rebuffer49 (.A(_06858_),
    .X(net573));
 sky130_fd_sc_hd__buf_1 rebuffer5 (.A(_06966_),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 rebuffer50 (.A(_07078_),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 rebuffer51 (.A(_06909_),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 rebuffer52 (.A(_06901_),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 rebuffer53 (.A(_06900_),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 rebuffer54 (.A(_06882_),
    .X(net578));
 sky130_fd_sc_hd__buf_6 rebuffer55 (.A(_06882_),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 rebuffer56 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 rebuffer57 (.A(net584),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 rebuffer58 (.A(_06780_),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_1 rebuffer59 (.A(_07106_),
    .X(net583));
 sky130_fd_sc_hd__buf_1 rebuffer6 (.A(net529),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_1 rebuffer60 (.A(_06781_),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_1 rebuffer61 (.A(_06945_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(_06884_),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_1 rebuffer63 (.A(net586),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_2 rebuffer64 (.A(_06827_),
    .X(net3132));
 sky130_fd_sc_hd__clkbuf_1 rebuffer65 (.A(_07145_),
    .X(net3163));
 sky130_fd_sc_hd__clkbuf_2 rebuffer66 (.A(_07114_),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer67 (.A(_06624_),
    .X(net3237));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer68 (.A(_06886_),
    .X(net3246));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(net3246),
    .X(net3333));
 sky130_fd_sc_hd__clkbuf_1 rebuffer7 (.A(net530),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(_06846_),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(_06868_),
    .X(net3405));
 sky130_fd_sc_hd__clkbuf_1 rebuffer72 (.A(_06846_),
    .X(net3408));
 sky130_fd_sc_hd__buf_1 rebuffer8 (.A(net531),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(net532),
    .X(net533));
 sky130_fd_sc_hd__buf_2 split34 (.A(_07464_),
    .X(net558));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_125 (.HI(net125));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_126 (.HI(net126));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_127 (.HI(net127));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_128 (.HI(net128));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_129 (.HI(net129));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_130 (.HI(net130));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_131 (.HI(net131));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_132 (.HI(net132));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_133 (.HI(net133));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_134 (.HI(net134));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_135 (.HI(net135));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_136 (.HI(net136));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_137 (.HI(net137));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_138 (.HI(net138));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_139 (.HI(net139));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__buf_1 wire1 (.A(_02826_),
    .X(net1580));
 sky130_fd_sc_hd__buf_4 wire79 (.A(_06856_),
    .X(net79));
 sky130_fd_sc_hd__buf_2 wire80 (.A(_05008_),
    .X(net80));
 sky130_fd_sc_hd__buf_2 wire81 (.A(_04977_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 wire85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 wire86 (.A(_05442_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 wire88 (.A(net3970),
    .X(net88));
 assign o_rgb[0] = net90;
 assign o_rgb[10] = net98;
 assign o_rgb[11] = net99;
 assign o_rgb[12] = net100;
 assign o_rgb[13] = net101;
 assign o_rgb[16] = net102;
 assign o_rgb[17] = net103;
 assign o_rgb[18] = net104;
 assign o_rgb[19] = net105;
 assign o_rgb[1] = net91;
 assign o_rgb[20] = net106;
 assign o_rgb[21] = net107;
 assign o_rgb[2] = net92;
 assign o_rgb[3] = net93;
 assign o_rgb[4] = net94;
 assign o_rgb[5] = net95;
 assign o_rgb[8] = net96;
 assign o_rgb[9] = net97;
 assign ones[0] = net124;
 assign ones[10] = net134;
 assign ones[11] = net135;
 assign ones[12] = net136;
 assign ones[13] = net137;
 assign ones[14] = net138;
 assign ones[15] = net139;
 assign ones[1] = net125;
 assign ones[2] = net126;
 assign ones[3] = net127;
 assign ones[4] = net128;
 assign ones[5] = net129;
 assign ones[6] = net130;
 assign ones[7] = net131;
 assign ones[8] = net132;
 assign ones[9] = net133;
 assign zeros[0] = net108;
 assign zeros[10] = net118;
 assign zeros[11] = net119;
 assign zeros[12] = net120;
 assign zeros[13] = net121;
 assign zeros[14] = net122;
 assign zeros[15] = net123;
 assign zeros[1] = net109;
 assign zeros[2] = net110;
 assign zeros[3] = net111;
 assign zeros[4] = net112;
 assign zeros[5] = net113;
 assign zeros[6] = net114;
 assign zeros[7] = net115;
 assign zeros[8] = net116;
 assign zeros[9] = net117;
endmodule

