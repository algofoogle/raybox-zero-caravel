VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 588.790 BY 599.510 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 584.790 27.240 588.790 27.840 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 353.640 588.790 354.240 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 258.440 588.790 259.040 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 95.240 588.790 95.840 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 108.840 588.790 109.440 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 122.440 588.790 123.040 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 136.040 588.790 136.640 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 149.640 588.790 150.240 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 163.240 588.790 163.840 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 176.840 588.790 177.440 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 190.440 588.790 191.040 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 204.040 588.790 204.640 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 217.640 588.790 218.240 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 231.240 588.790 231.840 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 244.840 588.790 245.440 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 272.040 588.790 272.640 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 584.790 285.640 588.790 286.240 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 299.240 588.790 299.840 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 312.840 588.790 313.440 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 326.440 588.790 327.040 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 340.040 588.790 340.640 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 367.240 588.790 367.840 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 380.840 588.790 381.440 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 394.440 588.790 395.040 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 408.040 588.790 408.640 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 421.640 588.790 422.240 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 435.240 588.790 435.840 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 448.840 588.790 449.440 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 462.440 588.790 463.040 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 584.790 476.040 588.790 476.640 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 489.640 588.790 490.240 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 503.240 588.790 503.840 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 516.840 588.790 517.440 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 530.440 588.790 531.040 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 584.790 544.040 588.790 544.640 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 584.790 557.640 588.790 558.240 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 40.840 588.790 41.440 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 54.440 588.790 55.040 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 68.040 588.790 68.640 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 584.790 81.640 588.790 82.240 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 584.790 571.240 588.790 571.840 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 595.510 7.270 599.510 ;
    END
  END i_spare_1
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 595.510 55.110 599.510 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 42.870 595.510 43.150 599.510 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 30.910 595.510 31.190 599.510 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 595.510 19.230 599.510 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 126.590 595.510 126.870 599.510 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 114.630 595.510 114.910 599.510 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 102.670 595.510 102.950 599.510 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 90.710 595.510 90.990 599.510 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 78.750 595.510 79.030 599.510 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 66.790 595.510 67.070 599.510 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 198.350 595.510 198.630 599.510 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 174.430 595.510 174.710 599.510 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 162.470 595.510 162.750 599.510 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.510 595.510 150.790 599.510 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 138.550 595.510 138.830 599.510 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 186.390 595.510 186.670 599.510 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 595.510 581.350 599.510 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 595.510 461.750 599.510 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 595.510 449.790 599.510 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 595.510 437.830 599.510 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 595.510 425.870 599.510 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 595.510 413.910 599.510 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 595.510 401.950 599.510 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 595.510 569.390 599.510 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 595.510 557.430 599.510 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 595.510 545.470 599.510 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 595.510 533.510 599.510 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 595.510 521.550 599.510 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 595.510 509.590 599.510 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 595.510 497.630 599.510 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 595.510 485.670 599.510 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 595.510 473.710 599.510 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 595.510 389.990 599.510 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 595.510 270.390 599.510 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 595.510 258.430 599.510 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 595.510 246.470 599.510 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 595.510 234.510 599.510 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 595.510 222.550 599.510 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 595.510 210.590 599.510 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 595.510 378.030 599.510 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 595.510 366.070 599.510 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 595.510 354.110 599.510 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 595.510 342.150 599.510 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 595.510 330.190 599.510 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 595.510 318.230 599.510 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 595.510 306.270 599.510 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 595.510 294.310 599.510 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 595.510 282.350 599.510 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 583.010 586.215 ;
        RECT 5.330 577.945 583.010 580.775 ;
        RECT 5.330 572.505 583.010 575.335 ;
        RECT 5.330 567.065 583.010 569.895 ;
        RECT 5.330 561.625 583.010 564.455 ;
        RECT 5.330 556.185 583.010 559.015 ;
        RECT 5.330 550.745 583.010 553.575 ;
        RECT 5.330 545.305 583.010 548.135 ;
        RECT 5.330 539.865 583.010 542.695 ;
        RECT 5.330 534.425 583.010 537.255 ;
        RECT 5.330 528.985 583.010 531.815 ;
        RECT 5.330 523.545 583.010 526.375 ;
        RECT 5.330 518.105 583.010 520.935 ;
        RECT 5.330 512.665 583.010 515.495 ;
        RECT 5.330 507.225 583.010 510.055 ;
        RECT 5.330 501.785 583.010 504.615 ;
        RECT 5.330 496.345 583.010 499.175 ;
        RECT 5.330 490.905 583.010 493.735 ;
        RECT 5.330 485.465 583.010 488.295 ;
        RECT 5.330 480.025 583.010 482.855 ;
        RECT 5.330 474.585 583.010 477.415 ;
        RECT 5.330 469.145 583.010 471.975 ;
        RECT 5.330 463.705 583.010 466.535 ;
        RECT 5.330 458.265 583.010 461.095 ;
        RECT 5.330 452.825 583.010 455.655 ;
        RECT 5.330 447.385 583.010 450.215 ;
        RECT 5.330 441.945 583.010 444.775 ;
        RECT 5.330 436.505 583.010 439.335 ;
        RECT 5.330 431.065 583.010 433.895 ;
        RECT 5.330 425.625 583.010 428.455 ;
        RECT 5.330 420.185 583.010 423.015 ;
        RECT 5.330 414.745 583.010 417.575 ;
        RECT 5.330 409.305 583.010 412.135 ;
        RECT 5.330 403.865 583.010 406.695 ;
        RECT 5.330 398.425 583.010 401.255 ;
        RECT 5.330 392.985 583.010 395.815 ;
        RECT 5.330 387.545 583.010 390.375 ;
        RECT 5.330 382.105 583.010 384.935 ;
        RECT 5.330 376.665 583.010 379.495 ;
        RECT 5.330 371.225 583.010 374.055 ;
        RECT 5.330 365.785 583.010 368.615 ;
        RECT 5.330 360.345 583.010 363.175 ;
        RECT 5.330 354.905 583.010 357.735 ;
        RECT 5.330 349.465 583.010 352.295 ;
        RECT 5.330 344.025 583.010 346.855 ;
        RECT 5.330 338.585 583.010 341.415 ;
        RECT 5.330 333.145 583.010 335.975 ;
        RECT 5.330 327.705 583.010 330.535 ;
        RECT 5.330 322.265 583.010 325.095 ;
        RECT 5.330 316.825 583.010 319.655 ;
        RECT 5.330 311.385 583.010 314.215 ;
        RECT 5.330 305.945 583.010 308.775 ;
        RECT 5.330 300.505 583.010 303.335 ;
        RECT 5.330 295.065 583.010 297.895 ;
        RECT 5.330 289.625 583.010 292.455 ;
        RECT 5.330 284.185 583.010 287.015 ;
        RECT 5.330 278.745 583.010 281.575 ;
        RECT 5.330 273.305 583.010 276.135 ;
        RECT 5.330 267.865 583.010 270.695 ;
        RECT 5.330 262.425 583.010 265.255 ;
        RECT 5.330 256.985 583.010 259.815 ;
        RECT 5.330 251.545 583.010 254.375 ;
        RECT 5.330 246.105 583.010 248.935 ;
        RECT 5.330 240.665 583.010 243.495 ;
        RECT 5.330 235.225 583.010 238.055 ;
        RECT 5.330 229.785 583.010 232.615 ;
        RECT 5.330 224.345 583.010 227.175 ;
        RECT 5.330 218.905 583.010 221.735 ;
        RECT 5.330 213.465 583.010 216.295 ;
        RECT 5.330 208.025 583.010 210.855 ;
        RECT 5.330 202.585 583.010 205.415 ;
        RECT 5.330 197.145 583.010 199.975 ;
        RECT 5.330 191.705 583.010 194.535 ;
        RECT 5.330 186.265 583.010 189.095 ;
        RECT 5.330 180.825 583.010 183.655 ;
        RECT 5.330 175.385 583.010 178.215 ;
        RECT 5.330 169.945 583.010 172.775 ;
        RECT 5.330 164.505 583.010 167.335 ;
        RECT 5.330 159.065 583.010 161.895 ;
        RECT 5.330 153.625 583.010 156.455 ;
        RECT 5.330 148.185 583.010 151.015 ;
        RECT 5.330 142.745 583.010 145.575 ;
        RECT 5.330 137.305 583.010 140.135 ;
        RECT 5.330 131.865 583.010 134.695 ;
        RECT 5.330 126.425 583.010 129.255 ;
        RECT 5.330 120.985 583.010 123.815 ;
        RECT 5.330 115.545 583.010 118.375 ;
        RECT 5.330 110.105 583.010 112.935 ;
        RECT 5.330 104.665 583.010 107.495 ;
        RECT 5.330 99.225 583.010 102.055 ;
        RECT 5.330 93.785 583.010 96.615 ;
        RECT 5.330 88.345 583.010 91.175 ;
        RECT 5.330 82.905 583.010 85.735 ;
        RECT 5.330 77.465 583.010 80.295 ;
        RECT 5.330 72.025 583.010 74.855 ;
        RECT 5.330 66.585 583.010 69.415 ;
        RECT 5.330 61.145 583.010 63.975 ;
        RECT 5.330 55.705 583.010 58.535 ;
        RECT 5.330 50.265 583.010 53.095 ;
        RECT 5.330 44.825 583.010 47.655 ;
        RECT 5.330 39.385 583.010 42.215 ;
        RECT 5.330 33.945 583.010 36.775 ;
        RECT 5.330 28.505 583.010 31.335 ;
        RECT 5.330 23.065 583.010 25.895 ;
        RECT 5.330 17.625 583.010 20.455 ;
        RECT 5.330 12.185 583.010 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 582.820 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 585.050 596.320 ;
      LAYER met2 ;
        RECT 13.500 595.230 18.670 596.350 ;
        RECT 19.510 595.230 30.630 596.350 ;
        RECT 31.470 595.230 42.590 596.350 ;
        RECT 43.430 595.230 54.550 596.350 ;
        RECT 55.390 595.230 66.510 596.350 ;
        RECT 67.350 595.230 78.470 596.350 ;
        RECT 79.310 595.230 90.430 596.350 ;
        RECT 91.270 595.230 102.390 596.350 ;
        RECT 103.230 595.230 114.350 596.350 ;
        RECT 115.190 595.230 126.310 596.350 ;
        RECT 127.150 595.230 138.270 596.350 ;
        RECT 139.110 595.230 150.230 596.350 ;
        RECT 151.070 595.230 162.190 596.350 ;
        RECT 163.030 595.230 174.150 596.350 ;
        RECT 174.990 595.230 186.110 596.350 ;
        RECT 186.950 595.230 198.070 596.350 ;
        RECT 198.910 595.230 210.030 596.350 ;
        RECT 210.870 595.230 221.990 596.350 ;
        RECT 222.830 595.230 233.950 596.350 ;
        RECT 234.790 595.230 245.910 596.350 ;
        RECT 246.750 595.230 257.870 596.350 ;
        RECT 258.710 595.230 269.830 596.350 ;
        RECT 270.670 595.230 281.790 596.350 ;
        RECT 282.630 595.230 293.750 596.350 ;
        RECT 294.590 595.230 305.710 596.350 ;
        RECT 306.550 595.230 317.670 596.350 ;
        RECT 318.510 595.230 329.630 596.350 ;
        RECT 330.470 595.230 341.590 596.350 ;
        RECT 342.430 595.230 353.550 596.350 ;
        RECT 354.390 595.230 365.510 596.350 ;
        RECT 366.350 595.230 377.470 596.350 ;
        RECT 378.310 595.230 389.430 596.350 ;
        RECT 390.270 595.230 401.390 596.350 ;
        RECT 402.230 595.230 413.350 596.350 ;
        RECT 414.190 595.230 425.310 596.350 ;
        RECT 426.150 595.230 437.270 596.350 ;
        RECT 438.110 595.230 449.230 596.350 ;
        RECT 450.070 595.230 461.190 596.350 ;
        RECT 462.030 595.230 473.150 596.350 ;
        RECT 473.990 595.230 485.110 596.350 ;
        RECT 485.950 595.230 497.070 596.350 ;
        RECT 497.910 595.230 509.030 596.350 ;
        RECT 509.870 595.230 520.990 596.350 ;
        RECT 521.830 595.230 532.950 596.350 ;
        RECT 533.790 595.230 544.910 596.350 ;
        RECT 545.750 595.230 556.870 596.350 ;
        RECT 557.710 595.230 568.830 596.350 ;
        RECT 569.670 595.230 580.790 596.350 ;
        RECT 581.630 595.230 585.020 596.350 ;
        RECT 13.500 4.280 585.020 595.230 ;
        RECT 13.990 3.670 28.330 4.280 ;
        RECT 29.170 3.670 43.510 4.280 ;
        RECT 44.350 3.670 58.690 4.280 ;
        RECT 59.530 3.670 73.870 4.280 ;
        RECT 74.710 3.670 89.050 4.280 ;
        RECT 89.890 3.670 104.230 4.280 ;
        RECT 105.070 3.670 119.410 4.280 ;
        RECT 120.250 3.670 134.590 4.280 ;
        RECT 135.430 3.670 149.770 4.280 ;
        RECT 150.610 3.670 164.950 4.280 ;
        RECT 165.790 3.670 180.130 4.280 ;
        RECT 180.970 3.670 195.310 4.280 ;
        RECT 196.150 3.670 210.490 4.280 ;
        RECT 211.330 3.670 225.670 4.280 ;
        RECT 226.510 3.670 240.850 4.280 ;
        RECT 241.690 3.670 256.030 4.280 ;
        RECT 256.870 3.670 271.210 4.280 ;
        RECT 272.050 3.670 286.390 4.280 ;
        RECT 287.230 3.670 301.570 4.280 ;
        RECT 302.410 3.670 316.750 4.280 ;
        RECT 317.590 3.670 331.930 4.280 ;
        RECT 332.770 3.670 347.110 4.280 ;
        RECT 347.950 3.670 362.290 4.280 ;
        RECT 363.130 3.670 377.470 4.280 ;
        RECT 378.310 3.670 392.650 4.280 ;
        RECT 393.490 3.670 407.830 4.280 ;
        RECT 408.670 3.670 423.010 4.280 ;
        RECT 423.850 3.670 438.190 4.280 ;
        RECT 439.030 3.670 453.370 4.280 ;
        RECT 454.210 3.670 468.550 4.280 ;
        RECT 469.390 3.670 483.730 4.280 ;
        RECT 484.570 3.670 498.910 4.280 ;
        RECT 499.750 3.670 514.090 4.280 ;
        RECT 514.930 3.670 529.270 4.280 ;
        RECT 530.110 3.670 544.450 4.280 ;
        RECT 545.290 3.670 559.630 4.280 ;
        RECT 560.470 3.670 574.810 4.280 ;
        RECT 575.650 3.670 585.020 4.280 ;
      LAYER met3 ;
        RECT 17.545 572.240 584.790 588.705 ;
        RECT 17.545 570.840 584.390 572.240 ;
        RECT 17.545 558.640 584.790 570.840 ;
        RECT 17.545 557.240 584.390 558.640 ;
        RECT 17.545 545.040 584.790 557.240 ;
        RECT 17.545 543.640 584.390 545.040 ;
        RECT 17.545 531.440 584.790 543.640 ;
        RECT 17.545 530.040 584.390 531.440 ;
        RECT 17.545 517.840 584.790 530.040 ;
        RECT 17.545 516.440 584.390 517.840 ;
        RECT 17.545 504.240 584.790 516.440 ;
        RECT 17.545 502.840 584.390 504.240 ;
        RECT 17.545 490.640 584.790 502.840 ;
        RECT 17.545 489.240 584.390 490.640 ;
        RECT 17.545 477.040 584.790 489.240 ;
        RECT 17.545 475.640 584.390 477.040 ;
        RECT 17.545 463.440 584.790 475.640 ;
        RECT 17.545 462.040 584.390 463.440 ;
        RECT 17.545 449.840 584.790 462.040 ;
        RECT 17.545 448.440 584.390 449.840 ;
        RECT 17.545 436.240 584.790 448.440 ;
        RECT 17.545 434.840 584.390 436.240 ;
        RECT 17.545 422.640 584.790 434.840 ;
        RECT 17.545 421.240 584.390 422.640 ;
        RECT 17.545 409.040 584.790 421.240 ;
        RECT 17.545 407.640 584.390 409.040 ;
        RECT 17.545 395.440 584.790 407.640 ;
        RECT 17.545 394.040 584.390 395.440 ;
        RECT 17.545 381.840 584.790 394.040 ;
        RECT 17.545 380.440 584.390 381.840 ;
        RECT 17.545 368.240 584.790 380.440 ;
        RECT 17.545 366.840 584.390 368.240 ;
        RECT 17.545 354.640 584.790 366.840 ;
        RECT 17.545 353.240 584.390 354.640 ;
        RECT 17.545 341.040 584.790 353.240 ;
        RECT 17.545 339.640 584.390 341.040 ;
        RECT 17.545 327.440 584.790 339.640 ;
        RECT 17.545 326.040 584.390 327.440 ;
        RECT 17.545 313.840 584.790 326.040 ;
        RECT 17.545 312.440 584.390 313.840 ;
        RECT 17.545 300.240 584.790 312.440 ;
        RECT 17.545 298.840 584.390 300.240 ;
        RECT 17.545 286.640 584.790 298.840 ;
        RECT 17.545 285.240 584.390 286.640 ;
        RECT 17.545 273.040 584.790 285.240 ;
        RECT 17.545 271.640 584.390 273.040 ;
        RECT 17.545 259.440 584.790 271.640 ;
        RECT 17.545 258.040 584.390 259.440 ;
        RECT 17.545 245.840 584.790 258.040 ;
        RECT 17.545 244.440 584.390 245.840 ;
        RECT 17.545 232.240 584.790 244.440 ;
        RECT 17.545 230.840 584.390 232.240 ;
        RECT 17.545 218.640 584.790 230.840 ;
        RECT 17.545 217.240 584.390 218.640 ;
        RECT 17.545 205.040 584.790 217.240 ;
        RECT 17.545 203.640 584.390 205.040 ;
        RECT 17.545 191.440 584.790 203.640 ;
        RECT 17.545 190.040 584.390 191.440 ;
        RECT 17.545 177.840 584.790 190.040 ;
        RECT 17.545 176.440 584.390 177.840 ;
        RECT 17.545 164.240 584.790 176.440 ;
        RECT 17.545 162.840 584.390 164.240 ;
        RECT 17.545 150.640 584.790 162.840 ;
        RECT 17.545 149.240 584.390 150.640 ;
        RECT 17.545 137.040 584.790 149.240 ;
        RECT 17.545 135.640 584.390 137.040 ;
        RECT 17.545 123.440 584.790 135.640 ;
        RECT 17.545 122.040 584.390 123.440 ;
        RECT 17.545 109.840 584.790 122.040 ;
        RECT 17.545 108.440 584.390 109.840 ;
        RECT 17.545 96.240 584.790 108.440 ;
        RECT 17.545 94.840 584.390 96.240 ;
        RECT 17.545 82.640 584.790 94.840 ;
        RECT 17.545 81.240 584.390 82.640 ;
        RECT 17.545 69.040 584.790 81.240 ;
        RECT 17.545 67.640 584.390 69.040 ;
        RECT 17.545 55.440 584.790 67.640 ;
        RECT 17.545 54.040 584.390 55.440 ;
        RECT 17.545 41.840 584.790 54.040 ;
        RECT 17.545 40.440 584.390 41.840 ;
        RECT 17.545 28.240 584.790 40.440 ;
        RECT 17.545 26.840 584.390 28.240 ;
        RECT 17.545 10.715 584.790 26.840 ;
      LAYER met4 ;
        RECT 32.495 13.095 97.440 581.225 ;
        RECT 99.840 13.095 174.240 581.225 ;
        RECT 176.640 13.095 251.040 581.225 ;
        RECT 253.440 13.095 327.840 581.225 ;
        RECT 330.240 13.095 404.640 581.225 ;
        RECT 407.040 13.095 481.440 581.225 ;
        RECT 483.840 13.095 558.240 581.225 ;
        RECT 560.640 13.095 573.785 581.225 ;
  END
END top_ew_algofoogle
END LIBRARY

