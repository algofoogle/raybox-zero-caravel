VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 587.350 BY 598.070 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 12.960 587.350 13.560 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 355.680 587.350 356.280 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 255.720 587.350 256.320 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 84.360 587.350 84.960 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 98.640 587.350 99.240 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 112.920 587.350 113.520 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 127.200 587.350 127.800 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 141.480 587.350 142.080 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 155.760 587.350 156.360 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 170.040 587.350 170.640 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 184.320 587.350 184.920 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 198.600 587.350 199.200 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 212.880 587.350 213.480 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 227.160 587.350 227.760 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 241.440 587.350 242.040 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 270.000 587.350 270.600 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 284.280 587.350 284.880 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 298.560 587.350 299.160 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 312.840 587.350 313.440 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 327.120 587.350 327.720 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 341.400 587.350 342.000 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 369.960 587.350 370.560 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 384.240 587.350 384.840 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 398.520 587.350 399.120 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 412.800 587.350 413.400 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 427.080 587.350 427.680 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 441.360 587.350 441.960 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 455.640 587.350 456.240 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 469.920 587.350 470.520 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 484.200 587.350 484.800 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 498.480 587.350 499.080 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 512.760 587.350 513.360 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 527.040 587.350 527.640 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 541.320 587.350 541.920 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 555.600 587.350 556.200 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 569.880 587.350 570.480 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 27.240 587.350 27.840 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 41.520 587.350 42.120 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 55.800 587.350 56.400 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 70.080 587.350 70.680 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.350 584.160 587.350 584.760 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 594.070 6.810 598.070 ;
    END
  END i_spare_1
  PIN i_test_wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END i_test_wb_clk_i
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 594.070 54.650 598.070 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 594.070 42.690 598.070 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 594.070 30.730 598.070 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 594.070 18.770 598.070 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 594.070 126.410 598.070 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 594.070 114.450 598.070 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 594.070 102.490 598.070 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 594.070 90.530 598.070 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 594.070 78.570 598.070 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 594.070 66.610 598.070 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 594.070 198.170 598.070 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 594.070 174.250 598.070 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 594.070 162.290 598.070 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 594.070 150.330 598.070 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 594.070 138.370 598.070 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 594.070 186.210 598.070 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 594.070 580.890 598.070 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 594.070 461.290 598.070 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 594.070 449.330 598.070 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 594.070 437.370 598.070 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 594.070 425.410 598.070 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 594.070 413.450 598.070 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 594.070 401.490 598.070 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 594.070 568.930 598.070 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 594.070 556.970 598.070 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 594.070 545.010 598.070 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 594.070 533.050 598.070 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 594.070 521.090 598.070 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 594.070 509.130 598.070 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 594.070 497.170 598.070 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 594.070 485.210 598.070 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 594.070 473.250 598.070 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 585.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 585.040 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 594.070 389.530 598.070 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 594.070 269.930 598.070 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 594.070 257.970 598.070 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 594.070 246.010 598.070 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 594.070 234.050 598.070 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 594.070 222.090 598.070 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 594.070 210.130 598.070 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 594.070 377.570 598.070 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 594.070 365.610 598.070 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 594.070 353.650 598.070 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 594.070 341.690 598.070 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 594.070 329.730 598.070 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 594.070 317.770 598.070 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 594.070 305.810 598.070 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 594.070 293.850 598.070 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 594.070 281.890 598.070 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 581.630 584.990 ;
        RECT 5.330 577.945 581.630 580.775 ;
        RECT 5.330 572.505 581.630 575.335 ;
        RECT 5.330 567.065 581.630 569.895 ;
        RECT 5.330 561.625 581.630 564.455 ;
        RECT 5.330 556.185 581.630 559.015 ;
        RECT 5.330 550.745 581.630 553.575 ;
        RECT 5.330 545.305 581.630 548.135 ;
        RECT 5.330 539.865 581.630 542.695 ;
        RECT 5.330 534.425 581.630 537.255 ;
        RECT 5.330 528.985 581.630 531.815 ;
        RECT 5.330 523.545 581.630 526.375 ;
        RECT 5.330 518.105 581.630 520.935 ;
        RECT 5.330 512.665 581.630 515.495 ;
        RECT 5.330 507.225 581.630 510.055 ;
        RECT 5.330 501.785 581.630 504.615 ;
        RECT 5.330 496.345 581.630 499.175 ;
        RECT 5.330 490.905 581.630 493.735 ;
        RECT 5.330 485.465 581.630 488.295 ;
        RECT 5.330 480.025 581.630 482.855 ;
        RECT 5.330 474.585 581.630 477.415 ;
        RECT 5.330 469.145 581.630 471.975 ;
        RECT 5.330 463.705 581.630 466.535 ;
        RECT 5.330 458.265 581.630 461.095 ;
        RECT 5.330 452.825 581.630 455.655 ;
        RECT 5.330 447.385 581.630 450.215 ;
        RECT 5.330 441.945 581.630 444.775 ;
        RECT 5.330 436.505 581.630 439.335 ;
        RECT 5.330 431.065 581.630 433.895 ;
        RECT 5.330 425.625 581.630 428.455 ;
        RECT 5.330 420.185 581.630 423.015 ;
        RECT 5.330 414.745 581.630 417.575 ;
        RECT 5.330 409.305 581.630 412.135 ;
        RECT 5.330 403.865 581.630 406.695 ;
        RECT 5.330 398.425 581.630 401.255 ;
        RECT 5.330 392.985 581.630 395.815 ;
        RECT 5.330 387.545 581.630 390.375 ;
        RECT 5.330 382.105 581.630 384.935 ;
        RECT 5.330 376.665 581.630 379.495 ;
        RECT 5.330 371.225 581.630 374.055 ;
        RECT 5.330 365.785 581.630 368.615 ;
        RECT 5.330 360.345 581.630 363.175 ;
        RECT 5.330 354.905 581.630 357.735 ;
        RECT 5.330 349.465 581.630 352.295 ;
        RECT 5.330 344.025 581.630 346.855 ;
        RECT 5.330 338.585 581.630 341.415 ;
        RECT 5.330 333.145 581.630 335.975 ;
        RECT 5.330 327.705 581.630 330.535 ;
        RECT 5.330 322.265 581.630 325.095 ;
        RECT 5.330 316.825 581.630 319.655 ;
        RECT 5.330 311.385 581.630 314.215 ;
        RECT 5.330 305.945 581.630 308.775 ;
        RECT 5.330 300.505 581.630 303.335 ;
        RECT 5.330 295.065 581.630 297.895 ;
        RECT 5.330 289.625 581.630 292.455 ;
        RECT 5.330 284.185 581.630 287.015 ;
        RECT 5.330 278.745 581.630 281.575 ;
        RECT 5.330 273.305 581.630 276.135 ;
        RECT 5.330 267.865 581.630 270.695 ;
        RECT 5.330 262.425 581.630 265.255 ;
        RECT 5.330 256.985 581.630 259.815 ;
        RECT 5.330 251.545 581.630 254.375 ;
        RECT 5.330 246.105 581.630 248.935 ;
        RECT 5.330 240.665 581.630 243.495 ;
        RECT 5.330 235.225 581.630 238.055 ;
        RECT 5.330 229.785 581.630 232.615 ;
        RECT 5.330 224.345 581.630 227.175 ;
        RECT 5.330 218.905 581.630 221.735 ;
        RECT 5.330 213.465 581.630 216.295 ;
        RECT 5.330 208.025 581.630 210.855 ;
        RECT 5.330 202.585 581.630 205.415 ;
        RECT 5.330 197.145 581.630 199.975 ;
        RECT 5.330 191.705 581.630 194.535 ;
        RECT 5.330 186.265 581.630 189.095 ;
        RECT 5.330 180.825 581.630 183.655 ;
        RECT 5.330 175.385 581.630 178.215 ;
        RECT 5.330 169.945 581.630 172.775 ;
        RECT 5.330 164.505 581.630 167.335 ;
        RECT 5.330 159.065 581.630 161.895 ;
        RECT 5.330 153.625 581.630 156.455 ;
        RECT 5.330 148.185 581.630 151.015 ;
        RECT 5.330 142.745 581.630 145.575 ;
        RECT 5.330 137.305 581.630 140.135 ;
        RECT 5.330 131.865 581.630 134.695 ;
        RECT 5.330 126.425 581.630 129.255 ;
        RECT 5.330 120.985 581.630 123.815 ;
        RECT 5.330 115.545 581.630 118.375 ;
        RECT 5.330 110.105 581.630 112.935 ;
        RECT 5.330 104.665 581.630 107.495 ;
        RECT 5.330 99.225 581.630 102.055 ;
        RECT 5.330 93.785 581.630 96.615 ;
        RECT 5.330 88.345 581.630 91.175 ;
        RECT 5.330 82.905 581.630 85.735 ;
        RECT 5.330 77.465 581.630 80.295 ;
        RECT 5.330 72.025 581.630 74.855 ;
        RECT 5.330 66.585 581.630 69.415 ;
        RECT 5.330 61.145 581.630 63.975 ;
        RECT 5.330 55.705 581.630 58.535 ;
        RECT 5.330 50.265 581.630 53.095 ;
        RECT 5.330 44.825 581.630 47.655 ;
        RECT 5.330 39.385 581.630 42.215 ;
        RECT 5.330 33.945 581.630 36.775 ;
        RECT 5.330 28.505 581.630 31.335 ;
        RECT 5.330 23.065 581.630 25.895 ;
        RECT 5.330 17.625 581.630 20.455 ;
        RECT 5.330 12.185 581.630 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 581.440 584.885 ;
      LAYER met1 ;
        RECT 5.520 9.220 581.440 585.040 ;
      LAYER met2 ;
        RECT 9.300 593.790 18.210 594.730 ;
        RECT 19.050 593.790 30.170 594.730 ;
        RECT 31.010 593.790 42.130 594.730 ;
        RECT 42.970 593.790 54.090 594.730 ;
        RECT 54.930 593.790 66.050 594.730 ;
        RECT 66.890 593.790 78.010 594.730 ;
        RECT 78.850 593.790 89.970 594.730 ;
        RECT 90.810 593.790 101.930 594.730 ;
        RECT 102.770 593.790 113.890 594.730 ;
        RECT 114.730 593.790 125.850 594.730 ;
        RECT 126.690 593.790 137.810 594.730 ;
        RECT 138.650 593.790 149.770 594.730 ;
        RECT 150.610 593.790 161.730 594.730 ;
        RECT 162.570 593.790 173.690 594.730 ;
        RECT 174.530 593.790 185.650 594.730 ;
        RECT 186.490 593.790 197.610 594.730 ;
        RECT 198.450 593.790 209.570 594.730 ;
        RECT 210.410 593.790 221.530 594.730 ;
        RECT 222.370 593.790 233.490 594.730 ;
        RECT 234.330 593.790 245.450 594.730 ;
        RECT 246.290 593.790 257.410 594.730 ;
        RECT 258.250 593.790 269.370 594.730 ;
        RECT 270.210 593.790 281.330 594.730 ;
        RECT 282.170 593.790 293.290 594.730 ;
        RECT 294.130 593.790 305.250 594.730 ;
        RECT 306.090 593.790 317.210 594.730 ;
        RECT 318.050 593.790 329.170 594.730 ;
        RECT 330.010 593.790 341.130 594.730 ;
        RECT 341.970 593.790 353.090 594.730 ;
        RECT 353.930 593.790 365.050 594.730 ;
        RECT 365.890 593.790 377.010 594.730 ;
        RECT 377.850 593.790 388.970 594.730 ;
        RECT 389.810 593.790 400.930 594.730 ;
        RECT 401.770 593.790 412.890 594.730 ;
        RECT 413.730 593.790 424.850 594.730 ;
        RECT 425.690 593.790 436.810 594.730 ;
        RECT 437.650 593.790 448.770 594.730 ;
        RECT 449.610 593.790 460.730 594.730 ;
        RECT 461.570 593.790 472.690 594.730 ;
        RECT 473.530 593.790 484.650 594.730 ;
        RECT 485.490 593.790 496.610 594.730 ;
        RECT 497.450 593.790 508.570 594.730 ;
        RECT 509.410 593.790 520.530 594.730 ;
        RECT 521.370 593.790 532.490 594.730 ;
        RECT 533.330 593.790 544.450 594.730 ;
        RECT 545.290 593.790 556.410 594.730 ;
        RECT 557.250 593.790 568.370 594.730 ;
        RECT 569.210 593.790 580.330 594.730 ;
        RECT 9.300 4.280 580.880 593.790 ;
        RECT 9.300 4.000 13.610 4.280 ;
        RECT 14.450 4.000 28.330 4.280 ;
        RECT 29.170 4.000 43.050 4.280 ;
        RECT 43.890 4.000 57.770 4.280 ;
        RECT 58.610 4.000 72.490 4.280 ;
        RECT 73.330 4.000 87.210 4.280 ;
        RECT 88.050 4.000 101.930 4.280 ;
        RECT 102.770 4.000 116.650 4.280 ;
        RECT 117.490 4.000 131.370 4.280 ;
        RECT 132.210 4.000 146.090 4.280 ;
        RECT 146.930 4.000 160.810 4.280 ;
        RECT 161.650 4.000 175.530 4.280 ;
        RECT 176.370 4.000 190.250 4.280 ;
        RECT 191.090 4.000 204.970 4.280 ;
        RECT 205.810 4.000 219.690 4.280 ;
        RECT 220.530 4.000 234.410 4.280 ;
        RECT 235.250 4.000 249.130 4.280 ;
        RECT 249.970 4.000 263.850 4.280 ;
        RECT 264.690 4.000 278.570 4.280 ;
        RECT 279.410 4.000 293.290 4.280 ;
        RECT 294.130 4.000 308.010 4.280 ;
        RECT 308.850 4.000 322.730 4.280 ;
        RECT 323.570 4.000 337.450 4.280 ;
        RECT 338.290 4.000 352.170 4.280 ;
        RECT 353.010 4.000 366.890 4.280 ;
        RECT 367.730 4.000 381.610 4.280 ;
        RECT 382.450 4.000 396.330 4.280 ;
        RECT 397.170 4.000 411.050 4.280 ;
        RECT 411.890 4.000 425.770 4.280 ;
        RECT 426.610 4.000 440.490 4.280 ;
        RECT 441.330 4.000 455.210 4.280 ;
        RECT 456.050 4.000 469.930 4.280 ;
        RECT 470.770 4.000 484.650 4.280 ;
        RECT 485.490 4.000 499.370 4.280 ;
        RECT 500.210 4.000 514.090 4.280 ;
        RECT 514.930 4.000 528.810 4.280 ;
        RECT 529.650 4.000 543.530 4.280 ;
        RECT 544.370 4.000 558.250 4.280 ;
        RECT 559.090 4.000 572.970 4.280 ;
        RECT 573.810 4.000 580.880 4.280 ;
      LAYER met3 ;
        RECT 21.050 583.760 582.950 584.965 ;
        RECT 21.050 570.880 583.350 583.760 ;
        RECT 21.050 569.480 582.950 570.880 ;
        RECT 21.050 556.600 583.350 569.480 ;
        RECT 21.050 555.200 582.950 556.600 ;
        RECT 21.050 542.320 583.350 555.200 ;
        RECT 21.050 540.920 582.950 542.320 ;
        RECT 21.050 528.040 583.350 540.920 ;
        RECT 21.050 526.640 582.950 528.040 ;
        RECT 21.050 513.760 583.350 526.640 ;
        RECT 21.050 512.360 582.950 513.760 ;
        RECT 21.050 499.480 583.350 512.360 ;
        RECT 21.050 498.080 582.950 499.480 ;
        RECT 21.050 485.200 583.350 498.080 ;
        RECT 21.050 483.800 582.950 485.200 ;
        RECT 21.050 470.920 583.350 483.800 ;
        RECT 21.050 469.520 582.950 470.920 ;
        RECT 21.050 456.640 583.350 469.520 ;
        RECT 21.050 455.240 582.950 456.640 ;
        RECT 21.050 442.360 583.350 455.240 ;
        RECT 21.050 440.960 582.950 442.360 ;
        RECT 21.050 428.080 583.350 440.960 ;
        RECT 21.050 426.680 582.950 428.080 ;
        RECT 21.050 413.800 583.350 426.680 ;
        RECT 21.050 412.400 582.950 413.800 ;
        RECT 21.050 399.520 583.350 412.400 ;
        RECT 21.050 398.120 582.950 399.520 ;
        RECT 21.050 385.240 583.350 398.120 ;
        RECT 21.050 383.840 582.950 385.240 ;
        RECT 21.050 370.960 583.350 383.840 ;
        RECT 21.050 369.560 582.950 370.960 ;
        RECT 21.050 356.680 583.350 369.560 ;
        RECT 21.050 355.280 582.950 356.680 ;
        RECT 21.050 342.400 583.350 355.280 ;
        RECT 21.050 341.000 582.950 342.400 ;
        RECT 21.050 328.120 583.350 341.000 ;
        RECT 21.050 326.720 582.950 328.120 ;
        RECT 21.050 313.840 583.350 326.720 ;
        RECT 21.050 312.440 582.950 313.840 ;
        RECT 21.050 299.560 583.350 312.440 ;
        RECT 21.050 298.160 582.950 299.560 ;
        RECT 21.050 285.280 583.350 298.160 ;
        RECT 21.050 283.880 582.950 285.280 ;
        RECT 21.050 271.000 583.350 283.880 ;
        RECT 21.050 269.600 582.950 271.000 ;
        RECT 21.050 256.720 583.350 269.600 ;
        RECT 21.050 255.320 582.950 256.720 ;
        RECT 21.050 242.440 583.350 255.320 ;
        RECT 21.050 241.040 582.950 242.440 ;
        RECT 21.050 228.160 583.350 241.040 ;
        RECT 21.050 226.760 582.950 228.160 ;
        RECT 21.050 213.880 583.350 226.760 ;
        RECT 21.050 212.480 582.950 213.880 ;
        RECT 21.050 199.600 583.350 212.480 ;
        RECT 21.050 198.200 582.950 199.600 ;
        RECT 21.050 185.320 583.350 198.200 ;
        RECT 21.050 183.920 582.950 185.320 ;
        RECT 21.050 171.040 583.350 183.920 ;
        RECT 21.050 169.640 582.950 171.040 ;
        RECT 21.050 156.760 583.350 169.640 ;
        RECT 21.050 155.360 582.950 156.760 ;
        RECT 21.050 142.480 583.350 155.360 ;
        RECT 21.050 141.080 582.950 142.480 ;
        RECT 21.050 128.200 583.350 141.080 ;
        RECT 21.050 126.800 582.950 128.200 ;
        RECT 21.050 113.920 583.350 126.800 ;
        RECT 21.050 112.520 582.950 113.920 ;
        RECT 21.050 99.640 583.350 112.520 ;
        RECT 21.050 98.240 582.950 99.640 ;
        RECT 21.050 85.360 583.350 98.240 ;
        RECT 21.050 83.960 582.950 85.360 ;
        RECT 21.050 71.080 583.350 83.960 ;
        RECT 21.050 69.680 582.950 71.080 ;
        RECT 21.050 56.800 583.350 69.680 ;
        RECT 21.050 55.400 582.950 56.800 ;
        RECT 21.050 42.520 583.350 55.400 ;
        RECT 21.050 41.120 582.950 42.520 ;
        RECT 21.050 28.240 583.350 41.120 ;
        RECT 21.050 26.840 582.950 28.240 ;
        RECT 21.050 13.960 583.350 26.840 ;
        RECT 21.050 12.560 582.950 13.960 ;
        RECT 21.050 10.715 583.350 12.560 ;
      LAYER met4 ;
        RECT 46.295 11.735 97.440 580.545 ;
        RECT 99.840 11.735 174.240 580.545 ;
        RECT 176.640 11.735 251.040 580.545 ;
        RECT 253.440 11.735 327.840 580.545 ;
        RECT 330.240 11.735 404.640 580.545 ;
        RECT 407.040 11.735 481.440 580.545 ;
        RECT 483.840 11.735 558.240 580.545 ;
        RECT 560.640 11.735 576.545 580.545 ;
  END
END top_ew_algofoogle
END LIBRARY

