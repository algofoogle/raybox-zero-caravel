magic
tech sky130A
magscale 1 2
timestamp 1699121585
<< nwell >>
rect 1066 116677 116510 117243
rect 1066 115589 116510 116155
rect 1066 114501 116510 115067
rect 1066 113413 116510 113979
rect 1066 112325 116510 112891
rect 1066 111237 116510 111803
rect 1066 110149 116510 110715
rect 1066 109061 116510 109627
rect 1066 107973 116510 108539
rect 1066 106885 116510 107451
rect 1066 105797 116510 106363
rect 1066 104709 116510 105275
rect 1066 103621 116510 104187
rect 1066 102533 116510 103099
rect 1066 101445 116510 102011
rect 1066 100357 116510 100923
rect 1066 99269 116510 99835
rect 1066 98181 116510 98747
rect 1066 97093 116510 97659
rect 1066 96005 116510 96571
rect 1066 94917 116510 95483
rect 1066 93829 116510 94395
rect 1066 92741 116510 93307
rect 1066 91653 116510 92219
rect 1066 90565 116510 91131
rect 1066 89477 116510 90043
rect 1066 88389 116510 88955
rect 1066 87301 116510 87867
rect 1066 86213 116510 86779
rect 1066 85125 116510 85691
rect 1066 84037 116510 84603
rect 1066 82949 116510 83515
rect 1066 81861 116510 82427
rect 1066 80773 116510 81339
rect 1066 79685 116510 80251
rect 1066 78597 116510 79163
rect 1066 77509 116510 78075
rect 1066 76421 116510 76987
rect 1066 75333 116510 75899
rect 1066 74245 116510 74811
rect 1066 73157 116510 73723
rect 1066 72069 116510 72635
rect 1066 70981 116510 71547
rect 1066 69893 116510 70459
rect 1066 68805 116510 69371
rect 1066 67717 116510 68283
rect 1066 66629 116510 67195
rect 1066 65541 116510 66107
rect 1066 64453 116510 65019
rect 1066 63365 116510 63931
rect 1066 62277 116510 62843
rect 1066 61189 116510 61755
rect 1066 60101 116510 60667
rect 1066 59013 116510 59579
rect 1066 57925 116510 58491
rect 1066 56837 116510 57403
rect 1066 55749 116510 56315
rect 1066 54661 116510 55227
rect 1066 53573 116510 54139
rect 1066 52485 116510 53051
rect 1066 51397 116510 51963
rect 1066 50309 116510 50875
rect 1066 49221 116510 49787
rect 1066 48133 116510 48699
rect 1066 47045 116510 47611
rect 1066 45957 116510 46523
rect 1066 44869 116510 45435
rect 1066 43781 116510 44347
rect 1066 42693 116510 43259
rect 1066 41605 116510 42171
rect 1066 40517 116510 41083
rect 1066 39429 116510 39995
rect 1066 38341 116510 38907
rect 1066 37253 116510 37819
rect 1066 36165 116510 36731
rect 1066 35077 116510 35643
rect 1066 33989 116510 34555
rect 1066 32901 116510 33467
rect 1066 31813 116510 32379
rect 1066 30725 116510 31291
rect 1066 29637 116510 30203
rect 1066 28549 116510 29115
rect 1066 27461 116510 28027
rect 1066 26373 116510 26939
rect 1066 25285 116510 25851
rect 1066 24197 116510 24763
rect 1066 23109 116510 23675
rect 1066 22021 116510 22587
rect 1066 20933 116510 21499
rect 1066 19845 116510 20411
rect 1066 18757 116510 19323
rect 1066 17669 116510 18235
rect 1066 16581 116510 17147
rect 1066 15493 116510 16059
rect 1066 14405 116510 14971
rect 1066 13317 116510 13883
rect 1066 12229 116510 12795
rect 1066 11141 116510 11707
rect 1066 10053 116510 10619
rect 1066 8965 116510 9531
rect 1066 7877 116510 8443
rect 1066 6789 116510 7355
rect 1066 5701 116510 6267
rect 1066 4613 116510 5179
rect 1066 3525 116510 4091
rect 1066 2437 116510 3003
<< obsli1 >>
rect 1104 2159 116472 117521
<< obsm1 >>
rect 1104 1980 116472 117552
<< metal2 >>
rect 2410 118933 2466 119733
rect 4710 118933 4766 119733
rect 7010 118933 7066 119733
rect 9310 118933 9366 119733
rect 11610 118933 11666 119733
rect 13910 118933 13966 119733
rect 16210 118933 16266 119733
rect 18510 118933 18566 119733
rect 20810 118933 20866 119733
rect 23110 118933 23166 119733
rect 25410 118933 25466 119733
rect 27710 118933 27766 119733
rect 30010 118933 30066 119733
rect 32310 118933 32366 119733
rect 34610 118933 34666 119733
rect 36910 118933 36966 119733
rect 39210 118933 39266 119733
rect 41510 118933 41566 119733
rect 43810 118933 43866 119733
rect 46110 118933 46166 119733
rect 48410 118933 48466 119733
rect 50710 118933 50766 119733
rect 53010 118933 53066 119733
rect 55310 118933 55366 119733
rect 57610 118933 57666 119733
rect 59910 118933 59966 119733
rect 62210 118933 62266 119733
rect 64510 118933 64566 119733
rect 66810 118933 66866 119733
rect 69110 118933 69166 119733
rect 71410 118933 71466 119733
rect 73710 118933 73766 119733
rect 76010 118933 76066 119733
rect 78310 118933 78366 119733
rect 80610 118933 80666 119733
rect 82910 118933 82966 119733
rect 85210 118933 85266 119733
rect 87510 118933 87566 119733
rect 89810 118933 89866 119733
rect 92110 118933 92166 119733
rect 94410 118933 94466 119733
rect 96710 118933 96766 119733
rect 99010 118933 99066 119733
rect 101310 118933 101366 119733
rect 103610 118933 103666 119733
rect 105910 118933 105966 119733
rect 108210 118933 108266 119733
rect 110510 118933 110566 119733
rect 112810 118933 112866 119733
rect 115110 118933 115166 119733
rect 2778 0 2834 800
rect 5722 0 5778 800
rect 8666 0 8722 800
rect 11610 0 11666 800
rect 14554 0 14610 800
rect 17498 0 17554 800
rect 20442 0 20498 800
rect 23386 0 23442 800
rect 26330 0 26386 800
rect 29274 0 29330 800
rect 32218 0 32274 800
rect 35162 0 35218 800
rect 38106 0 38162 800
rect 41050 0 41106 800
rect 43994 0 44050 800
rect 46938 0 46994 800
rect 49882 0 49938 800
rect 52826 0 52882 800
rect 55770 0 55826 800
rect 58714 0 58770 800
rect 61658 0 61714 800
rect 64602 0 64658 800
rect 67546 0 67602 800
rect 70490 0 70546 800
rect 73434 0 73490 800
rect 76378 0 76434 800
rect 79322 0 79378 800
rect 82266 0 82322 800
rect 85210 0 85266 800
rect 88154 0 88210 800
rect 91098 0 91154 800
rect 94042 0 94098 800
rect 96986 0 97042 800
rect 99930 0 99986 800
rect 102874 0 102930 800
rect 105818 0 105874 800
rect 108762 0 108818 800
rect 111706 0 111762 800
rect 114650 0 114706 800
<< obsm2 >>
rect 1584 118877 2354 119082
rect 2522 118877 4654 119082
rect 4822 118877 6954 119082
rect 7122 118877 9254 119082
rect 9422 118877 11554 119082
rect 11722 118877 13854 119082
rect 14022 118877 16154 119082
rect 16322 118877 18454 119082
rect 18622 118877 20754 119082
rect 20922 118877 23054 119082
rect 23222 118877 25354 119082
rect 25522 118877 27654 119082
rect 27822 118877 29954 119082
rect 30122 118877 32254 119082
rect 32422 118877 34554 119082
rect 34722 118877 36854 119082
rect 37022 118877 39154 119082
rect 39322 118877 41454 119082
rect 41622 118877 43754 119082
rect 43922 118877 46054 119082
rect 46222 118877 48354 119082
rect 48522 118877 50654 119082
rect 50822 118877 52954 119082
rect 53122 118877 55254 119082
rect 55422 118877 57554 119082
rect 57722 118877 59854 119082
rect 60022 118877 62154 119082
rect 62322 118877 64454 119082
rect 64622 118877 66754 119082
rect 66922 118877 69054 119082
rect 69222 118877 71354 119082
rect 71522 118877 73654 119082
rect 73822 118877 75954 119082
rect 76122 118877 78254 119082
rect 78422 118877 80554 119082
rect 80722 118877 82854 119082
rect 83022 118877 85154 119082
rect 85322 118877 87454 119082
rect 87622 118877 89754 119082
rect 89922 118877 92054 119082
rect 92222 118877 94354 119082
rect 94522 118877 96654 119082
rect 96822 118877 98954 119082
rect 99122 118877 101254 119082
rect 101422 118877 103554 119082
rect 103722 118877 105854 119082
rect 106022 118877 108154 119082
rect 108322 118877 110454 119082
rect 110622 118877 112754 119082
rect 112922 118877 115054 119082
rect 115222 118877 115992 119082
rect 1584 856 115992 118877
rect 1584 800 2722 856
rect 2890 800 5666 856
rect 5834 800 8610 856
rect 8778 800 11554 856
rect 11722 800 14498 856
rect 14666 800 17442 856
rect 17610 800 20386 856
rect 20554 800 23330 856
rect 23498 800 26274 856
rect 26442 800 29218 856
rect 29386 800 32162 856
rect 32330 800 35106 856
rect 35274 800 38050 856
rect 38218 800 40994 856
rect 41162 800 43938 856
rect 44106 800 46882 856
rect 47050 800 49826 856
rect 49994 800 52770 856
rect 52938 800 55714 856
rect 55882 800 58658 856
rect 58826 800 61602 856
rect 61770 800 64546 856
rect 64714 800 67490 856
rect 67658 800 70434 856
rect 70602 800 73378 856
rect 73546 800 76322 856
rect 76490 800 79266 856
rect 79434 800 82210 856
rect 82378 800 85154 856
rect 85322 800 88098 856
rect 88266 800 91042 856
rect 91210 800 93986 856
rect 94154 800 96930 856
rect 97098 800 99874 856
rect 100042 800 102818 856
rect 102986 800 105762 856
rect 105930 800 108706 856
rect 108874 800 111650 856
rect 111818 800 114594 856
rect 114762 800 115992 856
<< metal3 >>
rect 116789 116832 117589 116952
rect 116789 113976 117589 114096
rect 116789 111120 117589 111240
rect 116789 108264 117589 108384
rect 116789 105408 117589 105528
rect 116789 102552 117589 102672
rect 116789 99696 117589 99816
rect 116789 96840 117589 96960
rect 116789 93984 117589 94104
rect 116789 91128 117589 91248
rect 116789 88272 117589 88392
rect 116789 85416 117589 85536
rect 116789 82560 117589 82680
rect 116789 79704 117589 79824
rect 116789 76848 117589 76968
rect 116789 73992 117589 74112
rect 116789 71136 117589 71256
rect 116789 68280 117589 68400
rect 116789 65424 117589 65544
rect 116789 62568 117589 62688
rect 116789 59712 117589 59832
rect 116789 56856 117589 56976
rect 116789 54000 117589 54120
rect 116789 51144 117589 51264
rect 116789 48288 117589 48408
rect 116789 45432 117589 45552
rect 116789 42576 117589 42696
rect 116789 39720 117589 39840
rect 116789 36864 117589 36984
rect 116789 34008 117589 34128
rect 116789 31152 117589 31272
rect 116789 28296 117589 28416
rect 116789 25440 117589 25560
rect 116789 22584 117589 22704
rect 116789 19728 117589 19848
rect 116789 16872 117589 16992
rect 116789 14016 117589 14136
rect 116789 11160 117589 11280
rect 116789 8304 117589 8424
rect 116789 5448 117589 5568
rect 116789 2592 117589 2712
<< obsm3 >>
rect 2681 117032 116789 117537
rect 2681 116752 116709 117032
rect 2681 114176 116789 116752
rect 2681 113896 116709 114176
rect 2681 111320 116789 113896
rect 2681 111040 116709 111320
rect 2681 108464 116789 111040
rect 2681 108184 116709 108464
rect 2681 105608 116789 108184
rect 2681 105328 116709 105608
rect 2681 102752 116789 105328
rect 2681 102472 116709 102752
rect 2681 99896 116789 102472
rect 2681 99616 116709 99896
rect 2681 97040 116789 99616
rect 2681 96760 116709 97040
rect 2681 94184 116789 96760
rect 2681 93904 116709 94184
rect 2681 91328 116789 93904
rect 2681 91048 116709 91328
rect 2681 88472 116789 91048
rect 2681 88192 116709 88472
rect 2681 85616 116789 88192
rect 2681 85336 116709 85616
rect 2681 82760 116789 85336
rect 2681 82480 116709 82760
rect 2681 79904 116789 82480
rect 2681 79624 116709 79904
rect 2681 77048 116789 79624
rect 2681 76768 116709 77048
rect 2681 74192 116789 76768
rect 2681 73912 116709 74192
rect 2681 71336 116789 73912
rect 2681 71056 116709 71336
rect 2681 68480 116789 71056
rect 2681 68200 116709 68480
rect 2681 65624 116789 68200
rect 2681 65344 116709 65624
rect 2681 62768 116789 65344
rect 2681 62488 116709 62768
rect 2681 59912 116789 62488
rect 2681 59632 116709 59912
rect 2681 57056 116789 59632
rect 2681 56776 116709 57056
rect 2681 54200 116789 56776
rect 2681 53920 116709 54200
rect 2681 51344 116789 53920
rect 2681 51064 116709 51344
rect 2681 48488 116789 51064
rect 2681 48208 116709 48488
rect 2681 45632 116789 48208
rect 2681 45352 116709 45632
rect 2681 42776 116789 45352
rect 2681 42496 116709 42776
rect 2681 39920 116789 42496
rect 2681 39640 116709 39920
rect 2681 37064 116789 39640
rect 2681 36784 116709 37064
rect 2681 34208 116789 36784
rect 2681 33928 116709 34208
rect 2681 31352 116789 33928
rect 2681 31072 116709 31352
rect 2681 28496 116789 31072
rect 2681 28216 116709 28496
rect 2681 25640 116789 28216
rect 2681 25360 116709 25640
rect 2681 22784 116789 25360
rect 2681 22504 116709 22784
rect 2681 19928 116789 22504
rect 2681 19648 116709 19928
rect 2681 17072 116789 19648
rect 2681 16792 116709 17072
rect 2681 14216 116789 16792
rect 2681 13936 116709 14216
rect 2681 11360 116789 13936
rect 2681 11080 116709 11360
rect 2681 8504 116789 11080
rect 2681 8224 116709 8504
rect 2681 5648 116789 8224
rect 2681 5368 116709 5648
rect 2681 2792 116789 5368
rect 2681 2512 116709 2792
rect 2681 2143 116789 2512
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 9995 2347 19488 117061
rect 19968 2347 34848 117061
rect 35328 2347 50208 117061
rect 50688 2347 65568 117061
rect 66048 2347 80928 117061
rect 81408 2347 96288 117061
rect 96768 2347 111648 117061
rect 112128 2347 114021 117061
<< labels >>
rlabel metal2 s 115110 118933 115166 119733 6 i_clk
port 1 nsew signal input
rlabel metal3 s 116789 71136 117589 71256 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 116789 51144 117589 51264 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 116789 16872 117589 16992 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 116789 19728 117589 19848 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 116789 22584 117589 22704 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 116789 25440 117589 25560 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 116789 28296 117589 28416 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 116789 31152 117589 31272 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 116789 34008 117589 34128 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 116789 36864 117589 36984 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 116789 39720 117589 39840 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 116789 42576 117589 42696 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 116789 45432 117589 45552 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 116789 48288 117589 48408 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 116789 54000 117589 54120 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 116789 56856 117589 56976 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 116789 59712 117589 59832 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 116789 62568 117589 62688 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 116789 65424 117589 65544 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 116789 68280 117589 68400 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 116789 73992 117589 74112 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 116789 76848 117589 76968 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 116789 79704 117589 79824 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 116789 82560 117589 82680 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 116789 85416 117589 85536 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 116789 88272 117589 88392 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 116789 91128 117589 91248 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 116789 93984 117589 94104 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 116789 96840 117589 96960 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 116789 99696 117589 99816 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 116789 102552 117589 102672 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 116789 105408 117589 105528 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 116789 108264 117589 108384 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 116789 111120 117589 111240 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 116789 113976 117589 114096 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 116789 5448 117589 5568 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 116789 8304 117589 8424 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 116789 11160 117589 11280 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 116789 14016 117589 14136 6 i_reg_sclk
port 48 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal3 s 116789 116832 117589 116952 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 2410 118933 2466 119733 6 i_spare_1
port 52 nsew signal input
rlabel metal3 s 116789 2592 117589 2712 6 i_test_uc2
port 53 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 i_test_wci
port 54 nsew signal input
rlabel metal2 s 11610 118933 11666 119733 6 i_tex_in[0]
port 55 nsew signal input
rlabel metal2 s 9310 118933 9366 119733 6 i_tex_in[1]
port 56 nsew signal input
rlabel metal2 s 7010 118933 7066 119733 6 i_tex_in[2]
port 57 nsew signal input
rlabel metal2 s 4710 118933 4766 119733 6 i_tex_in[3]
port 58 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 i_vec_csb
port 59 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 i_vec_mosi
port 60 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 i_vec_sclk
port 61 nsew signal input
rlabel metal2 s 25410 118933 25466 119733 6 o_gpout[0]
port 62 nsew signal output
rlabel metal2 s 23110 118933 23166 119733 6 o_gpout[1]
port 63 nsew signal output
rlabel metal2 s 20810 118933 20866 119733 6 o_gpout[2]
port 64 nsew signal output
rlabel metal2 s 18510 118933 18566 119733 6 o_gpout[3]
port 65 nsew signal output
rlabel metal2 s 16210 118933 16266 119733 6 o_gpout[4]
port 66 nsew signal output
rlabel metal2 s 13910 118933 13966 119733 6 o_gpout[5]
port 67 nsew signal output
rlabel metal2 s 39210 118933 39266 119733 6 o_hsync
port 68 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 o_reset
port 69 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 o_rgb[0]
port 70 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 o_rgb[10]
port 71 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 o_rgb[11]
port 72 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 o_rgb[12]
port 73 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 o_rgb[13]
port 74 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 o_rgb[14]
port 75 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 o_rgb[15]
port 76 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 o_rgb[16]
port 77 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 o_rgb[17]
port 78 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 o_rgb[18]
port 79 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 o_rgb[19]
port 80 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 o_rgb[1]
port 81 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 o_rgb[20]
port 82 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 o_rgb[21]
port 83 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 o_rgb[22]
port 84 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 o_rgb[23]
port 85 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 o_rgb[2]
port 86 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 o_rgb[3]
port 87 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 o_rgb[4]
port 88 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 o_rgb[5]
port 89 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 o_rgb[6]
port 90 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 o_rgb[7]
port 91 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 o_rgb[8]
port 92 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 o_rgb[9]
port 93 nsew signal output
rlabel metal2 s 34610 118933 34666 119733 6 o_tex_csb
port 94 nsew signal output
rlabel metal2 s 32310 118933 32366 119733 6 o_tex_oeb0
port 95 nsew signal output
rlabel metal2 s 30010 118933 30066 119733 6 o_tex_out0
port 96 nsew signal output
rlabel metal2 s 27710 118933 27766 119733 6 o_tex_sclk
port 97 nsew signal output
rlabel metal2 s 36910 118933 36966 119733 6 o_vsync
port 98 nsew signal output
rlabel metal2 s 112810 118933 112866 119733 6 ones[0]
port 99 nsew signal output
rlabel metal2 s 89810 118933 89866 119733 6 ones[10]
port 100 nsew signal output
rlabel metal2 s 87510 118933 87566 119733 6 ones[11]
port 101 nsew signal output
rlabel metal2 s 85210 118933 85266 119733 6 ones[12]
port 102 nsew signal output
rlabel metal2 s 82910 118933 82966 119733 6 ones[13]
port 103 nsew signal output
rlabel metal2 s 80610 118933 80666 119733 6 ones[14]
port 104 nsew signal output
rlabel metal2 s 78310 118933 78366 119733 6 ones[15]
port 105 nsew signal output
rlabel metal2 s 110510 118933 110566 119733 6 ones[1]
port 106 nsew signal output
rlabel metal2 s 108210 118933 108266 119733 6 ones[2]
port 107 nsew signal output
rlabel metal2 s 105910 118933 105966 119733 6 ones[3]
port 108 nsew signal output
rlabel metal2 s 103610 118933 103666 119733 6 ones[4]
port 109 nsew signal output
rlabel metal2 s 101310 118933 101366 119733 6 ones[5]
port 110 nsew signal output
rlabel metal2 s 99010 118933 99066 119733 6 ones[6]
port 111 nsew signal output
rlabel metal2 s 96710 118933 96766 119733 6 ones[7]
port 112 nsew signal output
rlabel metal2 s 94410 118933 94466 119733 6 ones[8]
port 113 nsew signal output
rlabel metal2 s 92110 118933 92166 119733 6 ones[9]
port 114 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 116 nsew ground bidirectional
rlabel metal2 s 76010 118933 76066 119733 6 zeros[0]
port 117 nsew signal output
rlabel metal2 s 53010 118933 53066 119733 6 zeros[10]
port 118 nsew signal output
rlabel metal2 s 50710 118933 50766 119733 6 zeros[11]
port 119 nsew signal output
rlabel metal2 s 48410 118933 48466 119733 6 zeros[12]
port 120 nsew signal output
rlabel metal2 s 46110 118933 46166 119733 6 zeros[13]
port 121 nsew signal output
rlabel metal2 s 43810 118933 43866 119733 6 zeros[14]
port 122 nsew signal output
rlabel metal2 s 41510 118933 41566 119733 6 zeros[15]
port 123 nsew signal output
rlabel metal2 s 73710 118933 73766 119733 6 zeros[1]
port 124 nsew signal output
rlabel metal2 s 71410 118933 71466 119733 6 zeros[2]
port 125 nsew signal output
rlabel metal2 s 69110 118933 69166 119733 6 zeros[3]
port 126 nsew signal output
rlabel metal2 s 66810 118933 66866 119733 6 zeros[4]
port 127 nsew signal output
rlabel metal2 s 64510 118933 64566 119733 6 zeros[5]
port 128 nsew signal output
rlabel metal2 s 62210 118933 62266 119733 6 zeros[6]
port 129 nsew signal output
rlabel metal2 s 59910 118933 59966 119733 6 zeros[7]
port 130 nsew signal output
rlabel metal2 s 57610 118933 57666 119733 6 zeros[8]
port 131 nsew signal output
rlabel metal2 s 55310 118933 55366 119733 6 zeros[9]
port 132 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 117589 119733
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33513136
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_11_05_04_36/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1465168
<< end >>

