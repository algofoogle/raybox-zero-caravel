magic
tech sky130A
magscale 1 2
timestamp 1698582601
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 14 2128 119862 117552
<< metal2 >>
rect 1950 119200 2006 119800
rect 5814 119200 5870 119800
rect 9678 119200 9734 119800
rect 13542 119200 13598 119800
rect 16762 119200 16818 119800
rect 20626 119200 20682 119800
rect 24490 119200 24546 119800
rect 28354 119200 28410 119800
rect 32218 119200 32274 119800
rect 35438 119200 35494 119800
rect 39302 119200 39358 119800
rect 43166 119200 43222 119800
rect 47030 119200 47086 119800
rect 50894 119200 50950 119800
rect 54758 119200 54814 119800
rect 57978 119200 58034 119800
rect 61842 119200 61898 119800
rect 65706 119200 65762 119800
rect 69570 119200 69626 119800
rect 73434 119200 73490 119800
rect 77298 119200 77354 119800
rect 80518 119200 80574 119800
rect 84382 119200 84438 119800
rect 88246 119200 88302 119800
rect 92110 119200 92166 119800
rect 95974 119200 96030 119800
rect 99194 119200 99250 119800
rect 103058 119200 103114 119800
rect 106922 119200 106978 119800
rect 110786 119200 110842 119800
rect 114650 119200 114706 119800
rect 118514 119200 118570 119800
rect 18 200 74 800
rect 3238 200 3294 800
rect 7102 200 7158 800
rect 10966 200 11022 800
rect 14830 200 14886 800
rect 18694 200 18750 800
rect 21914 200 21970 800
rect 25778 200 25834 800
rect 29642 200 29698 800
rect 33506 200 33562 800
rect 37370 200 37426 800
rect 41234 200 41290 800
rect 44454 200 44510 800
rect 48318 200 48374 800
rect 52182 200 52238 800
rect 56046 200 56102 800
rect 59910 200 59966 800
rect 63774 200 63830 800
rect 66994 200 67050 800
rect 70858 200 70914 800
rect 74722 200 74778 800
rect 78586 200 78642 800
rect 82450 200 82506 800
rect 85670 200 85726 800
rect 89534 200 89590 800
rect 93398 200 93454 800
rect 97262 200 97318 800
rect 101126 200 101182 800
rect 104990 200 105046 800
rect 108210 200 108266 800
rect 112074 200 112130 800
rect 115938 200 115994 800
rect 119802 200 119858 800
<< obsm2 >>
rect 20 119856 119856 119898
rect 20 119144 1894 119856
rect 2062 119144 5758 119856
rect 5926 119144 9622 119856
rect 9790 119144 13486 119856
rect 13654 119144 16706 119856
rect 16874 119144 20570 119856
rect 20738 119144 24434 119856
rect 24602 119144 28298 119856
rect 28466 119144 32162 119856
rect 32330 119144 35382 119856
rect 35550 119144 39246 119856
rect 39414 119144 43110 119856
rect 43278 119144 46974 119856
rect 47142 119144 50838 119856
rect 51006 119144 54702 119856
rect 54870 119144 57922 119856
rect 58090 119144 61786 119856
rect 61954 119144 65650 119856
rect 65818 119144 69514 119856
rect 69682 119144 73378 119856
rect 73546 119144 77242 119856
rect 77410 119144 80462 119856
rect 80630 119144 84326 119856
rect 84494 119144 88190 119856
rect 88358 119144 92054 119856
rect 92222 119144 95918 119856
rect 96086 119144 99138 119856
rect 99306 119144 103002 119856
rect 103170 119144 106866 119856
rect 107034 119144 110730 119856
rect 110898 119144 114594 119856
rect 114762 119144 118458 119856
rect 118626 119144 119856 119856
rect 20 856 119856 119144
rect 130 800 3182 856
rect 3350 800 7046 856
rect 7214 800 10910 856
rect 11078 800 14774 856
rect 14942 800 18638 856
rect 18806 800 21858 856
rect 22026 800 25722 856
rect 25890 800 29586 856
rect 29754 800 33450 856
rect 33618 800 37314 856
rect 37482 800 41178 856
rect 41346 800 44398 856
rect 44566 800 48262 856
rect 48430 800 52126 856
rect 52294 800 55990 856
rect 56158 800 59854 856
rect 60022 800 63718 856
rect 63886 800 66938 856
rect 67106 800 70802 856
rect 70970 800 74666 856
rect 74834 800 78530 856
rect 78698 800 82394 856
rect 82562 800 85614 856
rect 85782 800 89478 856
rect 89646 800 93342 856
rect 93510 800 97206 856
rect 97374 800 101070 856
rect 101238 800 104934 856
rect 105102 800 108154 856
rect 108322 800 112018 856
rect 112186 800 115882 856
rect 116050 800 119746 856
<< metal3 >>
rect 200 118328 800 118448
rect 119200 118328 119800 118448
rect 200 114248 800 114368
rect 119200 114248 119800 114368
rect 200 110848 800 110968
rect 119200 110168 119800 110288
rect 200 106768 800 106888
rect 119200 106088 119800 106208
rect 200 102688 800 102808
rect 119200 102008 119800 102128
rect 200 98608 800 98728
rect 119200 97928 119800 98048
rect 200 94528 800 94648
rect 119200 94528 119800 94648
rect 200 90448 800 90568
rect 119200 90448 119800 90568
rect 200 87048 800 87168
rect 119200 86368 119800 86488
rect 200 82968 800 83088
rect 119200 82288 119800 82408
rect 200 78888 800 79008
rect 119200 78208 119800 78328
rect 200 74808 800 74928
rect 119200 74808 119800 74928
rect 200 70728 800 70848
rect 119200 70728 119800 70848
rect 200 67328 800 67448
rect 119200 66648 119800 66768
rect 200 63248 800 63368
rect 119200 62568 119800 62688
rect 200 59168 800 59288
rect 119200 58488 119800 58608
rect 200 55088 800 55208
rect 119200 54408 119800 54528
rect 200 51008 800 51128
rect 119200 51008 119800 51128
rect 200 46928 800 47048
rect 119200 46928 119800 47048
rect 200 43528 800 43648
rect 119200 42848 119800 42968
rect 200 39448 800 39568
rect 119200 38768 119800 38888
rect 200 35368 800 35488
rect 119200 34688 119800 34808
rect 200 31288 800 31408
rect 119200 30608 119800 30728
rect 200 27208 800 27328
rect 119200 27208 119800 27328
rect 200 23128 800 23248
rect 119200 23128 119800 23248
rect 200 19728 800 19848
rect 119200 19048 119800 19168
rect 200 15648 800 15768
rect 119200 14968 119800 15088
rect 200 11568 800 11688
rect 119200 10888 119800 11008
rect 200 7488 800 7608
rect 119200 7488 119800 7608
rect 200 3408 800 3528
rect 119200 3408 119800 3528
<< obsm3 >>
rect 880 118248 119120 118421
rect 800 114448 119200 118248
rect 880 114168 119120 114448
rect 800 111048 119200 114168
rect 880 110768 119200 111048
rect 800 110368 119200 110768
rect 800 110088 119120 110368
rect 800 106968 119200 110088
rect 880 106688 119200 106968
rect 800 106288 119200 106688
rect 800 106008 119120 106288
rect 800 102888 119200 106008
rect 880 102608 119200 102888
rect 800 102208 119200 102608
rect 800 101928 119120 102208
rect 800 98808 119200 101928
rect 880 98528 119200 98808
rect 800 98128 119200 98528
rect 800 97848 119120 98128
rect 800 94728 119200 97848
rect 880 94448 119120 94728
rect 800 90648 119200 94448
rect 880 90368 119120 90648
rect 800 87248 119200 90368
rect 880 86968 119200 87248
rect 800 86568 119200 86968
rect 800 86288 119120 86568
rect 800 83168 119200 86288
rect 880 82888 119200 83168
rect 800 82488 119200 82888
rect 800 82208 119120 82488
rect 800 79088 119200 82208
rect 880 78808 119200 79088
rect 800 78408 119200 78808
rect 800 78128 119120 78408
rect 800 75008 119200 78128
rect 880 74728 119120 75008
rect 800 70928 119200 74728
rect 880 70648 119120 70928
rect 800 67528 119200 70648
rect 880 67248 119200 67528
rect 800 66848 119200 67248
rect 800 66568 119120 66848
rect 800 63448 119200 66568
rect 880 63168 119200 63448
rect 800 62768 119200 63168
rect 800 62488 119120 62768
rect 800 59368 119200 62488
rect 880 59088 119200 59368
rect 800 58688 119200 59088
rect 800 58408 119120 58688
rect 800 55288 119200 58408
rect 880 55008 119200 55288
rect 800 54608 119200 55008
rect 800 54328 119120 54608
rect 800 51208 119200 54328
rect 880 50928 119120 51208
rect 800 47128 119200 50928
rect 880 46848 119120 47128
rect 800 43728 119200 46848
rect 880 43448 119200 43728
rect 800 43048 119200 43448
rect 800 42768 119120 43048
rect 800 39648 119200 42768
rect 880 39368 119200 39648
rect 800 38968 119200 39368
rect 800 38688 119120 38968
rect 800 35568 119200 38688
rect 880 35288 119200 35568
rect 800 34888 119200 35288
rect 800 34608 119120 34888
rect 800 31488 119200 34608
rect 880 31208 119200 31488
rect 800 30808 119200 31208
rect 800 30528 119120 30808
rect 800 27408 119200 30528
rect 880 27128 119120 27408
rect 800 23328 119200 27128
rect 880 23048 119120 23328
rect 800 19928 119200 23048
rect 880 19648 119200 19928
rect 800 19248 119200 19648
rect 800 18968 119120 19248
rect 800 15848 119200 18968
rect 880 15568 119200 15848
rect 800 15168 119200 15568
rect 800 14888 119120 15168
rect 800 11768 119200 14888
rect 880 11488 119200 11768
rect 800 11088 119200 11488
rect 800 10808 119120 11088
rect 800 7688 119200 10808
rect 880 7408 119120 7688
rect 800 3608 119200 7408
rect 880 3328 119120 3608
rect 800 2143 119200 3328
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 13123 2347 19488 109173
rect 19968 2347 34848 109173
rect 35328 2347 50208 109173
rect 50688 2347 65568 109173
rect 66048 2347 80928 109173
rect 81408 2347 96288 109173
rect 96768 2347 111629 109173
<< labels >>
rlabel metal3 s 119200 110168 119800 110288 6 i_clk
port 1 nsew signal input
rlabel metal3 s 119200 19048 119800 19168 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal2 s 29642 200 29698 800 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal3 s 119200 114248 119800 114368 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 44454 200 44510 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal3 s 119200 38768 119800 38888 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 57978 119200 58034 119800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal3 s 119200 34688 119800 34808 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal3 s 119200 62568 119800 62688 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal3 s 119200 97928 119800 98048 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal2 s 28354 119200 28410 119800 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal2 s 108210 200 108266 800 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal2 s 95974 119200 96030 119800 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal2 s 118514 119200 118570 119800 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 200 94528 800 94648 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal2 s 16762 119200 16818 119800 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal2 s 119802 200 119858 800 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal2 s 112074 200 112130 800 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 200 15648 800 15768 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal2 s 25778 200 25834 800 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal2 s 70858 200 70914 800 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 200 31288 800 31408 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal2 s 1950 119200 2006 119800 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 200 3408 800 3528 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal2 s 89534 200 89590 800 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 200 55088 800 55208 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 119200 70728 119800 70848 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal2 s 61842 119200 61898 119800 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 200 70728 800 70848 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 200 19728 800 19848 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 200 98608 800 98728 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal2 s 48318 200 48374 800 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 119200 118328 119800 118448 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal2 s 32218 119200 32274 119800 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal2 s 54758 119200 54814 119800 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal2 s 114650 119200 114706 119800 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal2 s 33506 200 33562 800 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal2 s 84382 119200 84438 119800 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal2 s 69570 119200 69626 119800 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 200 74808 800 74928 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 119200 7488 119800 7608 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 200 7488 800 7608 6 i_mode[1]
port 43 nsew signal input
rlabel metal2 s 97262 200 97318 800 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 200 87048 800 87168 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 200 67328 800 67448 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 119200 82288 119800 82408 6 i_reg_sclk
port 47 nsew signal input
rlabel metal3 s 119200 66648 119800 66768 6 i_reset_lock_a
port 48 nsew signal input
rlabel metal2 s 43166 119200 43222 119800 6 i_reset_lock_b
port 49 nsew signal input
rlabel metal2 s 47030 119200 47086 119800 6 i_tex_in[0]
port 50 nsew signal input
rlabel metal2 s 14830 200 14886 800 6 i_tex_in[1]
port 51 nsew signal input
rlabel metal3 s 119200 106088 119800 106208 6 i_tex_in[2]
port 52 nsew signal input
rlabel metal2 s 59910 200 59966 800 6 i_tex_in[3]
port 53 nsew signal input
rlabel metal2 s 74722 200 74778 800 6 i_vec_csb
port 54 nsew signal input
rlabel metal3 s 119200 46928 119800 47048 6 i_vec_mosi
port 55 nsew signal input
rlabel metal2 s 103058 119200 103114 119800 6 i_vec_sclk
port 56 nsew signal input
rlabel metal2 s 77298 119200 77354 119800 6 o_gpout[0]
port 57 nsew signal output
rlabel metal3 s 119200 86368 119800 86488 6 o_gpout[1]
port 58 nsew signal output
rlabel metal3 s 119200 90448 119800 90568 6 o_gpout[2]
port 59 nsew signal output
rlabel metal2 s 20626 119200 20682 119800 6 o_gpout[3]
port 60 nsew signal output
rlabel metal2 s 106922 119200 106978 119800 6 o_gpout[4]
port 61 nsew signal output
rlabel metal3 s 200 27208 800 27328 6 o_gpout[5]
port 62 nsew signal output
rlabel metal2 s 37370 200 37426 800 6 o_hsync
port 63 nsew signal output
rlabel metal3 s 119200 42848 119800 42968 6 o_reset
port 64 nsew signal output
rlabel metal3 s 119200 27208 119800 27328 6 o_rgb[0]
port 65 nsew signal output
rlabel metal2 s 13542 119200 13598 119800 6 o_rgb[10]
port 66 nsew signal output
rlabel metal2 s 50894 119200 50950 119800 6 o_rgb[11]
port 67 nsew signal output
rlabel metal2 s 115938 200 115994 800 6 o_rgb[12]
port 68 nsew signal output
rlabel metal3 s 119200 30608 119800 30728 6 o_rgb[13]
port 69 nsew signal output
rlabel metal3 s 200 78888 800 79008 6 o_rgb[14]
port 70 nsew signal output
rlabel metal3 s 200 63248 800 63368 6 o_rgb[15]
port 71 nsew signal output
rlabel metal2 s 101126 200 101182 800 6 o_rgb[16]
port 72 nsew signal output
rlabel metal2 s 52182 200 52238 800 6 o_rgb[17]
port 73 nsew signal output
rlabel metal2 s 35438 119200 35494 119800 6 o_rgb[18]
port 74 nsew signal output
rlabel metal3 s 200 90448 800 90568 6 o_rgb[19]
port 75 nsew signal output
rlabel metal3 s 200 51008 800 51128 6 o_rgb[1]
port 76 nsew signal output
rlabel metal3 s 119200 10888 119800 11008 6 o_rgb[20]
port 77 nsew signal output
rlabel metal3 s 200 11568 800 11688 6 o_rgb[21]
port 78 nsew signal output
rlabel metal2 s 9678 119200 9734 119800 6 o_rgb[22]
port 79 nsew signal output
rlabel metal2 s 65706 119200 65762 119800 6 o_rgb[23]
port 80 nsew signal output
rlabel metal2 s 85670 200 85726 800 6 o_rgb[2]
port 81 nsew signal output
rlabel metal2 s 10966 200 11022 800 6 o_rgb[3]
port 82 nsew signal output
rlabel metal3 s 200 46928 800 47048 6 o_rgb[4]
port 83 nsew signal output
rlabel metal3 s 119200 3408 119800 3528 6 o_rgb[5]
port 84 nsew signal output
rlabel metal3 s 119200 78208 119800 78328 6 o_rgb[6]
port 85 nsew signal output
rlabel metal3 s 119200 51008 119800 51128 6 o_rgb[7]
port 86 nsew signal output
rlabel metal2 s 93398 200 93454 800 6 o_rgb[8]
port 87 nsew signal output
rlabel metal3 s 200 82968 800 83088 6 o_rgb[9]
port 88 nsew signal output
rlabel metal3 s 119200 23128 119800 23248 6 o_tex_csb
port 89 nsew signal output
rlabel metal3 s 200 110848 800 110968 6 o_tex_oeb0
port 90 nsew signal output
rlabel metal3 s 119200 58488 119800 58608 6 o_tex_out0
port 91 nsew signal output
rlabel metal3 s 119200 94528 119800 94648 6 o_tex_sclk
port 92 nsew signal output
rlabel metal2 s 104990 200 105046 800 6 o_vsync
port 93 nsew signal output
rlabel metal3 s 119200 102008 119800 102128 6 ones[0]
port 94 nsew signal output
rlabel metal3 s 200 59168 800 59288 6 ones[10]
port 95 nsew signal output
rlabel metal3 s 200 118328 800 118448 6 ones[11]
port 96 nsew signal output
rlabel metal3 s 200 43528 800 43648 6 ones[12]
port 97 nsew signal output
rlabel metal2 s 18 200 74 800 6 ones[13]
port 98 nsew signal output
rlabel metal2 s 78586 200 78642 800 6 ones[14]
port 99 nsew signal output
rlabel metal3 s 200 23128 800 23248 6 ones[15]
port 100 nsew signal output
rlabel metal2 s 39302 119200 39358 119800 6 ones[1]
port 101 nsew signal output
rlabel metal2 s 80518 119200 80574 119800 6 ones[2]
port 102 nsew signal output
rlabel metal3 s 200 102688 800 102808 6 ones[3]
port 103 nsew signal output
rlabel metal2 s 18694 200 18750 800 6 ones[4]
port 104 nsew signal output
rlabel metal2 s 7102 200 7158 800 6 ones[5]
port 105 nsew signal output
rlabel metal2 s 99194 119200 99250 119800 6 ones[6]
port 106 nsew signal output
rlabel metal2 s 73434 119200 73490 119800 6 ones[7]
port 107 nsew signal output
rlabel metal2 s 56046 200 56102 800 6 ones[8]
port 108 nsew signal output
rlabel metal2 s 110786 119200 110842 119800 6 ones[9]
port 109 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 111 nsew ground bidirectional
rlabel metal3 s 119200 14968 119800 15088 6 zeros[0]
port 112 nsew signal output
rlabel metal3 s 200 114248 800 114368 6 zeros[10]
port 113 nsew signal output
rlabel metal3 s 200 39448 800 39568 6 zeros[11]
port 114 nsew signal output
rlabel metal2 s 21914 200 21970 800 6 zeros[12]
port 115 nsew signal output
rlabel metal2 s 41234 200 41290 800 6 zeros[13]
port 116 nsew signal output
rlabel metal2 s 63774 200 63830 800 6 zeros[14]
port 117 nsew signal output
rlabel metal3 s 119200 74808 119800 74928 6 zeros[15]
port 118 nsew signal output
rlabel metal2 s 66994 200 67050 800 6 zeros[1]
port 119 nsew signal output
rlabel metal2 s 92110 119200 92166 119800 6 zeros[2]
port 120 nsew signal output
rlabel metal2 s 88246 119200 88302 119800 6 zeros[3]
port 121 nsew signal output
rlabel metal2 s 5814 119200 5870 119800 6 zeros[4]
port 122 nsew signal output
rlabel metal2 s 24490 119200 24546 119800 6 zeros[5]
port 123 nsew signal output
rlabel metal2 s 82450 200 82506 800 6 zeros[6]
port 124 nsew signal output
rlabel metal3 s 200 35368 800 35488 6 zeros[7]
port 125 nsew signal output
rlabel metal3 s 200 106768 800 106888 6 zeros[8]
port 126 nsew signal output
rlabel metal3 s 119200 54408 119800 54528 6 zeros[9]
port 127 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32119276
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_10_29_22_55/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1541948
<< end >>

