magic
tech sky130A
magscale 1 2
timestamp 1698805415
<< nwell >>
rect 1066 111237 111266 111803
rect 1066 110149 111266 110715
rect 1066 109061 111266 109627
rect 1066 107973 111266 108539
rect 1066 106885 111266 107451
rect 1066 105797 111266 106363
rect 1066 104709 111266 105275
rect 1066 103621 111266 104187
rect 1066 102533 111266 103099
rect 1066 101445 111266 102011
rect 1066 100357 111266 100923
rect 1066 99269 111266 99835
rect 1066 98181 111266 98747
rect 1066 97093 111266 97659
rect 1066 96005 111266 96571
rect 1066 94917 111266 95483
rect 1066 93829 111266 94395
rect 1066 92741 111266 93307
rect 1066 91653 111266 92219
rect 1066 90565 111266 91131
rect 1066 89477 111266 90043
rect 1066 88389 111266 88955
rect 1066 87301 111266 87867
rect 1066 86213 111266 86779
rect 1066 85125 111266 85691
rect 1066 84037 111266 84603
rect 1066 82949 111266 83515
rect 1066 81861 111266 82427
rect 1066 80773 111266 81339
rect 1066 79685 111266 80251
rect 1066 78597 111266 79163
rect 1066 77509 111266 78075
rect 1066 76421 111266 76987
rect 1066 75333 111266 75899
rect 1066 74245 111266 74811
rect 1066 73157 111266 73723
rect 1066 72069 111266 72635
rect 1066 70981 111266 71547
rect 1066 69893 111266 70459
rect 1066 68805 111266 69371
rect 1066 67717 111266 68283
rect 1066 66629 111266 67195
rect 1066 65541 111266 66107
rect 1066 64453 111266 65019
rect 1066 63365 111266 63931
rect 1066 62277 111266 62843
rect 1066 61189 111266 61755
rect 1066 60101 111266 60667
rect 1066 59013 111266 59579
rect 1066 57925 111266 58491
rect 1066 56837 111266 57403
rect 1066 55749 111266 56315
rect 1066 54661 111266 55227
rect 1066 53573 111266 54139
rect 1066 52485 111266 53051
rect 1066 51397 111266 51963
rect 1066 50309 111266 50875
rect 1066 49221 111266 49787
rect 1066 48133 111266 48699
rect 1066 47045 111266 47611
rect 1066 45957 111266 46523
rect 1066 44869 111266 45435
rect 1066 43781 111266 44347
rect 1066 42693 111266 43259
rect 1066 41605 111266 42171
rect 1066 40517 111266 41083
rect 1066 39429 111266 39995
rect 1066 38341 111266 38907
rect 1066 37253 111266 37819
rect 1066 36165 111266 36731
rect 1066 35077 111266 35643
rect 1066 33989 111266 34555
rect 1066 32901 111266 33467
rect 1066 31813 111266 32379
rect 1066 30725 111266 31291
rect 1066 29637 111266 30203
rect 1066 28549 111266 29115
rect 1066 27461 111266 28027
rect 1066 26373 111266 26939
rect 1066 25285 111266 25851
rect 1066 24197 111266 24763
rect 1066 23109 111266 23675
rect 1066 22021 111266 22587
rect 1066 20933 111266 21499
rect 1066 19845 111266 20411
rect 1066 18757 111266 19323
rect 1066 17669 111266 18235
rect 1066 16581 111266 17147
rect 1066 15493 111266 16059
rect 1066 14405 111266 14971
rect 1066 13317 111266 13883
rect 1066 12229 111266 12795
rect 1066 11141 111266 11707
rect 1066 10053 111266 10619
rect 1066 8965 111266 9531
rect 1066 7877 111266 8443
rect 1066 6789 111266 7355
rect 1066 5701 111266 6267
rect 1066 4613 111266 5179
rect 1066 3525 111266 4091
rect 1066 2437 111266 3003
<< obsli1 >>
rect 1104 2159 111228 112081
<< obsm1 >>
rect 1104 1912 111228 112112
<< metal2 >>
rect 2042 113686 2098 114486
rect 4342 113686 4398 114486
rect 6642 113686 6698 114486
rect 8942 113686 8998 114486
rect 11242 113686 11298 114486
rect 13542 113686 13598 114486
rect 15842 113686 15898 114486
rect 18142 113686 18198 114486
rect 20442 113686 20498 114486
rect 22742 113686 22798 114486
rect 25042 113686 25098 114486
rect 27342 113686 27398 114486
rect 29642 113686 29698 114486
rect 31942 113686 31998 114486
rect 34242 113686 34298 114486
rect 36542 113686 36598 114486
rect 38842 113686 38898 114486
rect 41142 113686 41198 114486
rect 43442 113686 43498 114486
rect 45742 113686 45798 114486
rect 48042 113686 48098 114486
rect 50342 113686 50398 114486
rect 52642 113686 52698 114486
rect 54942 113686 54998 114486
rect 57242 113686 57298 114486
rect 59542 113686 59598 114486
rect 61842 113686 61898 114486
rect 64142 113686 64198 114486
rect 66442 113686 66498 114486
rect 68742 113686 68798 114486
rect 71042 113686 71098 114486
rect 73342 113686 73398 114486
rect 75642 113686 75698 114486
rect 77942 113686 77998 114486
rect 80242 113686 80298 114486
rect 82542 113686 82598 114486
rect 84842 113686 84898 114486
rect 87142 113686 87198 114486
rect 89442 113686 89498 114486
rect 91742 113686 91798 114486
rect 94042 113686 94098 114486
rect 96342 113686 96398 114486
rect 98642 113686 98698 114486
rect 100942 113686 100998 114486
rect 103242 113686 103298 114486
rect 105542 113686 105598 114486
rect 107842 113686 107898 114486
rect 110142 113686 110198 114486
rect 1674 0 1730 800
rect 4618 0 4674 800
rect 7562 0 7618 800
rect 10506 0 10562 800
rect 13450 0 13506 800
rect 16394 0 16450 800
rect 19338 0 19394 800
rect 22282 0 22338 800
rect 25226 0 25282 800
rect 28170 0 28226 800
rect 31114 0 31170 800
rect 34058 0 34114 800
rect 37002 0 37058 800
rect 39946 0 40002 800
rect 42890 0 42946 800
rect 45834 0 45890 800
rect 48778 0 48834 800
rect 51722 0 51778 800
rect 54666 0 54722 800
rect 57610 0 57666 800
rect 60554 0 60610 800
rect 63498 0 63554 800
rect 66442 0 66498 800
rect 69386 0 69442 800
rect 72330 0 72386 800
rect 75274 0 75330 800
rect 78218 0 78274 800
rect 81162 0 81218 800
rect 84106 0 84162 800
rect 87050 0 87106 800
rect 89994 0 90050 800
rect 92938 0 92994 800
rect 95882 0 95938 800
rect 98826 0 98882 800
rect 101770 0 101826 800
rect 104714 0 104770 800
rect 107658 0 107714 800
rect 110602 0 110658 800
<< obsm2 >>
rect 1676 113630 1986 113778
rect 2154 113630 4286 113778
rect 4454 113630 6586 113778
rect 6754 113630 8886 113778
rect 9054 113630 11186 113778
rect 11354 113630 13486 113778
rect 13654 113630 15786 113778
rect 15954 113630 18086 113778
rect 18254 113630 20386 113778
rect 20554 113630 22686 113778
rect 22854 113630 24986 113778
rect 25154 113630 27286 113778
rect 27454 113630 29586 113778
rect 29754 113630 31886 113778
rect 32054 113630 34186 113778
rect 34354 113630 36486 113778
rect 36654 113630 38786 113778
rect 38954 113630 41086 113778
rect 41254 113630 43386 113778
rect 43554 113630 45686 113778
rect 45854 113630 47986 113778
rect 48154 113630 50286 113778
rect 50454 113630 52586 113778
rect 52754 113630 54886 113778
rect 55054 113630 57186 113778
rect 57354 113630 59486 113778
rect 59654 113630 61786 113778
rect 61954 113630 64086 113778
rect 64254 113630 66386 113778
rect 66554 113630 68686 113778
rect 68854 113630 70986 113778
rect 71154 113630 73286 113778
rect 73454 113630 75586 113778
rect 75754 113630 77886 113778
rect 78054 113630 80186 113778
rect 80354 113630 82486 113778
rect 82654 113630 84786 113778
rect 84954 113630 87086 113778
rect 87254 113630 89386 113778
rect 89554 113630 91686 113778
rect 91854 113630 93986 113778
rect 94154 113630 96286 113778
rect 96454 113630 98586 113778
rect 98754 113630 100886 113778
rect 101054 113630 103186 113778
rect 103354 113630 105486 113778
rect 105654 113630 107786 113778
rect 107954 113630 110086 113778
rect 110254 113630 110932 113778
rect 1676 856 110932 113630
rect 1786 734 4562 856
rect 4730 734 7506 856
rect 7674 734 10450 856
rect 10618 734 13394 856
rect 13562 734 16338 856
rect 16506 734 19282 856
rect 19450 734 22226 856
rect 22394 734 25170 856
rect 25338 734 28114 856
rect 28282 734 31058 856
rect 31226 734 34002 856
rect 34170 734 36946 856
rect 37114 734 39890 856
rect 40058 734 42834 856
rect 43002 734 45778 856
rect 45946 734 48722 856
rect 48890 734 51666 856
rect 51834 734 54610 856
rect 54778 734 57554 856
rect 57722 734 60498 856
rect 60666 734 63442 856
rect 63610 734 66386 856
rect 66554 734 69330 856
rect 69498 734 72274 856
rect 72442 734 75218 856
rect 75386 734 78162 856
rect 78330 734 81106 856
rect 81274 734 84050 856
rect 84218 734 86994 856
rect 87162 734 89938 856
rect 90106 734 92882 856
rect 93050 734 95826 856
rect 95994 734 98770 856
rect 98938 734 101714 856
rect 101882 734 104658 856
rect 104826 734 107602 856
rect 107770 734 110546 856
rect 110714 734 110932 856
<< metal3 >>
rect 111542 111392 112342 111512
rect 111542 108536 112342 108656
rect 111542 105680 112342 105800
rect 111542 102824 112342 102944
rect 111542 99968 112342 100088
rect 111542 97112 112342 97232
rect 111542 94256 112342 94376
rect 111542 91400 112342 91520
rect 111542 88544 112342 88664
rect 111542 85688 112342 85808
rect 111542 82832 112342 82952
rect 111542 79976 112342 80096
rect 111542 77120 112342 77240
rect 111542 74264 112342 74384
rect 111542 71408 112342 71528
rect 111542 68552 112342 68672
rect 111542 65696 112342 65816
rect 111542 62840 112342 62960
rect 111542 59984 112342 60104
rect 111542 57128 112342 57248
rect 111542 54272 112342 54392
rect 111542 51416 112342 51536
rect 111542 48560 112342 48680
rect 111542 45704 112342 45824
rect 111542 42848 112342 42968
rect 111542 39992 112342 40112
rect 111542 37136 112342 37256
rect 111542 34280 112342 34400
rect 111542 31424 112342 31544
rect 111542 28568 112342 28688
rect 111542 25712 112342 25832
rect 111542 22856 112342 22976
rect 111542 20000 112342 20120
rect 111542 17144 112342 17264
rect 111542 14288 112342 14408
rect 111542 11432 112342 11552
rect 111542 8576 112342 8696
rect 111542 5720 112342 5840
rect 111542 2864 112342 2984
<< obsm3 >>
rect 4210 111592 111542 112097
rect 4210 111312 111462 111592
rect 4210 108736 111542 111312
rect 4210 108456 111462 108736
rect 4210 105880 111542 108456
rect 4210 105600 111462 105880
rect 4210 103024 111542 105600
rect 4210 102744 111462 103024
rect 4210 100168 111542 102744
rect 4210 99888 111462 100168
rect 4210 97312 111542 99888
rect 4210 97032 111462 97312
rect 4210 94456 111542 97032
rect 4210 94176 111462 94456
rect 4210 91600 111542 94176
rect 4210 91320 111462 91600
rect 4210 88744 111542 91320
rect 4210 88464 111462 88744
rect 4210 85888 111542 88464
rect 4210 85608 111462 85888
rect 4210 83032 111542 85608
rect 4210 82752 111462 83032
rect 4210 80176 111542 82752
rect 4210 79896 111462 80176
rect 4210 77320 111542 79896
rect 4210 77040 111462 77320
rect 4210 74464 111542 77040
rect 4210 74184 111462 74464
rect 4210 71608 111542 74184
rect 4210 71328 111462 71608
rect 4210 68752 111542 71328
rect 4210 68472 111462 68752
rect 4210 65896 111542 68472
rect 4210 65616 111462 65896
rect 4210 63040 111542 65616
rect 4210 62760 111462 63040
rect 4210 60184 111542 62760
rect 4210 59904 111462 60184
rect 4210 57328 111542 59904
rect 4210 57048 111462 57328
rect 4210 54472 111542 57048
rect 4210 54192 111462 54472
rect 4210 51616 111542 54192
rect 4210 51336 111462 51616
rect 4210 48760 111542 51336
rect 4210 48480 111462 48760
rect 4210 45904 111542 48480
rect 4210 45624 111462 45904
rect 4210 43048 111542 45624
rect 4210 42768 111462 43048
rect 4210 40192 111542 42768
rect 4210 39912 111462 40192
rect 4210 37336 111542 39912
rect 4210 37056 111462 37336
rect 4210 34480 111542 37056
rect 4210 34200 111462 34480
rect 4210 31624 111542 34200
rect 4210 31344 111462 31624
rect 4210 28768 111542 31344
rect 4210 28488 111462 28768
rect 4210 25912 111542 28488
rect 4210 25632 111462 25912
rect 4210 23056 111542 25632
rect 4210 22776 111462 23056
rect 4210 20200 111542 22776
rect 4210 19920 111462 20200
rect 4210 17344 111542 19920
rect 4210 17064 111462 17344
rect 4210 14488 111542 17064
rect 4210 14208 111462 14488
rect 4210 11632 111542 14208
rect 4210 11352 111462 11632
rect 4210 8776 111542 11352
rect 4210 8496 111462 8776
rect 4210 5920 111542 8496
rect 4210 5640 111462 5920
rect 4210 3064 111542 5640
rect 4210 2784 111462 3064
rect 4210 2143 111542 2784
<< metal4 >>
rect 4208 2128 4528 112112
rect 19568 2128 19888 112112
rect 34928 2128 35248 112112
rect 50288 2128 50608 112112
rect 65648 2128 65968 112112
rect 81008 2128 81328 112112
rect 96368 2128 96688 112112
<< obsm4 >>
rect 23059 2483 34848 111893
rect 35328 2483 50208 111893
rect 50688 2483 65568 111893
rect 66048 2483 80928 111893
rect 81408 2483 96288 111893
rect 96768 2483 97829 111893
<< labels >>
rlabel metal3 s 111542 2864 112342 2984 6 i_clk
port 1 nsew signal input
rlabel metal3 s 111542 68552 112342 68672 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 111542 48560 112342 48680 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 111542 14288 112342 14408 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 111542 17144 112342 17264 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 111542 20000 112342 20120 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 111542 22856 112342 22976 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 111542 25712 112342 25832 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 111542 28568 112342 28688 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 111542 31424 112342 31544 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 111542 34280 112342 34400 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 111542 37136 112342 37256 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 111542 39992 112342 40112 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 111542 42848 112342 42968 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 111542 45704 112342 45824 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 111542 51416 112342 51536 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 111542 54272 112342 54392 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 111542 57128 112342 57248 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 111542 59984 112342 60104 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 111542 62840 112342 62960 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 111542 65696 112342 65816 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 111542 71408 112342 71528 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 111542 74264 112342 74384 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 111542 77120 112342 77240 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 111542 79976 112342 80096 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 111542 82832 112342 82952 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 111542 85688 112342 85808 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 111542 88544 112342 88664 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 111542 91400 112342 91520 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 111542 94256 112342 94376 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 111542 97112 112342 97232 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 111542 99968 112342 100088 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 111542 102824 112342 102944 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 111542 105680 112342 105800 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 111542 108536 112342 108656 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 111542 111392 112342 111512 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 111542 5720 112342 5840 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 111542 8576 112342 8696 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 111542 11432 112342 11552 6 i_reg_sclk
port 47 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 i_reset_lock_a
port 48 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 i_reset_lock_b
port 49 nsew signal input
rlabel metal2 s 8942 113686 8998 114486 6 i_tex_in[0]
port 50 nsew signal input
rlabel metal2 s 6642 113686 6698 114486 6 i_tex_in[1]
port 51 nsew signal input
rlabel metal2 s 4342 113686 4398 114486 6 i_tex_in[2]
port 52 nsew signal input
rlabel metal2 s 2042 113686 2098 114486 6 i_tex_in[3]
port 53 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 i_vec_csb
port 54 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 i_vec_mosi
port 55 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 i_vec_sclk
port 56 nsew signal input
rlabel metal2 s 22742 113686 22798 114486 6 o_gpout[0]
port 57 nsew signal output
rlabel metal2 s 20442 113686 20498 114486 6 o_gpout[1]
port 58 nsew signal output
rlabel metal2 s 18142 113686 18198 114486 6 o_gpout[2]
port 59 nsew signal output
rlabel metal2 s 15842 113686 15898 114486 6 o_gpout[3]
port 60 nsew signal output
rlabel metal2 s 13542 113686 13598 114486 6 o_gpout[4]
port 61 nsew signal output
rlabel metal2 s 11242 113686 11298 114486 6 o_gpout[5]
port 62 nsew signal output
rlabel metal2 s 36542 113686 36598 114486 6 o_hsync
port 63 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 o_reset
port 64 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 o_rgb[0]
port 65 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 o_rgb[10]
port 66 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 o_rgb[11]
port 67 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 o_rgb[12]
port 68 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 o_rgb[13]
port 69 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 o_rgb[14]
port 70 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 o_rgb[15]
port 71 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 o_rgb[16]
port 72 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 o_rgb[17]
port 73 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 o_rgb[18]
port 74 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 o_rgb[19]
port 75 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 o_rgb[1]
port 76 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 o_rgb[20]
port 77 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 o_rgb[21]
port 78 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 o_rgb[22]
port 79 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 o_rgb[23]
port 80 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 o_rgb[2]
port 81 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 o_rgb[3]
port 82 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 o_rgb[4]
port 83 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 o_rgb[5]
port 84 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 o_rgb[6]
port 85 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 o_rgb[7]
port 86 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 o_rgb[8]
port 87 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 o_rgb[9]
port 88 nsew signal output
rlabel metal2 s 31942 113686 31998 114486 6 o_tex_csb
port 89 nsew signal output
rlabel metal2 s 29642 113686 29698 114486 6 o_tex_oeb0
port 90 nsew signal output
rlabel metal2 s 27342 113686 27398 114486 6 o_tex_out0
port 91 nsew signal output
rlabel metal2 s 25042 113686 25098 114486 6 o_tex_sclk
port 92 nsew signal output
rlabel metal2 s 34242 113686 34298 114486 6 o_vsync
port 93 nsew signal output
rlabel metal2 s 110142 113686 110198 114486 6 ones[0]
port 94 nsew signal output
rlabel metal2 s 87142 113686 87198 114486 6 ones[10]
port 95 nsew signal output
rlabel metal2 s 84842 113686 84898 114486 6 ones[11]
port 96 nsew signal output
rlabel metal2 s 82542 113686 82598 114486 6 ones[12]
port 97 nsew signal output
rlabel metal2 s 80242 113686 80298 114486 6 ones[13]
port 98 nsew signal output
rlabel metal2 s 77942 113686 77998 114486 6 ones[14]
port 99 nsew signal output
rlabel metal2 s 75642 113686 75698 114486 6 ones[15]
port 100 nsew signal output
rlabel metal2 s 107842 113686 107898 114486 6 ones[1]
port 101 nsew signal output
rlabel metal2 s 105542 113686 105598 114486 6 ones[2]
port 102 nsew signal output
rlabel metal2 s 103242 113686 103298 114486 6 ones[3]
port 103 nsew signal output
rlabel metal2 s 100942 113686 100998 114486 6 ones[4]
port 104 nsew signal output
rlabel metal2 s 98642 113686 98698 114486 6 ones[5]
port 105 nsew signal output
rlabel metal2 s 96342 113686 96398 114486 6 ones[6]
port 106 nsew signal output
rlabel metal2 s 94042 113686 94098 114486 6 ones[7]
port 107 nsew signal output
rlabel metal2 s 91742 113686 91798 114486 6 ones[8]
port 108 nsew signal output
rlabel metal2 s 89442 113686 89498 114486 6 ones[9]
port 109 nsew signal output
rlabel metal4 s 4208 2128 4528 112112 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 112112 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 112112 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 112112 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 112112 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 112112 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 112112 6 vssd1
port 111 nsew ground bidirectional
rlabel metal2 s 73342 113686 73398 114486 6 zeros[0]
port 112 nsew signal output
rlabel metal2 s 50342 113686 50398 114486 6 zeros[10]
port 113 nsew signal output
rlabel metal2 s 48042 113686 48098 114486 6 zeros[11]
port 114 nsew signal output
rlabel metal2 s 45742 113686 45798 114486 6 zeros[12]
port 115 nsew signal output
rlabel metal2 s 43442 113686 43498 114486 6 zeros[13]
port 116 nsew signal output
rlabel metal2 s 41142 113686 41198 114486 6 zeros[14]
port 117 nsew signal output
rlabel metal2 s 38842 113686 38898 114486 6 zeros[15]
port 118 nsew signal output
rlabel metal2 s 71042 113686 71098 114486 6 zeros[1]
port 119 nsew signal output
rlabel metal2 s 68742 113686 68798 114486 6 zeros[2]
port 120 nsew signal output
rlabel metal2 s 66442 113686 66498 114486 6 zeros[3]
port 121 nsew signal output
rlabel metal2 s 64142 113686 64198 114486 6 zeros[4]
port 122 nsew signal output
rlabel metal2 s 61842 113686 61898 114486 6 zeros[5]
port 123 nsew signal output
rlabel metal2 s 59542 113686 59598 114486 6 zeros[6]
port 124 nsew signal output
rlabel metal2 s 57242 113686 57298 114486 6 zeros[7]
port 125 nsew signal output
rlabel metal2 s 54942 113686 54998 114486 6 zeros[8]
port 126 nsew signal output
rlabel metal2 s 52642 113686 52698 114486 6 zeros[9]
port 127 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 112342 114486
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30335970
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_11_01_12_48/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1472938
<< end >>

