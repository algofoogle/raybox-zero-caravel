* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_la_invalid i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_outs_enb i_reg_sclk i_reset_lock_a i_reset_lock_b i_spare_0 i_spare_1 i_tex_in[0]
+ i_tex_in[1] i_tex_in[2] i_tex_in[3] i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1]
+ o_gpout[2] o_gpout[3] o_gpout[4] o_gpout[5] o_hsync o_reset o_rgb[10] o_rgb[11]
+ o_rgb[12] o_rgb[13] o_rgb[14] o_rgb[15] o_rgb[17] o_rgb[18] o_rgb[21] o_rgb[22]
+ o_rgb[23] o_rgb[6] o_rgb[7] o_rgb[9] o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk
+ o_vsync ones[0] ones[11] ones[12] ones[1] ones[2] ones[5] ones[6] ones[7] ones[8]
+ ones[9] vccd1 vssd1 zeros[0] zeros[10] zeros[11] zeros[12] zeros[13] zeros[14] zeros[15]
+ zeros[1] zeros[2] zeros[3] zeros[4] zeros[5] zeros[6] zeros[7] zeros[9] o_rgb[16]
+ ones[10] ones[4] ones[15] ones[3] ones[14] ones[13] o_rgb[8] o_rgb[5] o_rgb[4] o_rgb[3]
+ o_rgb[2] o_rgb[1] o_rgb[0] o_rgb[20] o_rgb[19] zeros[8]
XFILLER_0_59_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18869_ net6695 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20900_ clknet_leaf_32_i_clk net5533 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_21880_ net322 net1784 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20831_ net3628 net5923 vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__nor2_1
X_20762_ _03878_ net8181 _03935_ _03883_ net5448 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20693_ _03874_ _03875_ _03876_ _03877_ net4968 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a32o_1
Xhold7401 rbzero.wall_tracer.stepDistX\[-4\] vssd1 vssd1 vccd1 vccd1 net7928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7412 net3427 vssd1 vssd1 vccd1 vccd1 net7939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7423 net4540 vssd1 vssd1 vccd1 vccd1 net7950 sky130_fd_sc_hd__dlygate4sd3_1
X_20633__362 clknet_1_0__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__inv_2
Xhold7434 rbzero.wall_tracer.trackDistX\[1\] vssd1 vssd1 vccd1 vccd1 net7961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6700 rbzero.tex_g0\[16\] vssd1 vssd1 vccd1 vccd1 net7227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7445 net3846 vssd1 vssd1 vccd1 vccd1 net7972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6711 net2755 vssd1 vssd1 vccd1 vccd1 net7238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7456 rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1 vccd1 net7983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6722 rbzero.tex_g1\[23\] vssd1 vssd1 vccd1 vccd1 net7249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7467 net3834 vssd1 vssd1 vccd1 vccd1 net7994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6733 net2833 vssd1 vssd1 vccd1 vccd1 net7260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7478 rbzero.wall_tracer.trackDistX\[7\] vssd1 vssd1 vccd1 vccd1 net8005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7489 _00515_ vssd1 vssd1 vccd1 vccd1 net8016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6744 rbzero.pov.sclk_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net7271 sky130_fd_sc_hd__dlygate4sd3_1
X_21314_ clknet_leaf_3_i_clk net5167 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6755 _04446_ vssd1 vssd1 vccd1 vccd1 net7282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6766 net2638 vssd1 vssd1 vccd1 vccd1 net7293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6777 _03409_ vssd1 vssd1 vccd1 vccd1 net7304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6788 rbzero.tex_g0\[24\] vssd1 vssd1 vccd1 vccd1 net7315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6799 net2950 vssd1 vssd1 vccd1 vccd1 net7326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 net5253 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
X_21245_ clknet_leaf_11_i_clk net3747 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold351 net5283 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold362 net7523 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 net5656 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_1
Xhold384 net5291 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21176_ clknet_leaf_97_i_clk net2127 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold395 net5255 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20127_ net7595 _03707_ net4477 _03679_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20058_ net41 _03605_ _03140_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o21ai_4
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 net3008 vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 _01270_ vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _01403_ vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ net3517 _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__or2_2
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1073 net6161 vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ net4864 vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__buf_1
Xhold1084 net5530 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 net3898 vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__buf_4
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ net87 _04976_ _04851_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a31o_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _07708_ _07720_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__xor2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _04951_ vssd1 vssd1 vccd1 vccd1 _04952_
+ sky130_fd_sc_hd__mux2_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13501_ _06666_ _06668_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__and3_1
X_10713_ net2593 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__clkbuf_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _07610_ _07651_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__nor2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ net3388 _04861_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ _09311_ _09312_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ _06516_ _06599_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__or3_1
X_10644_ net6828 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16151_ _09123_ _09121_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ net2325 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ net561 net560 _06498_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer7 _06981_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
X_15102_ net5887 _08169_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__nand2_1
X_12314_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _04913_ vssd1 vssd1 vccd1 vccd1 _05500_
+ sky130_fd_sc_hd__mux2_1
X_16082_ net8065 _08128_ _08491_ _09035_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__or4_1
X_13294_ _06351_ _06435_ _06442_ _06454_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__nor4_1
XFILLER_0_106_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15033_ _06121_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19910_ net3261 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
X_12245_ _04967_ _05419_ _05423_ _04818_ _05431_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03510_ _03510_ vssd1 vssd1 vccd1 vccd1 clknet_0__03510_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _05239_ vssd1 vssd1 vccd1 vccd1 _05364_
+ sky130_fd_sc_hd__mux2_1
X_19841_ net3146 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ net51 net6904 _04309_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__mux2_1
X_16984_ _10004_ _10005_ vssd1 vssd1 vccd1 vccd1 _10006_ sky130_fd_sc_hd__nand2_4
XFILLER_0_208_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11058_ net5589 net5634 _04342_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
X_15935_ _09028_ _09029_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__xnor2_2
X_18723_ _02846_ _02872_ _02873_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18654_ net3619 net4423 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__nand2_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _08958_ _08960_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__nand2_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14817_ _07977_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
X_17605_ _01845_ net4659 _10260_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_135_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18585_ _06060_ _09103_ _09774_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a21oi_1
Xtop_ew_algofoogle_120 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_120/HI zeros[9] sky130_fd_sc_hd__conb_1
X_15797_ _08858_ _08891_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_131 vssd1 vssd1 vccd1 vccd1 ones[4] top_ew_algofoogle_131/LO sky130_fd_sc_hd__conb_1
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_142 vssd1 vssd1 vccd1 vccd1 ones[15] top_ew_algofoogle_142/LO sky130_fd_sc_hd__conb_1
X_17536_ _01677_ _01745_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14748_ net7823 vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17467_ _10428_ _01708_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14679_ _07780_ _07783_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ _08308_ _08403_ _09508_ vssd1 vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__or3_1
XFILLER_0_171_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19206_ net5065 _03182_ _03191_ _03189_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__o211a_1
X_17398_ _10414_ _10415_ vssd1 vssd1 vccd1 vccd1 _10416_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19137_ net1238 _03147_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__or2_1
Xhold6007 net1499 vssd1 vssd1 vccd1 vccd1 net6534 sky130_fd_sc_hd__dlygate4sd3_1
X_16349_ _09311_ _09312_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6018 rbzero.spi_registers.new_leak\[1\] vssd1 vssd1 vccd1 vccd1 net6545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6029 net1384 vssd1 vssd1 vccd1 vccd1 net6556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5306 _00599_ vssd1 vssd1 vccd1 vccd1 net5833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5317 rbzero.spi_registers.spi_counter\[0\] vssd1 vssd1 vccd1 vccd1 net5844 sky130_fd_sc_hd__dlygate4sd3_1
X_19068_ net3771 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__clkbuf_1
Xhold5328 _02844_ vssd1 vssd1 vccd1 vccd1 net5855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5339 net3487 vssd1 vssd1 vccd1 vccd1 net5866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4605 rbzero.spi_registers.texadd2\[18\] vssd1 vssd1 vccd1 vccd1 net5132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019_ _02230_ _02231_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4616 net739 vssd1 vssd1 vccd1 vccd1 net5143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4627 _00871_ vssd1 vssd1 vccd1 vccd1 net5154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4638 net907 vssd1 vssd1 vccd1 vccd1 net5165 sky130_fd_sc_hd__dlygate4sd3_1
X_21030_ clknet_leaf_53_i_clk net4227 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4649 rbzero.spi_registers.texadd2\[15\] vssd1 vssd1 vccd1 vccd1 net5176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3904 net8175 vssd1 vssd1 vccd1 vccd1 net4431 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3915 _03624_ vssd1 vssd1 vccd1 vccd1 net4442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3926 net637 vssd1 vssd1 vccd1 vccd1 net4453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3937 _01200_ vssd1 vssd1 vccd1 vccd1 net4464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3948 net1114 vssd1 vssd1 vccd1 vccd1 net4475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21932_ net374 net1175 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21863_ net305 net2672 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20814_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__nor2_1
X_21794_ net236 net2932 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20745_ net834 net4972 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20557__293 clknet_1_0__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__inv_2
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7220 rbzero.wall_hot\[1\] vssd1 vssd1 vccd1 vccd1 net7747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7242 _09085_ vssd1 vssd1 vccd1 vccd1 net7769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7253 rbzero.debug_overlay.playerY\[-4\] vssd1 vssd1 vccd1 vccd1 net7780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6530 net2235 vssd1 vssd1 vccd1 vccd1 net7057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6541 _04114_ vssd1 vssd1 vccd1 vccd1 net7068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7286 _07859_ vssd1 vssd1 vccd1 vccd1 net7813 sky130_fd_sc_hd__buf_2
Xhold6552 net2750 vssd1 vssd1 vccd1 vccd1 net7079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7297 _07916_ vssd1 vssd1 vccd1 vccd1 net7824 sky130_fd_sc_hd__clkbuf_4
Xhold6563 rbzero.tex_g1\[42\] vssd1 vssd1 vccd1 vccd1 net7090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6574 net2113 vssd1 vssd1 vccd1 vccd1 net7101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6585 rbzero.tex_b0\[4\] vssd1 vssd1 vccd1 vccd1 net7112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5840 net1374 vssd1 vssd1 vccd1 vccd1 net6367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6596 net2688 vssd1 vssd1 vccd1 vccd1 net7123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5851 net1441 vssd1 vssd1 vccd1 vccd1 net6378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5862 rbzero.spi_registers.new_texadd\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net6389
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ _04984_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__or2_1
Xhold5873 rbzero.spi_registers.new_texadd\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 net6400
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21228_ clknet_leaf_121_i_clk net3281 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5884 net1429 vssd1 vssd1 vccd1 vccd1 net6411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5895 net1496 vssd1 vssd1 vccd1 vccd1 net6422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold170 net5004 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 net5070 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 net5064 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
X_21159_ clknet_4_1__leaf_i_clk net3698 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13981_ _07105_ _07106_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__nand2_1
X_19813__88 clknet_1_1__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__inv_2
X_15720_ net7836 _08252_ _08254_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_52_i_clk clknet_4_11__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12932_ net4420 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__inv_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15651_ _08688_ _08727_ _08744_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__a21o_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12863_ net5937 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__buf_2
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _07729_ _07733_ _07771_ _07772_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__and4_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _04976_ _05003_ _04828_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18370_ _02551_ _02555_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__xnor2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15582_ _08640_ _08659_ _08675_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__a21o_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _05957_ _05966_ _05965_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_i_clk clknet_4_13__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17321_ _10211_ _10096_ _10220_ _08918_ vssd1 vssd1 vccd1 vccd1 _10340_ sky130_fd_sc_hd__o22ai_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _07033_ _07457_ _07703_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__or3_1
X_11745_ _04910_ _04934_ _04829_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__o21a_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _10181_ _10147_ vssd1 vssd1 vccd1 vccd1 _10271_ sky130_fd_sc_hd__or2b_1
X_14464_ _07592_ _07591_ _07590_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__a21o_1
X_11676_ net3488 _04857_ net3151 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16203_ _08421_ _09294_ _09295_ _08442_ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__a31o_1
X_13415_ _06550_ _06584_ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__or3_4
X_10627_ net2818 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17183_ _10192_ _10202_ vssd1 vssd1 vccd1 vccd1 _10203_ sky130_fd_sc_hd__xnor2_1
X_14395_ _07564_ _07565_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _09112_ _09117_ _09111_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__a21bo_1
X_13346_ _06424_ _06432_ _06426_ _06430_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__and4bb_1
X_10558_ net6922 net2880 _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16065_ _08509_ _08392_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ net8217 _06321_ _06323_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a21oi_2
X_10489_ net6882 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__clkbuf_1
X_15016_ net4183 _08037_ _08034_ _01633_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o211a_1
X_12228_ _04942_ _05402_ _05406_ _04844_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__o311a_1
XFILLER_0_208_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20385__138 clknet_1_1__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__inv_2
X_19824_ net3231 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
X_12159_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _05239_ vssd1 vssd1 vccd1 vccd1 _05347_
+ sky130_fd_sc_hd__mux2_1
Xhold1809 net6897 vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19755_ clknet_1_0__leaf__03506_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__buf_1
XFILLER_0_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16967_ _09663_ _09689_ _09688_ vssd1 vssd1 vccd1 vccd1 _09989_ sky130_fd_sc_hd__a21boi_2
X_18706_ rbzero.wall_tracer.rayAddendY\[2\] rbzero.wall_tracer.rayAddendY\[1\] rbzero.debug_overlay.vplaneY\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15918_ _08397_ _08994_ _09011_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__nand3_1
X_16898_ _09918_ _09919_ vssd1 vssd1 vccd1 vccd1 _09920_ sky130_fd_sc_hd__nor2_1
X_19686_ net6325 net3745 _03468_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15849_ _08529_ _08474_ _08494_ _08277_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__o22a_1
X_18637_ _02793_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18568_ _08103_ _09755_ _02733_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17519_ _08461_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18499_ _02626_ net3494 net4554 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__or3b_2
XFILLER_0_28_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20461_ clknet_1_0__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__buf_1
XFILLER_0_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5103 net1748 vssd1 vssd1 vccd1 vccd1 net5630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5114 _04316_ vssd1 vssd1 vccd1 vccd1 net5641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5125 rbzero.tex_b1\[61\] vssd1 vssd1 vccd1 vccd1 net5652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5136 _04244_ vssd1 vssd1 vccd1 vccd1 net5663 sky130_fd_sc_hd__dlygate4sd3_1
X_22131_ clknet_leaf_52_i_clk net5728 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4402 _01659_ vssd1 vssd1 vccd1 vccd1 net4929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5147 _04372_ vssd1 vssd1 vccd1 vccd1 net5674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5158 _04385_ vssd1 vssd1 vccd1 vccd1 net5685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4413 net604 vssd1 vssd1 vccd1 vccd1 net4940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5169 net3114 vssd1 vssd1 vccd1 vccd1 net5696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4424 rbzero.color_floor\[3\] vssd1 vssd1 vccd1 vccd1 net4951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4435 net620 vssd1 vssd1 vccd1 vccd1 net4962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4446 _01609_ vssd1 vssd1 vccd1 vccd1 net4973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3701 net7854 vssd1 vssd1 vccd1 vccd1 net4228 sky130_fd_sc_hd__dlygate4sd3_1
X_22062_ net504 net2743 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold4457 net658 vssd1 vssd1 vccd1 vccd1 net4984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3712 rbzero.wall_tracer.visualWallDist\[-2\] vssd1 vssd1 vccd1 vccd1 net4239
+ sky130_fd_sc_hd__buf_1
Xhold3723 rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1 vccd1 vccd1 net4250
+ sky130_fd_sc_hd__buf_1
X_21013_ clknet_leaf_62_i_clk net4244 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3734 net1155 vssd1 vssd1 vccd1 vccd1 net4261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4479 _00786_ vssd1 vssd1 vccd1 vccd1 net5006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3745 _00497_ vssd1 vssd1 vccd1 vccd1 net4272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3756 rbzero.debug_overlay.playerY\[-1\] vssd1 vssd1 vccd1 vccd1 net4283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3767 net8124 vssd1 vssd1 vccd1 vccd1 net4294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3778 net3151 vssd1 vssd1 vccd1 vccd1 net4305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3789 _00758_ vssd1 vssd1 vccd1 vccd1 net4316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21915_ net357 net2828 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21846_ net288 net1528 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21777_ clknet_leaf_8_i_clk net1476 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ net4347 _04501_ _04600_ _04718_ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20728_ _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20490__233 clknet_1_0__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__inv_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ _04466_ _04493_ _04499_ _04603_ _04652_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__a32o_4
XFILLER_0_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7050 net3448 vssd1 vssd1 vccd1 vccd1 net7577 sky130_fd_sc_hd__dlygate4sd3_1
X_13200_ net4446 net4828 vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__nor2_1
Xhold7061 rbzero.spi_registers.spi_buffer\[16\] vssd1 vssd1 vccd1 vccd1 net7588 sky130_fd_sc_hd__dlygate4sd3_1
X_14180_ _07314_ _07315_ _07317_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__a21oi_1
Xhold7072 net3584 vssd1 vssd1 vccd1 vccd1 net7599 sky130_fd_sc_hd__dlygate4sd3_1
X_11392_ net3857 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__clkinv_4
Xhold7083 _09749_ vssd1 vssd1 vccd1 vccd1 net7610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7094 net3592 vssd1 vssd1 vccd1 vccd1 net7621 sky130_fd_sc_hd__buf_1
Xhold6360 rbzero.tex_r1\[58\] vssd1 vssd1 vccd1 vccd1 net6887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6371 net2336 vssd1 vssd1 vccd1 vccd1 net6898 sky130_fd_sc_hd__dlygate4sd3_1
X_13131_ net4446 net5952 vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__nor2_1
Xhold6382 rbzero.tex_g1\[56\] vssd1 vssd1 vccd1 vccd1 net6909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6393 net2406 vssd1 vssd1 vccd1 vccd1 net6920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5670 net1130 vssd1 vssd1 vccd1 vccd1 net6197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5681 _03482_ vssd1 vssd1 vccd1 vccd1 net6208 sky130_fd_sc_hd__dlygate4sd3_1
X_13062_ _06163_ _06235_ _06237_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5692 net1185 vssd1 vssd1 vccd1 vccd1 net6219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12013_ _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__inv_2
X_17870_ _02104_ _02106_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__and2_1
Xhold4980 net1135 vssd1 vssd1 vccd1 vccd1 net5507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4991 net1550 vssd1 vssd1 vccd1 vccd1 net5518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ net4634 _09846_ _09847_ vssd1 vssd1 vccd1 vccd1 _09848_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_206_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19798__76 clknet_1_0__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__05847_ clknet_0__05847_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05847_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19540_ net6613 net1622 _03388_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__mux2_1
X_16752_ _09103_ _09784_ vssd1 vssd1 vccd1 vccd1 _09786_ sky130_fd_sc_hd__or2_1
X_13964_ _07134_ _07132_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__nor2_2
X_15703_ _08787_ _08791_ _08790_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__a21bo_1
X_12915_ net4777 net4674 _06088_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__or4_1
XFILLER_0_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16683_ net967 _09741_ _09742_ rbzero.wall_tracer.visualWallDist\[-9\] vssd1 vssd1
+ vccd1 vccd1 _00501_ sky130_fd_sc_hd__a22o_1
X_19471_ net1426 net6003 _03345_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__mux2_1
X_13895_ _07064_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15634_ _08210_ _08457_ _08663_ _08662_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__or4b_1
X_18422_ _02598_ _02603_ _02526_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12846_ _05961_ _05962_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__nand2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ net4733 _02528_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__or2_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15565_ _08631_ _08633_ _08632_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__a21o_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__xor2_4
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _08326_ _09403_ vssd1 vssd1 vccd1 vccd1 _10323_ sky130_fd_sc_hd__nor2_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _07666_ _07686_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_1
X_11728_ _04915_ _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18284_ net6454 net3816 _02477_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
X_15496_ _08588_ _08590_ vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _10004_ _10254_ _10129_ vssd1 vssd1 vccd1 vccd1 _10255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14447_ _07033_ _07391_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__nor2_1
X_11659_ _04821_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17166_ _08408_ _08409_ vssd1 vssd1 vccd1 vccd1 _10186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14378_ _07536_ _07547_ _07548_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold906 net6431 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ _09209_ net3420 vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__xnor2_1
Xhold917 net6379 vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _06499_ _06461_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__nand2_1
Xhold928 _01002_ vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ _10114_ _10116_ vssd1 vssd1 vccd1 vccd1 _10118_ sky130_fd_sc_hd__nand2_1
Xhold939 net6451 vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _09140_ _09141_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3008 net4773 vssd1 vssd1 vccd1 vccd1 net3535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3019 net5905 vssd1 vssd1 vccd1 vccd1 net3546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2307 _01029_ vssd1 vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2318 net2682 vssd1 vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2329 _01044_ vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1606 _01587_ vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1617 net6964 vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 net7298 vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ _02234_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__nor2_1
Xhold1639 _01025_ vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
X_19738_ net3823 net7649 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ net6504 net4074 _03457_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
X_21700_ clknet_leaf_115_i_clk net4365 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21631_ clknet_leaf_129_i_clk net3258 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21562_ net196 net2529 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21493_ clknet_leaf_9_i_clk net1772 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4210 net4253 vssd1 vssd1 vccd1 vccd1 net4737 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4221 net4052 vssd1 vssd1 vccd1 vccd1 net4748 sky130_fd_sc_hd__clkbuf_4
X_22114_ clknet_leaf_54_i_clk net4986 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4232 _00428_ vssd1 vssd1 vccd1 vccd1 net4759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4254 _06160_ vssd1 vssd1 vccd1 vccd1 net4781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4265 _02622_ vssd1 vssd1 vccd1 vccd1 net4792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3520 rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 net4047 sky130_fd_sc_hd__dlygate4sd3_1
X_22045_ net487 net2305 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold4276 net674 vssd1 vssd1 vccd1 vccd1 net4803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3531 _05059_ vssd1 vssd1 vccd1 vccd1 net4058 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3542 _00458_ vssd1 vssd1 vccd1 vccd1 net4069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4287 net5894 vssd1 vssd1 vccd1 vccd1 net4814 sky130_fd_sc_hd__clkbuf_2
Xhold3553 net5969 vssd1 vssd1 vccd1 vccd1 net4080 sky130_fd_sc_hd__buf_4
Xhold4298 net1941 vssd1 vssd1 vccd1 vccd1 net4825 sky130_fd_sc_hd__buf_1
Xhold3564 net7715 vssd1 vssd1 vccd1 vccd1 net4091 sky130_fd_sc_hd__buf_2
Xhold2830 _04162_ vssd1 vssd1 vccd1 vccd1 net3357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3575 net3969 vssd1 vssd1 vccd1 vccd1 net4102 sky130_fd_sc_hd__clkbuf_4
Xhold3586 _03800_ vssd1 vssd1 vccd1 vccd1 net4113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2841 _03380_ vssd1 vssd1 vccd1 vccd1 net3368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 net4680 vssd1 vssd1 vccd1 vccd1 net3379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3597 _09720_ vssd1 vssd1 vccd1 vccd1 net4124 sky130_fd_sc_hd__buf_2
Xhold2863 net4456 vssd1 vssd1 vccd1 vccd1 net3390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2874 rbzero.spi_registers.spi_buffer\[8\] vssd1 vssd1 vccd1 vccd1 net3401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2885 _03061_ vssd1 vssd1 vccd1 vccd1 net3412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2896 net4360 vssd1 vssd1 vccd1 vccd1 net3423 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10961_ net7230 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12700_ net31 net30 net32 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a21o_1
X_13680_ _06828_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10892_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ net27 net26 _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and3_1
X_21829_ net271 net2335 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15350_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1 vccd1 vccd1 _08445_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12562_ reg_gpout\[1\] clknet_1_0__leaf__05742_ _05054_ vssd1 vssd1 vccd1 vccd1 _05743_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14301_ _07240_ _07326_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11513_ net3642 _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__or2_1
X_15281_ _08374_ _08375_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ net7716 vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__clkbuf_1
X_17020_ _09373_ _09354_ vssd1 vssd1 vccd1 vccd1 _10041_ sky130_fd_sc_hd__nand2_1
X_14232_ _07033_ _07232_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__or2_1
X_11444_ _04554_ _04555_ rbzero.spi_registers.texadd3\[3\] vssd1 vssd1 vccd1 vccd1
+ _04636_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14163_ _07239_ _07322_ _07333_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11375_ _04555_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__clkbuf_4
Xhold6190 net1840 vssd1 vssd1 vccd1 vccd1 net6717 sky130_fd_sc_hd__dlygate4sd3_1
X_13114_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
X_14094_ _07256_ _07264_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__xor2_1
X_18971_ net2829 net7465 net2874 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _06173_ _06178_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__nor2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _01966_ _02144_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17853_ _02072_ _02090_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16804_ _09826_ _09824_ net4631 vssd1 vssd1 vccd1 vccd1 _09832_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_156_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17784_ _10327_ _10346_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__nor2_1
X_14996_ net4142 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
X_19523_ net4016 net5535 net3086 vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ _06855_ _06859_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__or2b_1
X_16735_ _09770_ _09771_ vssd1 vssd1 vccd1 vccd1 _09772_ sky130_fd_sc_hd__xor2_1
XFILLER_0_205_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20497__239 clknet_1_0__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__inv_2
XFILLER_0_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19454_ net1851 _03334_ net5563 _03339_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16666_ net4303 _09737_ _09740_ _07947_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13878_ _07042_ _07048_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15617_ _08180_ _08245_ _08709_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__and3_1
X_18405_ net4698 net4733 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__and2_1
X_12829_ _05952_ _05955_ _05950_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16597_ _09539_ _09554_ _09686_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__a21bo_1
X_19385_ net5197 _03283_ _03295_ _03288_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15548_ _08283_ _08269_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__xnor2_4
X_18336_ _02524_ _08038_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__nor2_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7808 net4523 vssd1 vssd1 vccd1 vccd1 net8335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7819 rbzero.texu_hot\[2\] vssd1 vssd1 vccd1 vccd1 net8346 sky130_fd_sc_hd__dlygate4sd3_1
X_18267_ net4028 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__clkbuf_1
X_15479_ _08374_ net4877 _08573_ _08366_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17218_ _10111_ _10112_ vssd1 vssd1 vccd1 vccd1 _10238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18198_ _02418_ net3811 _02393_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03856_ clknet_0__03856_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03856_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold703 net6356 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ _10167_ _10168_ vssd1 vssd1 vccd1 vccd1 _10169_ sky130_fd_sc_hd__xnor2_1
Xhold714 net6298 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold725 net5801 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 net6282 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 _01351_ vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 net5523 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
X_20160_ net3505 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold769 _03437_ vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20091_ net4901 _03485_ _03662_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a211o_1
Xhold2104 rbzero.tex_b1\[31\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 _04082_ vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2126 _01428_ vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2137 net7074 vssd1 vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1403 net7026 vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 _01062_ vssd1 vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _04254_ vssd1 vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 net4824 vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 net6767 vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1436 _01425_ vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _04312_ vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1458 net6783 vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _01464_ vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20993_ clknet_leaf_112_i_clk net4136 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21614_ clknet_leaf_97_i_clk net2809 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21545_ net179 net2894 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21476_ clknet_leaf_18_i_clk net4837 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20427_ clknet_1_0__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__buf_1
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ net7246 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4040 net3755 vssd1 vssd1 vccd1 vccd1 net4567 sky130_fd_sc_hd__clkbuf_2
Xhold4051 _00423_ vssd1 vssd1 vccd1 vccd1 net4578 sky130_fd_sc_hd__dlygate4sd3_1
X_11091_ net7385 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
Xhold4062 net3806 vssd1 vssd1 vccd1 vccd1 net4589 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4073 _04011_ vssd1 vssd1 vccd1 vccd1 net4600 sky130_fd_sc_hd__dlygate4sd3_1
X_20289_ net6376 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4084 net8457 vssd1 vssd1 vccd1 vccd1 net4611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4095 net3830 vssd1 vssd1 vccd1 vccd1 net4622 sky130_fd_sc_hd__clkbuf_2
Xhold3350 net3862 vssd1 vssd1 vccd1 vccd1 net3877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3361 net3797 vssd1 vssd1 vccd1 vccd1 net3888 sky130_fd_sc_hd__clkbuf_2
X_22028_ net470 net2819 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3372 net1622 vssd1 vssd1 vccd1 vccd1 net3899 sky130_fd_sc_hd__buf_1
XFILLER_0_175_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3383 _02974_ vssd1 vssd1 vccd1 vccd1 net3910 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3394 net7647 vssd1 vssd1 vccd1 vccd1 net3921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2660 _03541_ vssd1 vssd1 vccd1 vccd1 net3187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2671 rbzero.pov.ss_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net3198 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _07966_ _07978_ _07913_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__mux2_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold63 net5990 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2682 _00677_ vssd1 vssd1 vccd1 vccd1 net3209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 net4937 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold85 net4955 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2693 net7501 vssd1 vssd1 vccd1 vccd1 net3220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 net6025 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _06708_ _06832_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__nor2_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1970 _04046_ vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1981 _01089_ vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14781_ _07943_ _07945_ _07934_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__mux2_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1992 _04190_ vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ net4138 _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__nor2_1
X_16520_ _09607_ _09608_ vssd1 vssd1 vccd1 vccd1 _09610_ sky130_fd_sc_hd__and2_1
X_13732_ _06872_ _06880_ _06881_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__or3_1
X_10944_ net7318 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _09540_ _09541_ _08905_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_196_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ _06831_ _06833_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__xnor2_1
X_10875_ net2886 net7355 _04253_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__mux2_1
X_15402_ _08418_ _08458_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__nor2_2
XFILLER_0_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ net21 net20 net4156 _05746_ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__o41a_2
X_19170_ net5093 _03168_ _03171_ _03160_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16382_ _08611_ _09472_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__nor2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13594_ _06762_ _06763_ _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nand3_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18121_ net3847 net4415 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__nor2_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ net3599 _08119_ _08137_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__o21a_2
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _05708_ _05724_ _05725_ _05718_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18052_ _02284_ _02287_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__xnor2_1
X_15264_ _08355_ _08358_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__nand2_1
X_12476_ net5 net6 net7 vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17003_ _09907_ _09925_ _09923_ vssd1 vssd1 vccd1 vccd1 _10024_ sky130_fd_sc_hd__a21o_1
X_14215_ _06696_ _07327_ _07323_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__o21ai_1
XANTENNA_5 _05630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _04503_ _04534_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15195_ _08133_ _08289_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__nand2_1
X_14146_ _07313_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ rbzero.spi_registers.texadd0\[14\] _04545_ _04548_ _04549_ vssd1 vssd1 vccd1
+ vccd1 _04550_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14077_ _07209_ _07219_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__or2b_1
X_18954_ net6744 net5750 _03036_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
X_11289_ net4083 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__inv_2
X_17905_ _01968_ _02042_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a21oi_2
X_13028_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__inv_2
X_18885_ net6247 net2079 _03003_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _02004_ _02001_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__or2b_1
XFILLER_0_207_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer17 net540 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17767_ _01818_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__nand2_1
Xrebuffer28 _06681_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_1
XFILLER_0_89_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14979_ _08087_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer39 _06988_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_2
X_19506_ net1635 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16718_ net4034 _09102_ _09755_ vssd1 vssd1 vccd1 vccd1 _09756_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17698_ _01935_ _01936_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19437_ net3549 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16649_ _04466_ _04664_ _05184_ net4133 vssd1 vssd1 vccd1 vccd1 _09730_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ net5009 _03283_ _03286_ _03275_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__o211a_1
Xhold7605 net1048 vssd1 vssd1 vccd1 vccd1 net8132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _09735_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__clkbuf_4
Xhold7616 rbzero.floor_leak\[3\] vssd1 vssd1 vccd1 vccd1 net8143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7627 _00496_ vssd1 vssd1 vccd1 vccd1 net8154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19299_ net5117 _03236_ _03245_ _03246_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__o211a_1
Xhold7638 rbzero.map_overlay.i_mapdy\[4\] vssd1 vssd1 vccd1 vccd1 net8165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6904 net2826 vssd1 vssd1 vccd1 vccd1 net7431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6915 rbzero.pov.spi_buffer\[22\] vssd1 vssd1 vccd1 vccd1 net7442 sky130_fd_sc_hd__dlygate4sd3_1
X_21330_ clknet_leaf_8_i_clk net5390 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6926 net3134 vssd1 vssd1 vccd1 vccd1 net7453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6937 rbzero.pov.ready_buffer\[55\] vssd1 vssd1 vccd1 vccd1 net7464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6948 net2066 vssd1 vssd1 vccd1 vccd1 net7475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6959 net3107 vssd1 vssd1 vccd1 vccd1 net7486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold500 net4464 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
X_21261_ clknet_leaf_23_i_clk net3853 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold511 net8208 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold522 net4269 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold533 net4468 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
X_20212_ net4591 _03743_ _03766_ _03765_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold544 _01293_ vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
X_21192_ clknet_leaf_129_i_clk net3082 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold555 _01383_ vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 net6123 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _00685_ vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 net6194 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20143_ _03709_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 _01480_ vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20074_ net4344 _03660_ net3415 _03628_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__o211a_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 net6610 vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _00926_ vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 net5631 vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 _01045_ vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1244 _03446_ vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 net6722 vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 net4333 vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1277 net5537 vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _03518_ vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _01042_ vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ clknet_leaf_42_i_clk net3989 vssd1 vssd1 vccd1 vccd1 rbzero.wall_hot\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ net7224 net6277 _04138_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ net2947 net7287 _04105_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12330_ _04991_ _05507_ _05515_ _04821_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a31o_1
X_21528_ clknet_leaf_124_i_clk net5282 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20610__341 clknet_1_1__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__inv_2
X_12261_ _04955_ _05443_ _05445_ _05447_ _04824_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21459_ clknet_leaf_42_i_clk net1999 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14000_ _07122_ _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__xnor2_1
X_11212_ net6852 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12192_ reg_rgb\[14\] _05379_ _05054_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__mux2_2
X_11143_ net6806 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__clkbuf_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__clkbuf_4
X_11074_ net6130 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
X_15951_ _09043_ _09045_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3180 net7672 vssd1 vssd1 vccd1 vccd1 net3707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3191 net7931 vssd1 vssd1 vccd1 vccd1 net3718 sky130_fd_sc_hd__dlygate4sd3_1
X_14902_ net4547 _08034_ _08036_ net3847 net8238 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__o221a_1
X_15882_ _08925_ _08931_ _08974_ _08976_ _08895_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__o2111a_1
X_18670_ net8093 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2490 _00718_ vssd1 vssd1 vccd1 vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _01748_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__xnor2_1
X_14833_ net4435 _07991_ _07976_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__mux2_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03859_ clknet_0__03859_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03859_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17552_ _01791_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__xnor2_1
X_14764_ _07930_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__clkbuf_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _05164_ _05113_ _05102_ net3538 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _09475_ _09592_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__xor2_1
X_13715_ _06780_ _06782_ _06781_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21o_1
X_17483_ _10266_ _01724_ _10376_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a21o_1
X_10927_ net6074 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ net7813 net7811 _07865_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19222_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__buf_2
X_16434_ _08246_ _08430_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13646_ _06721_ _06673_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__nor2_1
X_10858_ net50 net2503 _04171_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ net4357 _03144_ net837 _03160_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__o211a_1
X_16365_ net7779 _09456_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__nor2_1
X_13577_ _06731_ _06740_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__xnor2_1
X_10789_ net2408 net6456 _04205_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__clkbuf_4
X_18104_ net3787 net4539 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12528_ net54 _05698_ _05708_ net15 vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a31o_1
X_16296_ _09379_ _09387_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__xor2_2
X_19084_ net2182 net6792 _09725_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15247_ _08322_ _08341_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__nor2_1
X_18035_ _02200_ _02214_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12459_ net7 net6 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4809 net913 vssd1 vssd1 vccd1 vccd1 net5336 sky130_fd_sc_hd__dlygate4sd3_1
X_15178_ _08270_ _08272_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ _07200_ _07230_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19986_ net3306 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18937_ _02992_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18868_ net1682 net6693 _02993_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _02055_ _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__nand2_1
X_18799_ _04490_ _02942_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20830_ net3628 net5923 _01633_ _04476_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20761_ _03934_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20692_ _03109_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_175_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7402 net4788 vssd1 vssd1 vccd1 vccd1 net7929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7413 rbzero.wall_tracer.stepDistY\[-4\] vssd1 vssd1 vccd1 vccd1 net7940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7424 rbzero.wall_tracer.trackDistY\[-7\] vssd1 vssd1 vccd1 vccd1 net7951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7435 net4588 vssd1 vssd1 vccd1 vccd1 net7962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6701 net2017 vssd1 vssd1 vccd1 vccd1 net7228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7446 rbzero.wall_tracer.trackDistX\[8\] vssd1 vssd1 vccd1 vccd1 net7973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6712 rbzero.tex_b1\[55\] vssd1 vssd1 vccd1 vccd1 net7239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7457 net3750 vssd1 vssd1 vccd1 vccd1 net7984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6723 net2651 vssd1 vssd1 vccd1 vccd1 net7250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7468 rbzero.wall_tracer.trackDistX\[-1\] vssd1 vssd1 vccd1 vccd1 net7995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6734 rbzero.tex_g1\[52\] vssd1 vssd1 vccd1 vccd1 net7261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7479 net4722 vssd1 vssd1 vccd1 vccd1 net8006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6745 net3305 vssd1 vssd1 vccd1 vccd1 net7272 sky130_fd_sc_hd__dlygate4sd3_1
X_21313_ clknet_leaf_6_i_clk net5151 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6756 net2912 vssd1 vssd1 vccd1 vccd1 net7283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6767 rbzero.tex_r1\[34\] vssd1 vssd1 vccd1 vccd1 net7294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6778 rbzero.tex_b1\[19\] vssd1 vssd1 vccd1 vccd1 net7305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6789 net2300 vssd1 vssd1 vccd1 vccd1 net7316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold330 net5301 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
X_21244_ clknet_leaf_11_i_clk net3840 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold341 net5331 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 net5285 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _03131_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 net5658 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21175_ clknet_leaf_97_i_clk net2163 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold385 net5293 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold396 net5257 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
X_20126_ rbzero.debug_overlay.facingX\[-8\] _03711_ vssd1 vssd1 vccd1 vccd1 _03713_
+ sky130_fd_sc_hd__or2_1
X_20057_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__clkbuf_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1030 _01255_ vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _03592_ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 net6660 vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 net6079 vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 _00594_ vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 net5532 vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ net4271 net4335 net4259 vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__nor3_1
Xhold1096 _03389_ vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__buf_4
XFILLER_0_178_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ clknet_leaf_65_i_clk _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _06493_ _06669_ _06670_ _06557_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ net7252 net5991 _04160_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _07624_ _07649_ _07650_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__a21oi_2
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _04022_ _04860_ _04863_ net4132 _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13431_ _06600_ _06601_ _06492_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643_ net6826 net2950 _04127_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ _09222_ _09242_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__xor2_2
X_13362_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__buf_6
XFILLER_0_134_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10574_ net6554 net6967 _04086_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer8 _07071_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_2
X_15101_ net5887 _08169_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__or2_2
X_12313_ _04818_ _05473_ _05481_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ net8041 _08128_ _08491_ _09174_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__or4_1
X_13293_ _06455_ _06459_ _06461_ _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15032_ _08126_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__clkbuf_4
X_12244_ _05213_ _05426_ _05430_ _04825_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19840_ net3145 net3111 _03528_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12175_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _05239_ vssd1 vssd1 vccd1 vccd1 _05363_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11126_ net6269 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
X_16983_ _09707_ _10003_ vssd1 vssd1 vccd1 vccd1 _10005_ sky130_fd_sc_hd__or2_1
X_18722_ _02872_ _02873_ _02846_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a21oi_1
X_11057_ net1956 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
X_15934_ _08417_ _08403_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18653_ net3575 _05164_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__xor2_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _08942_ _08959_ vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__xor2_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _06058_ _01736_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14816_ net3777 _07975_ _07976_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18584_ net4050 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
X_15796_ _08859_ _08890_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__and2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_110 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_110/HI o_rgb[21]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_121 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_121/HI zeros[10]
+ sky130_fd_sc_hd__conb_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_132 vssd1 vssd1 vccd1 vccd1 ones[5] top_ew_algofoogle_132/LO sky130_fd_sc_hd__conb_1
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17535_ _01758_ _01775_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__xnor2_1
X_11959_ rbzero.debug_overlay.facingY\[-6\] _05102_ _05090_ rbzero.debug_overlay.facingY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a22o_1
X_14747_ net7785 _07913_ _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__xor2_1
X_14678_ _07779_ _07655_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__xnor2_2
X_20617__347 clknet_1_1__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__inv_2
X_19205_ net6301 _03183_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16417_ _08306_ _08418_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__or2_1
X_13629_ _06794_ _06799_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__xnor2_1
X_17397_ _10187_ _10317_ _10319_ vssd1 vssd1 vccd1 vccd1 _10415_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19136_ net4420 _03145_ net1204 _03149_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__o211a_1
Xhold6008 _04398_ vssd1 vssd1 vccd1 vccd1 net6535 sky130_fd_sc_hd__dlygate4sd3_1
X_16348_ _09370_ _09439_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6019 net1643 vssd1 vssd1 vccd1 vccd1 net6546 sky130_fd_sc_hd__dlygate4sd3_1
X_16279_ _09258_ _09268_ _09266_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__a21o_1
X_19067_ _02472_ net3770 _03104_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
Xhold5307 rbzero.pov.ready_buffer\[61\] vssd1 vssd1 vccd1 vccd1 net5834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5318 net2198 vssd1 vssd1 vccd1 vccd1 net5845 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5329 net3753 vssd1 vssd1 vccd1 vccd1 net5856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4606 net773 vssd1 vssd1 vccd1 vccd1 net5133 sky130_fd_sc_hd__dlygate4sd3_1
X_18018_ _02150_ _02153_ _02236_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4617 rbzero.spi_registers.texadd1\[12\] vssd1 vssd1 vccd1 vccd1 net5144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4628 net786 vssd1 vssd1 vccd1 vccd1 net5155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4639 _00801_ vssd1 vssd1 vccd1 vccd1 net5166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3905 _00770_ vssd1 vssd1 vccd1 vccd1 net4432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3916 _03625_ vssd1 vssd1 vccd1 vccd1 net4443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3927 rbzero.pov.ready_buffer\[70\] vssd1 vssd1 vccd1 vccd1 net4454 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3938 net1027 vssd1 vssd1 vccd1 vccd1 net4465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19969_ net6327 net1869 net2312 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__mux2_1
X_20362__117 clknet_1_0__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__inv_2
X_21931_ net373 net3251 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21862_ net304 net2717 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20813_ net5739 _03877_ _03874_ _03978_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_188_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21793_ net235 net2705 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20744_ net834 net4972 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7210 rbzero.debug_overlay.vplaneX\[-9\] vssd1 vssd1 vccd1 vccd1 net7737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7221 rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 net7748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7243 rbzero.debug_overlay.playerX\[-2\] vssd1 vssd1 vccd1 vccd1 net7770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7254 net3317 vssd1 vssd1 vccd1 vccd1 net7781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6520 net2126 vssd1 vssd1 vccd1 vccd1 net7047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6531 rbzero.tex_b0\[37\] vssd1 vssd1 vccd1 vccd1 net7058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6542 net2328 vssd1 vssd1 vccd1 vccd1 net7069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7287 rbzero.wall_tracer.stepDistX\[8\] vssd1 vssd1 vccd1 vccd1 net7814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6553 _04198_ vssd1 vssd1 vccd1 vccd1 net7080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7298 _07957_ vssd1 vssd1 vccd1 vccd1 net7825 sky130_fd_sc_hd__buf_1
Xhold6564 net2432 vssd1 vssd1 vccd1 vccd1 net7091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5830 net1230 vssd1 vssd1 vccd1 vccd1 net6357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6575 rbzero.tex_r0\[60\] vssd1 vssd1 vccd1 vccd1 net7102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6586 net2164 vssd1 vssd1 vccd1 vccd1 net7113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5841 _03436_ vssd1 vssd1 vccd1 vccd1 net6368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6597 rbzero.tex_b0\[19\] vssd1 vssd1 vccd1 vccd1 net7124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5852 rbzero.spi_registers.new_texadd\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net6379
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5863 net1419 vssd1 vssd1 vccd1 vccd1 net6390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5874 net1331 vssd1 vssd1 vccd1 vccd1 net6401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5885 rbzero.pov.spi_buffer\[4\] vssd1 vssd1 vccd1 vccd1 net6412 sky130_fd_sc_hd__dlygate4sd3_1
X_21227_ clknet_leaf_121_i_clk net1705 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold160 net5012 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 net5006 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5896 _03474_ vssd1 vssd1 vccd1 vccd1 net6423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 net5040 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 net5066 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
X_21158_ clknet_leaf_2_i_clk net5802 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20109_ _03483_ _03698_ _03661_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a21o_1
X_13980_ _07116_ _07103_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__or2b_1
X_21089_ clknet_leaf_46_i_clk net1243 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__05794_ clknet_0__05794_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05794_
+ sky130_fd_sc_hd__clkbuf_16
X_12931_ net3964 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__clkbuf_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15650_ _08688_ _08727_ _08744_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__nand3_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ net4642 _06033_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nor2_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11813_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _04978_ vssd1 vssd1 vccd1 vccd1 _05003_
+ sky130_fd_sc_hd__mux2_1
X_14601_ _07706_ _07721_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__xor2_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _08640_ _08659_ _08675_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _05949_ _05956_ _05960_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__or4_4
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _08918_ _10211_ _10096_ _10220_ vssd1 vssd1 vccd1 vccd1 _10339_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _07284_ _07457_ _07701_ _07702_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__o31a_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _04933_ vssd1 vssd1 vccd1 vccd1 _04934_
+ sky130_fd_sc_hd__mux2_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _10021_ _10249_ vssd1 vssd1 vccd1 vccd1 _10270_ sky130_fd_sc_hd__nand2_1
X_14463_ _07592_ _07590_ _07591_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__nand3_1
XFILLER_0_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ _04859_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13414_ net561 net560 _06459_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a21oi_1
X_16202_ _08024_ net75 vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__nand2_1
X_10626_ net7469 net2817 _04116_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__mux2_1
X_17182_ _10199_ _10201_ vssd1 vssd1 vccd1 vccd1 _10202_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14394_ _07284_ _07198_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__nor2_1
X_16133_ _08611_ _09225_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13345_ _06503_ _06511_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__nor3_4
XFILLER_0_148_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ net2768 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16064_ _09156_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__nand2_1
X_13276_ _06327_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__xor2_4
X_10488_ net2229 net6880 _04042_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__mux2_1
X_15015_ net4182 vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__buf_4
X_12227_ _04955_ _05409_ _05413_ _04824_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19823_ net3351 net7554 _03517_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__mux2_1
X_12158_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _05239_ vssd1 vssd1 vccd1 vccd1 _05346_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11109_ net2578 net6637 _04375_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16966_ _09986_ _09987_ vssd1 vssd1 vccd1 vccd1 _09988_ sky130_fd_sc_hd__or2_2
X_12089_ _05276_ _05277_ _04988_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__o21a_1
X_18705_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__or2_1
X_15917_ _08397_ _08994_ _09011_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19685_ net1490 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__clkbuf_1
X_16897_ _09917_ _09914_ vssd1 vssd1 vccd1 vccd1 _09919_ sky130_fd_sc_hd__and2b_1
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ net3677 rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _02794_
+ sky130_fd_sc_hd__and2_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _08329_ _08458_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18567_ _06104_ net7713 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15779_ _08862_ _08867_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17518_ _10409_ _10410_ _10412_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18498_ _02673_ _02674_ _02656_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17449_ _01681_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19119_ net3374 vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5104 _04173_ vssd1 vssd1 vccd1 vccd1 net5631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5115 net656 vssd1 vssd1 vccd1 vccd1 net5642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5126 net2134 vssd1 vssd1 vccd1 vccd1 net5653 sky130_fd_sc_hd__dlygate4sd3_1
X_22130_ clknet_leaf_53_i_clk net5524 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold5137 net2463 vssd1 vssd1 vccd1 vccd1 net5664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5148 net2307 vssd1 vssd1 vccd1 vccd1 net5675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4403 net594 vssd1 vssd1 vccd1 vccd1 net4930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5159 net2704 vssd1 vssd1 vccd1 vccd1 net5686 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__05688_ clknet_0__05688_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05688_
+ sky130_fd_sc_hd__clkbuf_16
Xhold4414 _01655_ vssd1 vssd1 vccd1 vccd1 net4941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4425 net606 vssd1 vssd1 vccd1 vccd1 net4952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22061_ net503 net2344 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold4436 rbzero.color_sky\[2\] vssd1 vssd1 vccd1 vccd1 net4963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4447 net649 vssd1 vssd1 vccd1 vccd1 net4974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3702 net7856 vssd1 vssd1 vccd1 vccd1 net4229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3713 net8019 vssd1 vssd1 vccd1 vccd1 net4240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4458 _01601_ vssd1 vssd1 vccd1 vccd1 net4985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3724 net8080 vssd1 vssd1 vccd1 vccd1 net4251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4469 rbzero.pov.ready vssd1 vssd1 vccd1 vccd1 net4996 sky130_fd_sc_hd__dlygate4sd3_1
X_21012_ clknet_leaf_62_i_clk net4289 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3735 rbzero.wall_tracer.visualWallDist\[4\] vssd1 vssd1 vccd1 vccd1 net4262 sky130_fd_sc_hd__buf_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3746 net1586 vssd1 vssd1 vccd1 vccd1 net4273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3757 net4188 vssd1 vssd1 vccd1 vccd1 net4284 sky130_fd_sc_hd__buf_1
Xhold3768 net897 vssd1 vssd1 vccd1 vccd1 net4295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3779 net8156 vssd1 vssd1 vccd1 vccd1 net4306 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21914_ net356 net2293 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21845_ net287 net2255 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21776_ clknet_leaf_12_i_clk net1324 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20727_ net1120 net5252 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _04466_ _04601_ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7040 net2396 vssd1 vssd1 vccd1 vccd1 net7567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7051 rbzero.spi_registers.spi_buffer\[20\] vssd1 vssd1 vccd1 vccd1 net7578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7062 net3556 vssd1 vssd1 vccd1 vccd1 net7589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7073 rbzero.spi_registers.spi_buffer\[22\] vssd1 vssd1 vccd1 vccd1 net7600 sky130_fd_sc_hd__dlygate4sd3_1
X_11391_ _04577_ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7084 net3649 vssd1 vssd1 vccd1 vccd1 net7611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6350 rbzero.pov.ready_buffer\[39\] vssd1 vssd1 vccd1 vccd1 net6877 sky130_fd_sc_hd__dlygate4sd3_1
X_13130_ net4446 net4828 vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__and2_1
Xhold6361 net2297 vssd1 vssd1 vccd1 vccd1 net6888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6372 _04095_ vssd1 vssd1 vccd1 vccd1 net6899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6383 net2700 vssd1 vssd1 vccd1 vccd1 net6910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold6394 rbzero.tex_r1\[12\] vssd1 vssd1 vccd1 vccd1 net6921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5660 net1142 vssd1 vssd1 vccd1 vccd1 net6187 sky130_fd_sc_hd__dlygate4sd3_1
X_13061_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__buf_2
Xhold5671 _04305_ vssd1 vssd1 vccd1 vccd1 net6198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5682 net1524 vssd1 vssd1 vccd1 vccd1 net6209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5693 _04349_ vssd1 vssd1 vccd1 vccd1 net6220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12012_ net3569 net4960 _04845_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__mux2_1
Xhold4970 _01017_ vssd1 vssd1 vccd1 vccd1 net5497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4981 rbzero.floor_leak\[5\] vssd1 vssd1 vccd1 vccd1 net5508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4992 _00883_ vssd1 vssd1 vccd1 vccd1 net5519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ _09818_ _09209_ vssd1 vssd1 vccd1 vccd1 _09847_ sky130_fd_sc_hd__nand2_1
X_16751_ _09103_ _09784_ vssd1 vssd1 vccd1 vccd1 _09785_ sky130_fd_sc_hd__nand2_1
X_13963_ _06827_ _06863_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15702_ _08765_ _08796_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__xor2_1
X_19470_ net5998 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
X_12914_ net4576 net4550 net4293 _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__or4_1
X_16682_ net756 _09741_ _09742_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1
+ vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
X_13894_ _07063_ _07057_ _07061_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__nor3_1
XFILLER_0_186_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18421_ _02587_ _02602_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__xnor2_1
X_15633_ _08665_ _08673_ _08672_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _05997_ _06013_ _06016_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__or4b_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ net4733 _02528_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__nand2_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _08636_ _08637_ _08639_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__a21o_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _05950_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__nor2_4
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17303_ _08309_ _09170_ vssd1 vssd1 vccd1 vccd1 _10322_ sky130_fd_sc_hd__or2_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _04916_ vssd1 vssd1 vccd1 vccd1 _04917_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14515_ _07668_ _07684_ _07685_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__a21oi_1
X_15495_ _08589_ _08510_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18283_ net1539 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ _10017_ _10018_ _10127_ vssd1 vssd1 vccd1 vccd1 _10254_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ net7569 _04813_ _04834_ _04794_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__o211a_1
X_14446_ _07615_ _07616_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__or2b_1
Xclkbuf_1_1__f__03872_ clknet_0__03872_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03872_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _04104_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__clkbuf_4
X_17165_ _08338_ _08472_ _09135_ _08366_ vssd1 vssd1 vccd1 vccd1 _10185_ sky130_fd_sc_hd__a2bb2o_1
X_14377_ _07537_ _07546_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__or2_1
X_11589_ net1616 _04777_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__nand3_1
XFILLER_0_153_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold907 _00988_ vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold918 net6381 vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ _06456_ _06458_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__xnor2_1
X_16116_ net8216 net5904 _08111_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__mux2_1
X_17096_ _10114_ _10116_ vssd1 vssd1 vccd1 vccd1 _10117_ sky130_fd_sc_hd__nor2_1
Xhold929 net6406 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16047_ _08389_ _08308_ _08309_ _08211_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__o22ai_1
X_13259_ _06427_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3009 net8226 vssd1 vssd1 vccd1 vccd1 net3536 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2308 net5625 vssd1 vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2319 _04318_ vssd1 vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1607 net5652 vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 _01478_ vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _02158_ _02159_ _02233_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__and3_1
Xhold1629 _04142_ vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
X_19737_ net7655 net7648 _03496_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__and3_1
X_16949_ _08474_ _08494_ vssd1 vssd1 vccd1 vccd1 _09971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19668_ net6343 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18619_ net5927 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19599_ _03320_ net3843 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21630_ clknet_leaf_129_i_clk net3235 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_20474__218 clknet_1_0__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__inv_2
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21561_ net195 net2964 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21492_ clknet_leaf_5_i_clk net1407 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_i_clk clknet_4_14__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4200 net8077 vssd1 vssd1 vccd1 vccd1 net4727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22113_ clknet_leaf_62_i_clk net4970 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4211 _08057_ vssd1 vssd1 vccd1 vccd1 net4738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4222 _01192_ vssd1 vssd1 vccd1 vccd1 net4749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4233 net1681 vssd1 vssd1 vccd1 vccd1 net4760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4244 _02799_ vssd1 vssd1 vccd1 vccd1 net4771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3510 rbzero.spi_registers.spi_buffer\[4\] vssd1 vssd1 vccd1 vccd1 net4037 sky130_fd_sc_hd__dlygate4sd3_1
X_20368__123 clknet_1_1__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__inv_2
Xhold4255 _02319_ vssd1 vssd1 vccd1 vccd1 net4782 sky130_fd_sc_hd__clkbuf_2
X_22044_ net486 net2788 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
Xhold4266 _02624_ vssd1 vssd1 vccd1 vccd1 net4793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3521 net4006 vssd1 vssd1 vccd1 vccd1 net4048 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_66_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold4277 _01220_ vssd1 vssd1 vccd1 vccd1 net4804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3532 _09728_ vssd1 vssd1 vccd1 vccd1 net4059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4288 _02474_ vssd1 vssd1 vccd1 vccd1 net4815 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3543 net4137 vssd1 vssd1 vccd1 vccd1 net4070 sky130_fd_sc_hd__clkbuf_1
Xhold3554 _00482_ vssd1 vssd1 vccd1 vccd1 net4081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4299 _01231_ vssd1 vssd1 vccd1 vccd1 net4826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2820 _00719_ vssd1 vssd1 vccd1 vccd1 net3347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3565 _05675_ vssd1 vssd1 vccd1 vccd1 net4092 sky130_fd_sc_hd__clkbuf_4
Xhold2831 _01482_ vssd1 vssd1 vccd1 vccd1 net3358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3576 _05677_ vssd1 vssd1 vccd1 vccd1 net4103 sky130_fd_sc_hd__clkbuf_4
Xhold3587 _01246_ vssd1 vssd1 vccd1 vccd1 net4114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2842 _00930_ vssd1 vssd1 vccd1 vccd1 net3369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3598 _00472_ vssd1 vssd1 vccd1 vccd1 net4125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2853 net7994 vssd1 vssd1 vccd1 vccd1 net3380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2864 net8316 vssd1 vssd1 vccd1 vccd1 net3391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2875 net2003 vssd1 vssd1 vccd1 vccd1 net3402 sky130_fd_sc_hd__buf_2
XFILLER_0_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2886 _00708_ vssd1 vssd1 vccd1 vccd1 net3413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2897 net4911 vssd1 vssd1 vccd1 vccd1 net3424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ net7228 net3029 _04298_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10891_ _04103_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _05797_ net24 net25 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a21o_1
X_21828_ net270 net2708 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12561_ _05696_ _05740_ _05741_ net4141 vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__o22a_2
X_21759_ clknet_leaf_111_i_clk net4114 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14300_ _07469_ _07470_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__nand2_2
X_11512_ _04701_ _04460_ _04601_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or3b_1
X_15280_ net4397 _06120_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__nand2_1
X_12492_ net4138 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14231_ _07240_ _07198_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11443_ rbzero.spi_registers.texadd2\[3\] _04566_ _04567_ _04020_ vssd1 vssd1 vccd1
+ vccd1 _04635_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _07331_ _07332_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11374_ _04554_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6180 net1875 vssd1 vssd1 vccd1 vccd1 net6707 sky130_fd_sc_hd__dlygate4sd3_1
X_13113_ _06281_ _06282_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__and3_1
Xhold6191 rbzero.tex_g1\[37\] vssd1 vssd1 vccd1 vccd1 net6718 sky130_fd_sc_hd__dlygate4sd3_1
X_14093_ _07257_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__xnor2_1
X_18970_ net1559 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5490 net3735 vssd1 vssd1 vccd1 vccd1 net6017 sky130_fd_sc_hd__dlygate4sd3_1
X_17921_ _02141_ _02143_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__or2_1
X_13044_ _06211_ _06216_ _06218_ _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17852_ _02075_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16803_ _09831_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17783_ _08799_ _10220_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14995_ _08093_ net4141 vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19522_ net1427 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
X_16734_ net5554 _09103_ _09766_ vssd1 vssd1 vccd1 vccd1 _09771_ sky130_fd_sc_hd__a21bo_1
X_13946_ _07103_ _07116_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19453_ _03205_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__buf_4
XFILLER_0_202_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16665_ net4339 _09737_ _09740_ _07938_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ _07045_ _07046_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ net4698 net4733 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _08709_ _08710_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19384_ net6683 _03284_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or2_1
X_12828_ _05949_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or2b_1
X_16596_ _09551_ _09553_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18335_ net3565 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15547_ _08628_ _08641_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__xor2_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ net44 _05916_ _05915_ net46 vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__a22o_1
Xhold7809 rbzero.wall_tracer.stepDistX\[10\] vssd1 vssd1 vccd1 vccd1 net8336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ net1287 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__clkbuf_1
X_15478_ _08572_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17217_ _10235_ _10236_ vssd1 vssd1 vccd1 vccd1 _10237_ sky130_fd_sc_hd__nand2_2
X_14429_ _07584_ _07599_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__xor2_2
XFILLER_0_163_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03855_ clknet_0__03855_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03855_
+ sky130_fd_sc_hd__clkbuf_16
X_18197_ _09809_ _02416_ _02417_ _10380_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_170_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17148_ _09373_ _09600_ vssd1 vssd1 vccd1 vccd1 _10168_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 _03547_ vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 _02486_ vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 net5495 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 _03821_ vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold748 net5557 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _10098_ _10099_ vssd1 vssd1 vccd1 vccd1 _10100_ sky130_fd_sc_hd__xnor2_1
Xhold759 net6354 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20090_ _03682_ _03683_ _03610_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2105 net2214 vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2116 _01551_ vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2127 net7416 vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2138 net7076 vssd1 vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 _01060_ vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 net7183 vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 net4826 vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1426 net6769 vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1437 net7050 vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1448 _01347_ vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1459 net6785 vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20992_ clknet_leaf_111_i_clk net4119 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21613_ clknet_leaf_97_i_clk net1184 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21544_ net178 net1150 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21475_ clknet_leaf_21_i_clk net3845 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4030 net811 vssd1 vssd1 vccd1 vccd1 net4557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4041 net7957 vssd1 vssd1 vccd1 vccd1 net4568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4052 net3206 vssd1 vssd1 vccd1 vccd1 net4579 sky130_fd_sc_hd__dlygate4sd3_1
X_11090_ net2367 net7383 _04364_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
Xhold4063 rbzero.pov.ready_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net4590 sky130_fd_sc_hd__dlygate4sd3_1
X_20288_ net6374 net1492 _03814_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
Xhold4074 net8101 vssd1 vssd1 vccd1 vccd1 net4601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4085 net1154 vssd1 vssd1 vccd1 vccd1 net4612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3340 _03099_ vssd1 vssd1 vccd1 vccd1 net3867 sky130_fd_sc_hd__dlygate4sd3_1
X_22027_ net469 net1896 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
Xhold4096 net8338 vssd1 vssd1 vccd1 vccd1 net4623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3351 _03086_ vssd1 vssd1 vccd1 vccd1 net3878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3362 net8351 vssd1 vssd1 vccd1 vccd1 net3889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3373 _03079_ vssd1 vssd1 vccd1 vccd1 net3900 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3384 _02975_ vssd1 vssd1 vccd1 vccd1 net3911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2650 _04280_ vssd1 vssd1 vccd1 vccd1 net3177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3395 _03500_ vssd1 vssd1 vccd1 vccd1 net3922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2661 _01107_ vssd1 vssd1 vccd1 vccd1 net3188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold64 net5992 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2672 net3048 vssd1 vssd1 vccd1 vccd1 net3199 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2683 net3328 vssd1 vssd1 vccd1 vccd1 net3210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 _03603_ vssd1 vssd1 vccd1 vccd1 net3221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net4921 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 net4957 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _06715_ _06813_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__nand2_1
Xhold1960 _00672_ vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net6027 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1971 _01584_ vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _04467_ _05178_ _05180_ _04659_ net7716 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__o32a_1
X_14780_ _07926_ _07944_ _07913_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__mux2_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1982 net7038 vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1993 _01456_ vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
X_10943_ net7316 net2482 _04287_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__mux2_1
X_13731_ _06900_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__xnor2_1
X_20422__172 clknet_1_1__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__inv_2
X_16450_ net4520 _06123_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__nand2_2
XFILLER_0_211_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10874_ net6595 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__clkbuf_1
X_13662_ _06693_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _08492_ _08493_ _08495_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__a21oi_4
X_12613_ _05747_ net18 _05748_ _05754_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a41o_2
X_16381_ _09471_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__buf_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _06576_ _06754_ _06702_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ net3732 _02343_ _02344_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a21boi_1
X_15332_ _08421_ _08424_ _08426_ _08133_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__a211o_2
X_12544_ net44 _05700_ _05698_ net4147 vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a22o_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18051_ _02285_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15263_ _08207_ _08266_ _08357_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12475_ _05655_ _05656_ net7 vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17002_ _10021_ _10022_ vssd1 vssd1 vccd1 vccd1 _10023_ sky130_fd_sc_hd__nor2_2
X_14214_ _07372_ _07384_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__xnor2_1
X_11426_ _04521_ _04531_ _04533_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15194_ _08288_ net3445 _06027_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__mux2_2
XANTENNA_6 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14145_ _07314_ _07315_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__xor2_1
X_11357_ rbzero.spi_registers.texadd1\[14\] vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14076_ _07221_ _07222_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__or2_1
X_18953_ net3253 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
X_11288_ net3871 net3976 _04476_ _04482_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o31ai_2
X_17904_ _02040_ _02041_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__nor2_1
X_13027_ _06201_ net3790 _06202_ net4567 vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__o22a_1
X_18884_ net6233 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
X_17835_ _01807_ _02003_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17766_ _02001_ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__xnor2_1
Xrebuffer18 net557 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ net4624 _08021_ _08079_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__mux2_1
Xrebuffer29 net555 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19505_ net1426 net5500 _03365_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16717_ _06104_ net7713 vssd1 vssd1 vccd1 vccd1 _09755_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13929_ _06854_ _06860_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__a21bo_1
X_17697_ _01935_ _01936_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19436_ _03320_ net3548 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ net4133 _04664_ net5948 vssd1 vssd1 vccd1 vccd1 _09729_ sky130_fd_sc_hd__and3_1
X_19782__61 clknet_1_1__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
XFILLER_0_18_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19367_ net1785 _03284_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__or2_1
X_16579_ _09540_ _09541_ _08401_ vssd1 vssd1 vccd1 vccd1 _09669_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ net6333 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7606 _00504_ vssd1 vssd1 vccd1 vccd1 net8133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7617 rbzero.spi_registers.vshift\[3\] vssd1 vssd1 vccd1 vccd1 net8144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19298_ _03205_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__buf_4
Xhold7628 rbzero.spi_registers.vshift\[1\] vssd1 vssd1 vccd1 vccd1 net8155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7639 rbzero.map_overlay.i_mapdx\[0\] vssd1 vssd1 vccd1 vccd1 net8166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6905 rbzero.tex_g0\[29\] vssd1 vssd1 vccd1 vccd1 net7432 sky130_fd_sc_hd__dlygate4sd3_1
X_18249_ _02463_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6916 net3022 vssd1 vssd1 vccd1 vccd1 net7443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6927 rbzero.pov.spi_buffer\[59\] vssd1 vssd1 vccd1 vccd1 net7454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6938 net663 vssd1 vssd1 vccd1 vccd1 net7465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6949 rbzero.tex_g0\[48\] vssd1 vssd1 vccd1 vccd1 net7476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21260_ clknet_leaf_22_i_clk net3942 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold501 net8066 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20586__319 clknet_1_0__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__inv_2
XFILLER_0_29_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold512 net8011 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 net5439 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
X_20211_ net4423 _03744_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__or2_1
Xhold534 net6493 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 net6171 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03869_ _03869_ vssd1 vssd1 vccd1 vccd1 clknet_0__03869_ sky130_fd_sc_hd__clkbuf_16
X_21191_ clknet_leaf_129_i_clk net3278 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold556 net6167 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold567 _01646_ vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 net7909 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_1
X_20142_ net7334 _03707_ net4595 _03679_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__o211a_1
Xhold589 _04090_ vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20073_ net3414 _03485_ _03662_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a211o_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _03110_ vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 net6590 vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 _01472_ vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1234 net6745 vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1245 _00980_ vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 net6724 vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1267 net6358 vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1278 net6592 vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 _01086_ vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20975_ clknet_leaf_110_i_clk net4175 vssd1 vssd1 vccd1 vccd1 reg_rgb\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10590_ net2948 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21527_ clknet_leaf_119_i_clk net4999 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ _05206_ _05446_ _04829_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__o21a_1
X_21458_ clknet_leaf_42_i_clk net1431 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20452__198 clknet_1_1__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__inv_2
X_11211_ net6850 net2854 _04423_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12191_ net3976 _04653_ net4148 _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21389_ clknet_leaf_20_i_clk net5250 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11142_ net6804 net2512 _04390_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__clkbuf_4
X_11073_ net1797 net6128 _04353_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15950_ _08420_ _08469_ _09044_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__a21bo_1
Xhold3170 _02990_ vssd1 vssd1 vccd1 vccd1 net3697 sky130_fd_sc_hd__dlygate4sd3_1
X_14901_ net4268 _08037_ _08043_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__o21a_1
Xhold3181 _03497_ vssd1 vssd1 vccd1 vccd1 net3708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3192 rbzero.debug_overlay.facingX\[-1\] vssd1 vssd1 vccd1 vccd1 net3719 sky130_fd_sc_hd__buf_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _08928_ _08975_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__nor2_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2480 _01028_ vssd1 vssd1 vccd1 vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _10190_ _09225_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2491 rbzero.pov.spi_buffer\[8\] vssd1 vssd1 vccd1 vccd1 net3018 sky130_fd_sc_hd__dlygate4sd3_1
X_14832_ net8362 _07988_ _07990_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_204_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03858_ clknet_0__03858_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03858_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1790 _01027_ vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
X_17551_ _10327_ _10096_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__nor2_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14763_ net4403 _07929_ _07872_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ net4598 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16502_ _09467_ _09496_ _09591_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__a21boi_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ _06785_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17482_ _10269_ _10270_ _10374_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a21o_1
X_10926_ net6072 net3107 _04276_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14694_ _07860_ _07861_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__a21o_1
XFILLER_0_211_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19221_ net1030 _03140_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__and2_1
X_16433_ _09402_ _09406_ _09405_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__a21oi_1
X_10857_ net6295 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__clkbuf_1
X_13645_ _06719_ net572 vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__nor2_2
XFILLER_0_186_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ _09721_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__clkbuf_4
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__xnor2_1
X_10788_ net2460 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__clkbuf_1
X_13576_ _06742_ _06743_ _06746_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a21o_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _02328_ _02329_ net3730 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__o21a_1
X_15315_ net3600 _06121_ _08408_ _08409_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19083_ net2056 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__clkbuf_1
X_12527_ net13 net12 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__and2b_1
X_16295_ _09385_ _09386_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18034_ _02268_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__xor2_1
X_15246_ net3822 _08128_ _08139_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12458_ net9 net8 vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11409_ _04462_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nor2_2
X_15177_ _08271_ _08241_ _08252_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__or3b_2
X_12389_ _04949_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14128_ _07272_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__xnor2_1
X_19985_ net7272 net7502 _08092_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14059_ _07228_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__and2_4
X_18936_ net1103 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20429__178 clknet_1_1__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__inv_2
XFILLER_0_158_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18867_ net1971 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17818_ net4655 net4756 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ _02943_ _02929_ _04480_ _02866_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a211o_1
X_17749_ _01896_ _01900_ _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20760_ _03930_ _03931_ _03932_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19419_ net4964 _03310_ _03315_ _03316_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__a211o_1
X_20691_ net777 net4968 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7403 rbzero.wall_tracer.trackDistX\[-10\] vssd1 vssd1 vccd1 vccd1 net7930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7414 net4391 vssd1 vssd1 vccd1 vccd1 net7941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7425 net4564 vssd1 vssd1 vccd1 vccd1 net7952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7436 rbzero.wall_tracer.trackDistX\[3\] vssd1 vssd1 vccd1 vccd1 net7963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6702 _04301_ vssd1 vssd1 vccd1 vccd1 net7229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7447 net4654 vssd1 vssd1 vccd1 vccd1 net7974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6713 net2253 vssd1 vssd1 vccd1 vccd1 net7240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7458 rbzero.wall_tracer.trackDistX\[-2\] vssd1 vssd1 vccd1 vccd1 net7985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6724 rbzero.tex_r0\[5\] vssd1 vssd1 vccd1 vccd1 net7251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7469 net4580 vssd1 vssd1 vccd1 vccd1 net7996 sky130_fd_sc_hd__dlygate4sd3_1
X_21312_ clknet_leaf_7_i_clk net5067 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6735 net2820 vssd1 vssd1 vccd1 vccd1 net7262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6746 _03486_ vssd1 vssd1 vccd1 vccd1 net7273 sky130_fd_sc_hd__buf_2
Xhold6757 rbzero.tex_r0\[8\] vssd1 vssd1 vccd1 vccd1 net7284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6768 net2774 vssd1 vssd1 vccd1 vccd1 net7295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6779 net2694 vssd1 vssd1 vccd1 vccd1 net7306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold320 net5357 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
X_21243_ clknet_leaf_16_i_clk net3404 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 net5215 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold342 net5333 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 net5196 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 net4348 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
X_21174_ clknet_leaf_97_i_clk net2081 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold375 net5295 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold386 net5335 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 net6106 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
X_20125_ net3407 _03707_ net4626 _03679_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20056_ net41 _03605_ _03123_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__o21a_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 net7696 vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__buf_2
Xhold1031 net3120 vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 _01154_ vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 net6662 vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20640__368 clknet_1_0__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__inv_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 net6081 vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 net6527 vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 net6664 vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _00936_ vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _04836_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__buf_4
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20958_ clknet_leaf_66_i_clk _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ net7037 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__clkbuf_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _04467_ _04865_ _04860_ _04022_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__o221a_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ net6041 net4948 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__xnor2_1
X_19761__42 clknet_1_1__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_0_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10642_ net6824 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13430_ _06548_ _06464_ _06525_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ _06519_ _06521_ _06502_ _06524_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__and4bb_2
X_10573_ net6900 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20534__273 clknet_1_1__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__inv_2
XFILLER_0_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ net5887 _08194_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__nand2_1
X_12312_ _04825_ _05485_ _05489_ _05497_ _04844_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__o311a_1
Xrebuffer9 _07026_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_1
X_13292_ _06435_ _06442_ _06462_ _06450_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__or4_4
Xhold7970 _05999_ vssd1 vssd1 vccd1 vccd1 net8497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16080_ _08114_ _09172_ _09173_ _08441_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7992 rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 net8519 sky130_fd_sc_hd__dlygate4sd3_1
X_12243_ _04977_ _05427_ _05429_ _04988_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15031_ _08119_ _08121_ _08125_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12174_ _04910_ _05361_ _04828_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ net6267 net2351 _04030_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16982_ _09707_ _10003_ vssd1 vssd1 vccd1 vccd1 _10004_ sky130_fd_sc_hd__nand2_2
X_18721_ _02849_ _02853_ _02871_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a21o_1
X_11056_ net5634 net6766 _04342_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
X_15933_ _09026_ _09027_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18652_ _02559_ net8027 net4772 net3534 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__a31o_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _08126_ _08474_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__nor2_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _01841_ _01842_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a21o_2
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ net3775 vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__buf_4
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ net7706 net4049 net4648 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
X_15795_ _08885_ _08888_ _08889_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__a21oi_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_100 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_100/HI o_rgb[9] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_111 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_111/HI zeros[0] sky130_fd_sc_hd__conb_1
XFILLER_0_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_122 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_122/HI zeros[11]
+ sky130_fd_sc_hd__conb_1
X_17534_ _01773_ _01774_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__nor2_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_133 vssd1 vssd1 vccd1 vccd1 ones[6] top_ew_algofoogle_133/LO sky130_fd_sc_hd__conb_1
XFILLER_0_169_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _07821_ _07861_ _07888_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_197_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11958_ rbzero.debug_overlay.facingY\[-2\] _05080_ _05103_ rbzero.debug_overlay.facingY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10909_ net7397 net6762 _04265_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__mux2_1
X_17465_ _10336_ _10359_ _10357_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14677_ _07844_ _07847_ net8354 vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11889_ _05070_ _05077_ net3517 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_200_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19204_ net5232 _03182_ _03190_ _03189_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16416_ _09505_ _09506_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13628_ _06797_ _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17396_ _10412_ _10413_ vssd1 vssd1 vccd1 vccd1 _10414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19135_ net1203 _03147_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or2_1
X_16347_ _09436_ _09438_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ _06729_ _06727_ _06725_ _06726_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__nand4_1
Xhold6009 net1500 vssd1 vssd1 vccd1 vccd1 net6536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19066_ net3794 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16278_ _09340_ _09369_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5308 net3411 vssd1 vssd1 vccd1 vccd1 net5835 sky130_fd_sc_hd__buf_1
XFILLER_0_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20665__11 clknet_1_0__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
Xhold5319 _00640_ vssd1 vssd1 vccd1 vccd1 net5846 sky130_fd_sc_hd__dlygate4sd3_1
X_18017_ _02148_ _02252_ _02235_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a21oi_1
X_15229_ _08318_ _08323_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__or2_2
XFILLER_0_164_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4607 _00849_ vssd1 vssd1 vccd1 vccd1 net5134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4618 net771 vssd1 vssd1 vccd1 vccd1 net5145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4629 rbzero.mapdxw\[0\] vssd1 vssd1 vccd1 vccd1 net5156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3906 net1240 vssd1 vssd1 vccd1 vccd1 net4433 sky130_fd_sc_hd__dlygate4sd3_1
X_20680__25 clknet_1_0__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3917 _01172_ vssd1 vssd1 vccd1 vccd1 net4444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3928 _03645_ vssd1 vssd1 vccd1 vccd1 net4455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19968_ net2313 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
X_18919_ net3302 net7565 _03025_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19899_ net2935 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
X_21930_ net372 net3154 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21861_ net303 net2356 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20812_ net8222 _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__xnor2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21792_ net234 net2353 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20743_ _03914_ _03915_ _03916_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_175_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7200 net4173 vssd1 vssd1 vccd1 vccd1 net7727 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7211 gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 net7738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7222 rbzero.trace_state\[1\] vssd1 vssd1 vccd1 vccd1 net7749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7244 net3461 vssd1 vssd1 vccd1 vccd1 net7771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6510 net2762 vssd1 vssd1 vccd1 vccd1 net7037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6521 rbzero.tex_g1\[6\] vssd1 vssd1 vccd1 vccd1 net7048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7266 _06544_ vssd1 vssd1 vccd1 vccd1 net7793 sky130_fd_sc_hd__buf_1
XFILLER_0_104_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6532 net2211 vssd1 vssd1 vccd1 vccd1 net7059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6543 rbzero.tex_g0\[25\] vssd1 vssd1 vccd1 vccd1 net7070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7288 net4755 vssd1 vssd1 vccd1 vccd1 net7815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6554 net2751 vssd1 vssd1 vccd1 vccd1 net7081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7299 rbzero.wall_tracer.stepDistY\[2\] vssd1 vssd1 vccd1 vccd1 net7826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5820 net1325 vssd1 vssd1 vccd1 vccd1 net6347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6565 rbzero.pov.ready_buffer\[42\] vssd1 vssd1 vccd1 vccd1 net7092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6576 net1842 vssd1 vssd1 vccd1 vccd1 net7103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5831 rbzero.tex_r0\[0\] vssd1 vssd1 vccd1 vccd1 net6358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6587 _04454_ vssd1 vssd1 vccd1 vccd1 net7114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5842 rbzero.spi_registers.new_texadd\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net6369
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5853 net1444 vssd1 vssd1 vccd1 vccd1 net6380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6598 net2679 vssd1 vssd1 vccd1 vccd1 net7125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 net4711 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ clknet_leaf_121_i_clk net1711 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5864 _02488_ vssd1 vssd1 vccd1 vccd1 net6391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5875 _03452_ vssd1 vssd1 vccd1 vccd1 net6402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5886 net1316 vssd1 vssd1 vccd1 vccd1 net6413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 net5014 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5897 net1497 vssd1 vssd1 vccd1 vccd1 net6424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 net5028 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 net5042 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 net5128 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
X_21157_ clknet_leaf_2_i_clk net5866 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20108_ net3552 _03694_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21088_ clknet_leaf_13_i_clk net1283 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20564__299 clknet_1_0__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__inv_2
XFILLER_0_176_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20039_ net3389 _03607_ net4455 _03628_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__o211a_1
X_12930_ net4354 _06104_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__nand2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ net4641 vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__inv_2
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _07768_ _07769_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__or3_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04938_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__or2_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15580_ _08665_ _08674_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _05964_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__or2_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _07699_ _07700_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _04836_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__buf_4
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _10246_ _10248_ vssd1 vssd1 vccd1 vccd1 _10269_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14462_ _07632_ _07613_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ net3014 _04858_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16201_ _08024_ net75 vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__or2_1
X_13413_ _06522_ _06531_ _06533_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__and3_1
X_10625_ net7371 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17181_ _10068_ _10069_ _10200_ vssd1 vssd1 vccd1 vccd1 _10201_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14393_ _07561_ _07563_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16132_ _09224_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__clkbuf_4
X_10556_ net2880 net7226 _04086_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__mux2_1
X_13344_ net574 _06514_ _06485_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16063_ _08244_ _08414_ _08386_ _08246_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__a22o_1
X_10487_ net2985 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__clkbuf_1
X_13275_ _06404_ _06353_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__and2_2
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ net4013 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__clkbuf_1
X_12226_ _04921_ _05410_ _05412_ _04829_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__o211a_1
X_12157_ _04910_ _05344_ _04828_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__o21a_1
X_19822_ net3211 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11108_ net2602 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16965_ _09984_ _09985_ _09963_ vssd1 vssd1 vccd1 vccd1 _09987_ sky130_fd_sc_hd__a21oi_1
X_12088_ rbzero.tex_r1\[63\] rbzero.tex_r1\[62\] _04913_ vssd1 vssd1 vccd1 vccd1 _05277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11039_ _04193_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__clkbuf_4
X_15916_ _09001_ _09010_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__xnor2_1
X_18704_ _02856_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02857_
+ sky130_fd_sc_hd__nand2_1
X_19684_ net6417 net3838 _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__mux2_1
X_16896_ _09914_ _09917_ vssd1 vssd1 vccd1 vccd1 _09918_ sky130_fd_sc_hd__and2b_1
XFILLER_0_190_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18635_ net3678 rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _02793_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _08529_ _08494_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__nor2_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ net3962 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
X_15778_ _08869_ _08872_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__xor2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17517_ _01756_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__xor2_1
XFILLER_0_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14729_ _07843_ _07895_ _07897_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__a21oi_1
X_18497_ _02626_ net4554 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ _01688_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _08167_ net4914 _10278_ vssd1 vssd1 vccd1 vccd1 _10397_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19118_ net1803 _03125_ net5536 _03128_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5105 net1749 vssd1 vssd1 vccd1 vccd1 net5632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5116 _01343_ vssd1 vssd1 vccd1 vccd1 net5643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5127 _04322_ vssd1 vssd1 vccd1 vccd1 net5654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19049_ net3593 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5138 rbzero.wall_tracer.mapX\[7\] vssd1 vssd1 vccd1 vccd1 net5665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5149 rbzero.tex_r1\[38\] vssd1 vssd1 vccd1 vccd1 net5676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4404 gpout0.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4415 net605 vssd1 vssd1 vccd1 vccd1 net4942 sky130_fd_sc_hd__dlygate4sd3_1
X_22060_ net502 net2769 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold4426 _00894_ vssd1 vssd1 vccd1 vccd1 net4953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4437 net621 vssd1 vssd1 vccd1 vccd1 net4964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3703 net8144 vssd1 vssd1 vccd1 vccd1 net4230 sky130_fd_sc_hd__buf_1
Xhold4448 rbzero.spi_registers.texadd3\[23\] vssd1 vssd1 vccd1 vccd1 net4975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3714 net835 vssd1 vssd1 vccd1 vccd1 net4241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4459 net659 vssd1 vssd1 vccd1 vccd1 net4986 sky130_fd_sc_hd__dlygate4sd3_1
X_21011_ clknet_leaf_38_i_clk net1823 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3725 net851 vssd1 vssd1 vccd1 vccd1 net4252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3736 net8010 vssd1 vssd1 vccd1 vccd1 net4263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3747 rbzero.wall_tracer.visualWallDist\[0\] vssd1 vssd1 vccd1 vccd1 net4274 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3758 _01190_ vssd1 vssd1 vccd1 vccd1 net4285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21913_ net355 net2422 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21844_ net286 net2210 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21775_ clknet_leaf_46_i_clk net1216 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20726_ net1120 net5252 vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7030 rbzero.spi_registers.new_other\[8\] vssd1 vssd1 vccd1 vccd1 net7557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7041 rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 net7568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7052 net3478 vssd1 vssd1 vccd1 vccd1 net7579 sky130_fd_sc_hd__dlygate4sd3_1
X_11390_ _04578_ _04545_ _04581_ _04503_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__o211a_1
Xhold7063 _03097_ vssd1 vssd1 vccd1 vccd1 net7590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7074 net3583 vssd1 vssd1 vccd1 vccd1 net7601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6340 rbzero.tex_b0\[13\] vssd1 vssd1 vccd1 vccd1 net6867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7085 rbzero.pov.ready_buffer\[32\] vssd1 vssd1 vccd1 vccd1 net7612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6351 net1932 vssd1 vssd1 vccd1 vccd1 net6878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7096 _03737_ vssd1 vssd1 vccd1 vccd1 net7623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6362 rbzero.tex_b1\[7\] vssd1 vssd1 vccd1 vccd1 net6889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6373 net2337 vssd1 vssd1 vccd1 vccd1 net6900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6384 _04184_ vssd1 vssd1 vccd1 vccd1 net6911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6395 net2271 vssd1 vssd1 vccd1 vccd1 net6922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5650 _03839_ vssd1 vssd1 vccd1 vccd1 net6177 sky130_fd_sc_hd__dlygate4sd3_1
X_13060_ net4646 net4780 vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and2_1
Xhold5661 _04117_ vssd1 vssd1 vccd1 vccd1 net6188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5672 net1131 vssd1 vssd1 vccd1 vccd1 net6199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5683 rbzero.tex_g1\[14\] vssd1 vssd1 vccd1 vccd1 net6210 sky130_fd_sc_hd__dlygate4sd3_1
X_12011_ _05176_ _05199_ _04751_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__o21ba_1
Xhold5694 net1186 vssd1 vssd1 vccd1 vccd1 net6221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21209_ clknet_leaf_117_i_clk net1790 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4960 rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 net5487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4971 net1254 vssd1 vssd1 vccd1 vccd1 net5498 sky130_fd_sc_hd__dlygate4sd3_1
X_20646__374 clknet_1_1__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__inv_2
Xhold4982 net1414 vssd1 vssd1 vccd1 vccd1 net5509 sky130_fd_sc_hd__buf_1
XFILLER_0_100_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4993 net1551 vssd1 vssd1 vccd1 vccd1 net5520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20345__102 clknet_1_0__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__inv_2
X_16750_ net5328 _09783_ vssd1 vssd1 vccd1 vccd1 _09784_ sky130_fd_sc_hd__xnor2_1
X_13962_ _06864_ _06752_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__or2b_1
X_15701_ _08739_ _08766_ _08781_ _08793_ _08795_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__a32o_1
X_12913_ net4737 net4690 net4694 net4584 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__or4_1
X_16681_ net777 _09741_ _09742_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1
+ vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
X_13893_ _07057_ _07061_ _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o21a_1
X_18420_ _02600_ _02601_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__nand2_1
X_15632_ _08676_ _08677_ _08687_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__a21o_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__or2_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18351_ net5963 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__clkbuf_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15563_ _08642_ _08643_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__xnor2_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _10319_ _10320_ vssd1 vssd1 vccd1 vccd1 _10321_ sky130_fd_sc_hd__and2_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _07669_ _07670_ _07683_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__and3_1
X_11726_ _04835_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__clkbuf_8
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ net6492 net3863 _02477_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
X_15494_ _08511_ _08508_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _10250_ _10252_ vssd1 vssd1 vccd1 vccd1 _10253_ sky130_fd_sc_hd__xor2_4
XFILLER_0_65_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14445_ _07572_ _07574_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1__f__03871_ clknet_0__03871_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03871_
+ sky130_fd_sc_hd__clkbuf_16
X_11657_ net88 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__buf_4
X_20391__144 clknet_1_0__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__inv_2
X_10608_ net2385 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__clkbuf_1
X_17164_ _10083_ _10092_ _10091_ vssd1 vssd1 vccd1 vccd1 _10184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14376_ _07537_ _07546_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__xor2_4
X_11588_ net1075 net1658 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16115_ _09108_ _09208_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__xor2_4
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13327_ _06345_ _06497_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__xnor2_4
Xhold908 net6306 vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17095_ _09953_ _09990_ _10115_ vssd1 vssd1 vccd1 vccd1 _10116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10539_ net6752 net6754 _04075_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold919 _00587_ vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16046_ _08389_ _08211_ _08294_ _08306_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ _06410_ _06418_ _06428_ _06385_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ _04847_ _05395_ net86 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _06296_ _06299_ _06297_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a21o_1
Xhold2309 net5627 vssd1 vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1608 net5654 vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ _02158_ _02159_ _02233_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1619 net6738 vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19789__67 clknet_1_1__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
X_16948_ _08181_ _09673_ _09969_ vssd1 vssd1 vccd1 vccd1 _09970_ sky130_fd_sc_hd__a21oi_4
X_19736_ net3923 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ _09899_ _09900_ vssd1 vssd1 vccd1 vccd1 _09901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667_ net6341 net1492 _03457_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18618_ net5925 _02777_ _02664_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
X_19598_ net3770 _02472_ net1777 _03139_ net3842 vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18549_ _06034_ _06036_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21560_ net194 net2609 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21491_ clknet_leaf_8_i_clk net1485 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4201 net3640 vssd1 vssd1 vccd1 vccd1 net4728 sky130_fd_sc_hd__dlygate4sd3_1
X_22112_ clknet_leaf_87_i_clk net921 vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4212 _00427_ vssd1 vssd1 vccd1 vccd1 net4739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4223 net618 vssd1 vssd1 vccd1 vccd1 net4750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4234 net8273 vssd1 vssd1 vccd1 vccd1 net4761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4245 _02804_ vssd1 vssd1 vccd1 vccd1 net4772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3500 rbzero.spi_registers.spi_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net4027 sky130_fd_sc_hd__dlygate4sd3_1
X_22043_ net485 net2916 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
Xhold3511 net4015 vssd1 vssd1 vccd1 vccd1 net4038 sky130_fd_sc_hd__buf_1
Xhold4267 net8110 vssd1 vssd1 vccd1 vccd1 net4794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3522 _06060_ vssd1 vssd1 vccd1 vccd1 net4049 sky130_fd_sc_hd__buf_2
Xhold3533 _00476_ vssd1 vssd1 vccd1 vccd1 net4060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4278 net675 vssd1 vssd1 vccd1 vccd1 net4805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4289 _03427_ vssd1 vssd1 vccd1 vccd1 net4816 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3544 _05674_ vssd1 vssd1 vccd1 vccd1 net4071 sky130_fd_sc_hd__clkbuf_4
Xhold2810 net4187 vssd1 vssd1 vccd1 vccd1 net3337 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3555 net7749 vssd1 vssd1 vccd1 vccd1 net4082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2821 net7764 vssd1 vssd1 vccd1 vccd1 net3348 sky130_fd_sc_hd__clkbuf_2
Xhold3566 net7717 vssd1 vssd1 vccd1 vccd1 net4093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2832 net7968 vssd1 vssd1 vccd1 vccd1 net3359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3577 _01244_ vssd1 vssd1 vccd1 vccd1 net4104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2843 net5886 vssd1 vssd1 vccd1 vccd1 net3370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3588 net7709 vssd1 vssd1 vccd1 vccd1 net4115 sky130_fd_sc_hd__clkbuf_2
Xhold3599 net7618 vssd1 vssd1 vccd1 vccd1 net4126 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2854 net4676 vssd1 vssd1 vccd1 vccd1 net3381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2865 net7986 vssd1 vssd1 vccd1 vccd1 net3392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2876 _03088_ vssd1 vssd1 vccd1 vccd1 net3403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2887 net7572 vssd1 vssd1 vccd1 vccd1 net3414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2898 net4692 vssd1 vssd1 vccd1 vccd1 net3425 sky130_fd_sc_hd__dlygate4sd3_1
X_10890_ net7053 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21827_ net269 net2359 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12560_ _05701_ _05718_ _05713_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nand3_1
XFILLER_0_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21758_ clknet_leaf_111_i_clk net4026 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11511_ _04022_ _04467_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__or2_1
X_20709_ net754 net5400 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ net4095 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21689_ clknet_leaf_28_i_clk net5871 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _07399_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__nand2_2
X_11442_ rbzero.spi_registers.texadd1\[2\] _04548_ vssd1 vssd1 vccd1 vccd1 _04634_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_184_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14161_ _07239_ _07322_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__xor2_1
X_11373_ _04561_ _04562_ _04563_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6170 net1770 vssd1 vssd1 vccd1 vccd1 net6697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6181 _03013_ vssd1 vssd1 vccd1 vccd1 net6708 sky130_fd_sc_hd__dlygate4sd3_1
X_13112_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6192 net2429 vssd1 vssd1 vccd1 vccd1 net6719 sky130_fd_sc_hd__dlygate4sd3_1
X_14092_ _07258_ _07261_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__and3_1
Xhold5480 net2060 vssd1 vssd1 vccd1 vccd1 net6007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5491 rbzero.spi_registers.new_floor\[0\] vssd1 vssd1 vccd1 vccd1 net6018 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _02157_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__clkbuf_1
X_13043_ _06217_ net3766 _06209_ net4589 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o2bb2a_1
X_17851_ _02080_ _02088_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__xnor2_1
Xhold4790 _00844_ vssd1 vssd1 vccd1 vccd1 net5317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16802_ _09830_ net4541 net4649 vssd1 vssd1 vccd1 vccd1 _09831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17782_ _02019_ _02020_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__and2_1
X_14994_ net4150 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16733_ net5666 _09102_ vssd1 vssd1 vccd1 vccd1 _09770_ sky130_fd_sc_hd__xor2_1
X_19521_ net1426 net6486 net3086 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux2_1
X_13945_ _07114_ _07115_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19452_ net5562 _03335_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__or2_1
X_16664_ net4343 _09737_ _09740_ _07929_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
X_13876_ _07043_ _07044_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15615_ net8414 _08225_ _08227_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__or3_1
X_18403_ net8075 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__inv_2
X_19383_ net5189 _03283_ _03294_ _03288_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__o211a_1
X_12827_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16595_ _09682_ _09683_ _09671_ vssd1 vssd1 vccd1 vccd1 _09685_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _02519_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__xor2_1
X_15546_ _08636_ _08640_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__and2_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ net43 _05902_ net36 net37 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a211o_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11709_ net4132 _04889_ _04896_ net4115 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a22o_1
X_18265_ net6355 net1622 _02477_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
X_15477_ _06119_ net8033 vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__nor2_1
X_12689_ net55 _05864_ _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17216_ _10207_ _10234_ vssd1 vssd1 vccd1 vccd1 _10236_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ _07585_ _07597_ _07598_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_1_1__f__03854_ clknet_0__03854_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03854_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18196_ _02414_ _02415_ _02407_ _02411_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _10042_ _10165_ _10166_ vssd1 vssd1 vccd1 vccd1 _10167_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold705 _01113_ vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ _07461_ _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__nand2_1
Xhold716 _00576_ vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_14__f_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold727 net5497 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 _01260_ vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17078_ _09974_ _09975_ _08948_ vssd1 vssd1 vccd1 vccd1 _10099_ sky130_fd_sc_hd__a21oi_1
Xhold749 net5559 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
X_16029_ _09059_ _09065_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2106 _04355_ vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2117 net3877 vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2128 _04411_ vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2139 _01288_ vssd1 vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1405 net6877 vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 net6968 vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1427 _01038_ vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 net7052 vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1449 net6835 vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
X_19719_ net5280 net7273 _03488_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20991_ clknet_leaf_110_i_clk net3518 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_133_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21612_ clknet_leaf_133_i_clk net2773 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21543_ net177 net2074 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21474_ clknet_leaf_18_i_clk net888 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_mapd
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4020 net3854 vssd1 vssd1 vccd1 vccd1 net4547 sky130_fd_sc_hd__clkbuf_2
Xhold4031 net8340 vssd1 vssd1 vccd1 vccd1 net4558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4042 net3801 vssd1 vssd1 vccd1 vccd1 net4569 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4053 net7995 vssd1 vssd1 vccd1 vccd1 net4580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20287_ net1556 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
Xhold4064 net1171 vssd1 vssd1 vccd1 vccd1 net4591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4075 net682 vssd1 vssd1 vccd1 vccd1 net4602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3330 net7707 vssd1 vssd1 vccd1 vccd1 net3857 sky130_fd_sc_hd__clkbuf_2
X_22026_ net468 net1074 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3341 _00740_ vssd1 vssd1 vccd1 vccd1 net3868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4086 _09216_ vssd1 vssd1 vccd1 vccd1 net4613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3352 _00728_ vssd1 vssd1 vccd1 vccd1 net3879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4097 net3832 vssd1 vssd1 vccd1 vccd1 net4624 sky130_fd_sc_hd__clkbuf_2
Xhold3374 _00721_ vssd1 vssd1 vccd1 vccd1 net3901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2640 _03564_ vssd1 vssd1 vccd1 vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3385 _00641_ vssd1 vssd1 vccd1 vccd1 net3912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2651 _01376_ vssd1 vssd1 vccd1 vccd1 net3178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3396 net7650 vssd1 vssd1 vccd1 vccd1 net3923 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2662 net5738 vssd1 vssd1 vccd1 vccd1 net3189 sky130_fd_sc_hd__buf_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold65 _01473_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2673 _03600_ vssd1 vssd1 vccd1 vccd1 net3200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2684 _03519_ vssd1 vssd1 vccd1 vccd1 net3211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net4923 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
X_19768__48 clknet_1_1__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1950 _04248_ vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net4943 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2695 _01165_ vssd1 vssd1 vccd1 vccd1 net3222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1961 net7376 vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold98 _01081_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1972 net7164 vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net4160 _04462_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__o21ai_1
Xhold1983 net7040 vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1994 net7335 vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
X_13730_ _06788_ _06789_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__xnor2_1
X_10942_ net7073 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13661_ _06769_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__buf_4
XFILLER_0_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20457__203 clknet_1_0__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__inv_2
X_10873_ net6593 net2886 _04253_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15400_ _08494_ _08472_ _08366_ _08464_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_183_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12612_ _05774_ _05782_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nand3_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _06124_ _09413_ net7837 vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__or3b_2
XFILLER_0_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _06692_ _06755_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__nor2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _04511_ _05989_ _08114_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__o211a_2
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ net4066 _05701_ _05699_ net71 vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a22o_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ _01760_ net4908 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15262_ _08355_ _08356_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12474_ _04020_ _04495_ _04494_ _04500_ _05633_ net5 vssd1 vssd1 vccd1 vccd1 _05656_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17001_ _09927_ _10019_ _10020_ vssd1 vssd1 vccd1 vccd1 _10022_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14213_ _07378_ _07377_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _04614_ _04616_ _04503_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__mux2_1
X_15193_ net3445 _08256_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _05743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14144_ _07242_ _07281_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11356_ _04505_ _04504_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__and2b_2
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14075_ _07203_ _07220_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__nand2_1
X_18952_ net7453 net7471 _03036_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
X_11287_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13026_ net4665 vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__inv_2
X_17903_ _02064_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18883_ net6231 net638 _03003_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
X_17834_ _02021_ _02029_ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14977_ _08086_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
X_17765_ _01807_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer19 _06663_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_1
X_19504_ net2257 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ _06852_ _06861_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _06068_ _08194_ vssd1 vssd1 vccd1 vccd1 _09754_ sky130_fd_sc_hd__xnor2_1
X_17696_ _01780_ _01830_ _01828_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19435_ net1564 net3547 _03323_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16647_ net4118 net4124 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13859_ _07027_ net529 vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16578_ _09666_ _09667_ _08905_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__a21o_1
X_19366_ net5021 _03283_ _03285_ _03275_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_65_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15529_ _08608_ _08623_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18317_ net6331 net3631 _02476_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
X_19297_ net1538 _03238_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7607 rbzero.spi_registers.texadd1\[14\] vssd1 vssd1 vccd1 vccd1 net8134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7618 rbzero.row_render.texu\[1\] vssd1 vssd1 vccd1 vccd1 net8145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7629 rbzero.map_overlay.i_othery\[3\] vssd1 vssd1 vccd1 vccd1 net8156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18248_ _02462_ net3926 net4782 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_4
Xhold6906 net3089 vssd1 vssd1 vccd1 vccd1 net7433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6917 _03018_ vssd1 vssd1 vccd1 vccd1 net7444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6928 net2903 vssd1 vssd1 vccd1 vccd1 net7455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6939 _03054_ vssd1 vssd1 vccd1 vccd1 net7466 sky130_fd_sc_hd__dlygate4sd3_1
X_18179_ net3751 net4435 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold502 net4266 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 net6139 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20210_ net5476 _03743_ _03764_ _03765_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__o211a_1
Xhold524 net5441 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03868_ _03868_ vssd1 vssd1 vccd1 vccd1 clknet_0__03868_ sky130_fd_sc_hd__clkbuf_16
X_21190_ clknet_leaf_129_i_clk net3209 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold535 _03135_ vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 net6173 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 net6169 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20141_ rbzero.debug_overlay.facingX\[-2\] _03711_ vssd1 vssd1 vccd1 vccd1 _03722_
+ sky130_fd_sc_hd__or2_1
Xhold568 net6099 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 net8140 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20072_ _08214_ _03610_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__nor2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _00749_ vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _04297_ vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 rbzero.pov.spi_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 net6747 vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 net6941 vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1257 _01367_ vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1268 net6360 vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1279 net6594 vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
X_20406__157 clknet_1_0__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__inv_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20974_ clknet_leaf_110_i_clk net4166 vssd1 vssd1 vccd1 vccd1 reg_rgb\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21526_ clknet_leaf_19_i_clk net1525 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21457_ clknet_leaf_25_i_clk net3377 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ net6675 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12190_ net4163 _05377_ _04656_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a21o_1
X_21388_ clknet_leaf_20_i_clk net4990 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11141_ net6748 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
X_20339_ clknet_1_0__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__clkbuf_4
X_11072_ net2240 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3160 net7639 vssd1 vssd1 vccd1 vccd1 net3687 sky130_fd_sc_hd__dlygate4sd3_1
X_14900_ net4541 _08034_ _08036_ net4565 net4571 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__o221a_1
Xhold3171 _00646_ vssd1 vssd1 vccd1 vccd1 net3698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22009_ net451 net1847 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _08920_ _08927_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__nor2_1
Xhold3182 net7675 vssd1 vssd1 vccd1 vccd1 net3709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3193 net7741 vssd1 vssd1 vccd1 vccd1 net3720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2470 _04221_ vssd1 vssd1 vccd1 vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2481 rbzero.pov.spi_buffer\[67\] vssd1 vssd1 vccd1 vccd1 net3008 sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ net8354 _07921_ _07928_ net7794 net7806 vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__a221o_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2492 net1856 vssd1 vssd1 vccd1 vccd1 net3019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03857_ clknet_0__03857_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03857_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1780 net5674 vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _08799_ _09664_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nor2_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1791 net2660 vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
X_14762_ net7833 _07922_ _07928_ net7824 net4704 vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__a221o_2
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11974_ net3677 _05080_ _05103_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1
+ vccd1 _05163_ sky130_fd_sc_hd__a22o_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _09497_ _09465_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__or2b_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _06777_ _06786_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__or2_1
X_17481_ _01721_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__or2_1
X_10925_ net2617 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14693_ _07821_ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16432_ _08244_ _08430_ _09392_ _09394_ _09395_ vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__a32o_1
X_19220_ net5444 _03167_ _03198_ _03189_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _06683_ _06737_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__and2_4
X_10856_ net6293 net3104 _04238_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ net836 _03146_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or2_1
X_16363_ _09330_ _09331_ _09328_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ net582 _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__nor2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ net6456 net7210 _04205_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
X_18102_ _02334_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__clkbuf_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ net3532 _08119_ _08162_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__o21a_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ net46 net6792 _03109_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
X_12526_ net43 _05701_ _05699_ net46 _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a221o_1
X_16294_ _09260_ _09263_ _09259_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18033_ net8008 _09540_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15245_ _08330_ _08332_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12457_ net9 _05638_ net5 net6 vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and4b_1
XFILLER_0_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11408_ net7562 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__clkbuf_4
X_20511__252 clknet_1_0__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__inv_2
X_15176_ net4630 _08137_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__nor2_1
X_12388_ rbzero.tex_b1\[15\] rbzero.tex_b1\[14\] _04951_ vssd1 vssd1 vccd1 vccd1 _05573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _07285_ _07297_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ _04523_ _04528_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__a21o_1
X_19984_ net3221 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ _07135_ _07186_ _07227_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__a21o_1
X_18935_ net2934 net7481 _03025_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ net4500 _06169_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18866_ net6661 net7003 _02993_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17817_ net4655 net4756 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18797_ net4709 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19747__29 clknet_1_1__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
X_17748_ _01985_ _01986_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17679_ _09272_ _10346_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19418_ _04459_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__buf_4
X_20690_ net777 net4968 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19349_ net6409 _03271_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7404 net4505 vssd1 vssd1 vccd1 vccd1 net7931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7415 net3472 vssd1 vssd1 vccd1 vccd1 net7942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7426 rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 net7953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7437 net4609 vssd1 vssd1 vccd1 vccd1 net7964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6703 net2018 vssd1 vssd1 vccd1 vccd1 net7230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7448 rbzero.wall_tracer.trackDistX\[2\] vssd1 vssd1 vccd1 vccd1 net7975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6714 rbzero.tex_b0\[56\] vssd1 vssd1 vccd1 vccd1 net7241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7459 net4664 vssd1 vssd1 vccd1 vccd1 net7986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6725 net2592 vssd1 vssd1 vccd1 vccd1 net7252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21311_ clknet_leaf_7_i_clk net5234 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6736 _04189_ vssd1 vssd1 vccd1 vccd1 net7263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6747 rbzero.tex_g1\[51\] vssd1 vssd1 vccd1 vccd1 net7274 sky130_fd_sc_hd__dlygate4sd3_1
X_11462__1 clknet_4_9__leaf_i_clk vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
Xhold6758 net2143 vssd1 vssd1 vccd1 vccd1 net7285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6769 rbzero.tex_b0\[22\] vssd1 vssd1 vccd1 vccd1 net7296 sky130_fd_sc_hd__dlygate4sd3_1
X_21242_ clknet_leaf_43_i_clk net3818 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold310 _03159_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 net5383 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 net5217 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 net5231 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21173_ clknet_leaf_97_i_clk net1170 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold354 net5198 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 net4847 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold376 net5297 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold387 net5337 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 net6108 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
X_20124_ rbzero.debug_overlay.facingX\[-9\] _03711_ vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20055_ net4021 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 _00707_ vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _02977_ vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _03053_ vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 net6515 vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 _01092_ vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _01275_ vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 net6529 vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 net5785 vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 net6055 vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ clknet_leaf_65_i_clk _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ net7035 net2592 _04160_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__mux2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11690_ net4105 _04867_ _04865_ _04467_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20888_ net4948 net63 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10641_ net6822 net1517 _04127_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13360_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__buf_6
X_10572_ net2324 net6898 _04086_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12311_ _05491_ _05493_ _05496_ _04919_ net84 vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21509_ clknet_leaf_48_i_clk net1693 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20569__304 clknet_1_1__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__inv_2
XFILLER_0_146_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13291_ _06327_ _06446_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__xnor2_2
Xhold7971 _08370_ vssd1 vssd1 vccd1 vccd1 net8498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ net4351 _08124_ _06119_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__a21o_1
Xhold7993 _09451_ vssd1 vssd1 vccd1 vccd1 net8520 sky130_fd_sc_hd__dlygate4sd3_1
X_12242_ _04832_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04923_ vssd1 vssd1 vccd1 vccd1 _05361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ net5682 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16981_ _09888_ _10002_ vssd1 vssd1 vccd1 vccd1 _10003_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18720_ _02849_ _02853_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nand3_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ net6526 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
X_15932_ _08402_ _08411_ _08430_ net7836 vssd1 vssd1 vccd1 vccd1 _09027_ sky130_fd_sc_hd__a2bb2o_1
X_15863_ _08341_ _08905_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__nor2_1
X_18651_ _04490_ _02806_ _02807_ _09736_ rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a32o_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _01841_ _01842_ _06057_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__o21ai_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14814_ net8354 _07970_ _07973_ net7824 _07974_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__a221o_4
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _08829_ _08848_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18582_ net7705 _02744_ net91 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_101 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_101/HI o_rgb[10]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_112 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_112/HI zeros[1] sky130_fd_sc_hd__conb_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_123 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_123/HI zeros[12]
+ sky130_fd_sc_hd__conb_1
X_17533_ _01771_ _01772_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__and2_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ net7787 vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__clkbuf_4
Xtop_ew_algofoogle_134 vssd1 vssd1 vccd1 vccd1 ones[7] top_ew_algofoogle_134/LO sky130_fd_sc_hd__conb_1
XFILLER_0_157_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net3927 _05093_ _05095_ rbzero.debug_overlay.facingY\[-3\] _05145_ vssd1
+ vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net7169 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__clkbuf_1
X_17464_ _01680_ _01705_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14676_ _07843_ _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__nand2_1
X_11888_ net4132 _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16415_ _09249_ _09254_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19203_ net6520 _03183_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13627_ _06576_ _06771_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__nor2_1
X_10839_ net6034 net7043 _04227_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
X_17395_ _09915_ _09116_ _10411_ vssd1 vssd1 vccd1 vccd1 _10413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16346_ _09271_ _09310_ _09437_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_172_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19134_ net4369 _03145_ net1177 _03149_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__o211a_1
X_13558_ net555 vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19065_ net3770 net3793 _03104_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
X_12509_ net14 net13 vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__and2b_1
X_16277_ _09342_ _09368_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13489_ _06529_ _06535_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5309 _03618_ vssd1 vssd1 vccd1 vccd1 net5836 sky130_fd_sc_hd__dlygate4sd3_1
X_15228_ _08322_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18016_ _02158_ _02159_ _02233_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_2__f_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4608 net774 vssd1 vssd1 vccd1 vccd1 net5135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4619 _00819_ vssd1 vssd1 vccd1 vccd1 net5146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15159_ net4630 _08137_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__or2_2
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3907 net7788 vssd1 vssd1 vccd1 vccd1 net4434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3918 net3340 vssd1 vssd1 vccd1 vccd1 net4445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3929 _01178_ vssd1 vssd1 vccd1 vccd1 net4456 sky130_fd_sc_hd__dlygate4sd3_1
X_19967_ net5764 net6327 net2312 vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18918_ net3293 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
X_19898_ net6731 net2934 _03550_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18849_ net3695 _02986_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21860_ net302 net1975 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20811_ _03975_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21791_ net233 net1413 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20742_ net5376 _03877_ _03874_ _03918_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20338__96 clknet_1_0__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__inv_2
XFILLER_0_169_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20518__258 clknet_1_1__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__inv_2
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7201 rbzero.spi_registers.got_new_vinf vssd1 vssd1 vccd1 vccd1 net7728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7212 rbzero.debug_overlay.vplaneY\[-4\] vssd1 vssd1 vccd1 vccd1 net7739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7223 rbzero.spi_registers.spi_buffer\[5\] vssd1 vssd1 vccd1 vccd1 net7750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6500 net1930 vssd1 vssd1 vccd1 vccd1 net7027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7245 _09578_ vssd1 vssd1 vccd1 vccd1 net7772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6511 rbzero.tex_b1\[40\] vssd1 vssd1 vccd1 vccd1 net7038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7256 net8369 vssd1 vssd1 vccd1 vccd1 net7783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6522 net2399 vssd1 vssd1 vccd1 vccd1 net7049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7267 _07989_ vssd1 vssd1 vccd1 vccd1 net7794 sky130_fd_sc_hd__buf_2
Xhold6533 _04418_ vssd1 vssd1 vccd1 vccd1 net7060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7278 net550 vssd1 vssd1 vccd1 vccd1 net7805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6544 net2217 vssd1 vssd1 vccd1 vccd1 net7071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7289 net4890 vssd1 vssd1 vccd1 vccd1 net7816 sky130_fd_sc_hd__buf_1
Xhold6555 rbzero.pov.ready_buffer\[43\] vssd1 vssd1 vccd1 vccd1 net7082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5810 net1423 vssd1 vssd1 vccd1 vccd1 net6337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5821 _03475_ vssd1 vssd1 vccd1 vccd1 net6348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6566 net779 vssd1 vssd1 vccd1 vccd1 net7093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5832 net1794 vssd1 vssd1 vccd1 vccd1 net6359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6577 rbzero.tex_g1\[39\] vssd1 vssd1 vccd1 vccd1 net7104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6588 net2165 vssd1 vssd1 vccd1 vccd1 net7115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5843 net1453 vssd1 vssd1 vccd1 vccd1 net6370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6599 _04438_ vssd1 vssd1 vccd1 vccd1 net7126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5854 _02499_ vssd1 vssd1 vccd1 vccd1 net6381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 net5034 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ clknet_leaf_23_i_clk net3268 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5865 rbzero.spi_registers.new_texadd\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net6392
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5876 net1332 vssd1 vssd1 vccd1 vccd1 net6403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net6040 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 net5056 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5887 _03523_ vssd1 vssd1 vccd1 vccd1 net6414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net5030 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5898 rbzero.spi_registers.new_texadd\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net6425
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 net5080 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ clknet_leaf_122_i_clk net3938 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold195 net5130 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
X_20107_ net3473 _03662_ net4375 _03316_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21087_ clknet_leaf_12_i_clk net1424 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20038_ net4454 _03485_ _03609_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ net4044 _06028_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__or2_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11811_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _04978_ vssd1 vssd1 vccd1 vccd1 _05001_
+ sky130_fd_sc_hd__mux2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _05965_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__or2b_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ net431 net2320 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _07699_ _07700_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__xnor2_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _04930_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__or2_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14461_ _07614_ _07612_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__nand2_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _04861_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16200_ _08905_ _09292_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ _06461_ _06558_ _06534_ _06491_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__a211o_1
X_10624_ net7369 net2610 _04116_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__mux2_1
X_17180_ _10070_ _10071_ vssd1 vssd1 vccd1 vccd1 _10200_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14392_ _07308_ _07193_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _06124_ net4908 vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ _06479_ _06512_ _06475_ _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10555_ _04030_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16062_ _08880_ _08391_ _08403_ _08418_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__or4_1
Xhold7790 net3391 vssd1 vssd1 vccd1 vccd1 net8317 sky130_fd_sc_hd__dlygate4sd3_1
X_13274_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xnor2_1
X_10486_ net6880 net7268 _04042_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15013_ _08038_ net4012 vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__and2_1
X_12225_ net88 _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ net3329 net3351 _03517_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__mux2_1
X_12156_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _04912_ vssd1 vssd1 vccd1 vccd1 _05344_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11107_ net6637 net7097 _04375_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16964_ _09963_ _09984_ _09985_ vssd1 vssd1 vccd1 vccd1 _09986_ sky130_fd_sc_hd__and3_1
X_12087_ _04930_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_194_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18703_ net8241 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__clkbuf_4
X_11038_ net2938 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
X_15915_ _09008_ _09009_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__nor2_1
X_20623__353 clknet_1_1__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__inv_2
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19683_ _03456_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__buf_4
X_16895_ _08338_ _09915_ _09636_ _09916_ vssd1 vssd1 vccd1 vccd1 _09917_ sky130_fd_sc_hd__o31ai_1
X_18634_ net3677 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__clkbuf_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _08906_ _08940_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ net3961 _06104_ _10260_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
X_15777_ _08870_ _08871_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__or2b_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ net3945 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ _09249_ _10289_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14728_ _07841_ _07852_ _07896_ net7813 vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__o211a_1
X_18496_ _02626_ net4554 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__or2_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17447_ _10348_ _01682_ _01687_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ _07827_ _07829_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17378_ _09373_ net4914 vssd1 vssd1 vccd1 vccd1 _10396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19117_ net5535 _03126_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__or2_1
X_16329_ _09418_ _09420_ vssd1 vssd1 vccd1 vccd1 _09421_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5106 rbzero.tex_b1\[33\] vssd1 vssd1 vccd1 vccd1 net5633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5117 rbzero.tex_r1\[33\] vssd1 vssd1 vccd1 vccd1 net5644 sky130_fd_sc_hd__dlygate4sd3_1
X_19048_ net7621 net7589 net3398 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
Xhold5128 net2135 vssd1 vssd1 vccd1 vccd1 net5655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5139 net2379 vssd1 vssd1 vccd1 vccd1 net5666 sky130_fd_sc_hd__buf_1
XFILLER_0_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4405 net595 vssd1 vssd1 vccd1 vccd1 net4932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4416 rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 net4943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4427 net607 vssd1 vssd1 vccd1 vccd1 net4954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4438 _00887_ vssd1 vssd1 vccd1 vccd1 net4965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3704 _00900_ vssd1 vssd1 vccd1 vccd1 net4231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4449 net705 vssd1 vssd1 vccd1 vccd1 net4976 sky130_fd_sc_hd__dlygate4sd3_1
X_21010_ clknet_leaf_38_i_clk net4273 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3726 rbzero.wall_tracer.visualWallDist\[3\] vssd1 vssd1 vccd1 vccd1 net4253 sky130_fd_sc_hd__buf_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3737 net1039 vssd1 vssd1 vccd1 vccd1 net4264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3748 net8030 vssd1 vssd1 vccd1 vccd1 net4275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3759 net2398 vssd1 vssd1 vccd1 vccd1 net4286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19803__80 clknet_1_1__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__inv_2
X_21912_ net354 net2687 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
X_20598__330 clknet_1_0__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__inv_2
XFILLER_0_179_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21843_ net285 net2547 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21774_ clknet_leaf_48_i_clk net1443 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20725_ _03899_ _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7020 rbzero.pov.ready_buffer\[24\] vssd1 vssd1 vccd1 vccd1 net7547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7031 net2709 vssd1 vssd1 vccd1 vccd1 net7558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7042 net4450 vssd1 vssd1 vccd1 vccd1 net7569 sky130_fd_sc_hd__buf_1
Xhold7053 _03101_ vssd1 vssd1 vccd1 vccd1 net7580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7064 net3557 vssd1 vssd1 vccd1 vccd1 net7591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6330 rbzero.spi_registers.new_mapd\[14\] vssd1 vssd1 vccd1 vccd1 net6857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7075 _03103_ vssd1 vssd1 vccd1 vccd1 net7602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6341 net1909 vssd1 vssd1 vccd1 vccd1 net6868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7086 net3080 vssd1 vssd1 vccd1 vccd1 net7613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6352 rbzero.tex_r1\[46\] vssd1 vssd1 vccd1 vccd1 net6879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7097 net3881 vssd1 vssd1 vccd1 vccd1 net7624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6363 net2536 vssd1 vssd1 vccd1 vccd1 net6890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6374 rbzero.tex_r1\[59\] vssd1 vssd1 vccd1 vccd1 net6901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5640 rbzero.tex_g1\[28\] vssd1 vssd1 vccd1 vccd1 net6167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6385 net2245 vssd1 vssd1 vccd1 vccd1 net6912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6396 rbzero.tex_g0\[46\] vssd1 vssd1 vccd1 vccd1 net6923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5651 net1387 vssd1 vssd1 vccd1 vccd1 net6178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5662 net1143 vssd1 vssd1 vccd1 vccd1 net6189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5673 rbzero.pov.spi_buffer\[53\] vssd1 vssd1 vccd1 vccd1 net6200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5684 net1173 vssd1 vssd1 vccd1 vccd1 net6211 sky130_fd_sc_hd__dlygate4sd3_1
X_12010_ _04736_ _05189_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__and3b_1
Xhold5695 rbzero.tex_g1\[5\] vssd1 vssd1 vccd1 vccd1 net6222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4950 _01229_ vssd1 vssd1 vccd1 vccd1 net5477 sky130_fd_sc_hd__dlygate4sd3_1
X_21208_ clknet_leaf_127_i_clk net1147 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4961 net1217 vssd1 vssd1 vccd1 vccd1 net5488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4972 rbzero.spi_registers.new_leak\[3\] vssd1 vssd1 vccd1 vccd1 net5499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4983 _00884_ vssd1 vssd1 vccd1 vccd1 net5510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4994 rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 net5521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21139_ clknet_leaf_95_i_clk net3528 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_4
X_13961_ _07100_ _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15700_ _08794_ _08781_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__xnor2_1
X_12912_ net4705 net4718 net4751 net4757 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__or4_1
X_16680_ net5596 _09741_ _09742_ net4769 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
X_13892_ _07006_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15631_ _08690_ _08701_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__xnor2_4
X_12843_ _05948_ _05976_ _06017_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__and3_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15562_ _08646_ _08647_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_189_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18350_ net5961 _02535_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12774_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__and2_2
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _10163_ net8008 _10318_ vssd1 vssd1 vccd1 vccd1 _10320_ sky130_fd_sc_hd__o21ai_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _07669_ _07670_ _07683_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__a21o_1
X_11725_ _04831_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__buf_4
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _08580_ _08582_ _08579_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18281_ net1420 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17232_ _09891_ _10126_ _10251_ vssd1 vssd1 vccd1 vccd1 _10252_ sky130_fd_sc_hd__a21oi_2
X_14444_ _07612_ _07613_ _07614_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_182_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11656_ _04796_ _04814_ _04830_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nor3_1
Xclkbuf_1_1__f__03870_ clknet_0__03870_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03870_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10607_ net7141 net6187 _04105_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__mux2_1
X_17163_ _10067_ _10076_ _10075_ vssd1 vssd1 vccd1 vccd1 _10183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14375_ _07492_ _07538_ _07541_ _07543_ _07545_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__a32oi_4
X_11587_ net1075 net1658 vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ _09109_ _09207_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__xor2_4
XFILLER_0_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13326_ _06343_ _06404_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nand2_2
X_17094_ _09988_ _09989_ vssd1 vssd1 vccd1 vccd1 _10115_ sky130_fd_sc_hd__nor2_1
X_10538_ net2174 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold909 _02494_ vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16045_ _09137_ _09138_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ _06420_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__inv_2
X_10469_ net2131 net6689 _04031_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _04950_ vssd1 vssd1 vccd1 vccd1 _05395_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13188_ _06269_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12139_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _04837_ vssd1 vssd1 vccd1 vccd1 _05327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17996_ _02062_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__xnor2_1
Xhold1609 _01338_ vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19735_ net7649 net2310 net3922 vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__and3b_1
X_16947_ net4622 _06123_ vssd1 vssd1 vccd1 vccd1 _09969_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19666_ net1311 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
X_16878_ _08543_ _09472_ vssd1 vssd1 vccd1 vccd1 _09900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18617_ _02526_ _02769_ _02770_ _02775_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a32o_1
X_15829_ _08878_ _08883_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19597_ net1778 net887 _03312_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18548_ net5935 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18479_ _02626_ net3494 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21490_ clknet_leaf_8_i_clk net1925 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20372_ clknet_1_1__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__buf_1
XFILLER_0_71_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22111_ clknet_leaf_89_i_clk net4924 vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4213 net3296 vssd1 vssd1 vccd1 vccd1 net4740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4224 net4247 vssd1 vssd1 vccd1 vccd1 net4751 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4235 net3943 vssd1 vssd1 vccd1 vccd1 net4762 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3501 net1395 vssd1 vssd1 vccd1 vccd1 net4028 sky130_fd_sc_hd__dlygate4sd3_1
X_22042_ net484 net1844 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold4246 net8028 vssd1 vssd1 vccd1 vccd1 net4773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3512 _02485_ vssd1 vssd1 vccd1 vccd1 net4039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4257 _02561_ vssd1 vssd1 vccd1 vccd1 net4784 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4268 net1610 vssd1 vssd1 vccd1 vccd1 net4795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3523 _02746_ vssd1 vssd1 vccd1 vccd1 net4050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3534 rbzero.spi_registers.ss_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net4061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2800 net4903 vssd1 vssd1 vccd1 vccd1 net3327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3545 _01250_ vssd1 vssd1 vccd1 vccd1 net4072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2811 net5985 vssd1 vssd1 vccd1 vccd1 net3338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3556 net3773 vssd1 vssd1 vccd1 vccd1 net4083 sky130_fd_sc_hd__buf_2
Xhold2822 net5838 vssd1 vssd1 vccd1 vccd1 net3349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3567 net4159 vssd1 vssd1 vccd1 vccd1 net4094 sky130_fd_sc_hd__clkbuf_1
Xhold3578 net5910 vssd1 vssd1 vccd1 vccd1 net4105 sky130_fd_sc_hd__buf_2
Xhold2833 net4753 vssd1 vssd1 vccd1 vccd1 net3360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3589 _05061_ vssd1 vssd1 vccd1 vccd1 net4116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2844 net5888 vssd1 vssd1 vccd1 vccd1 net3371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 net8345 vssd1 vssd1 vccd1 vccd1 net3382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2866 net4552 vssd1 vssd1 vccd1 vccd1 net3393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2877 _00730_ vssd1 vssd1 vccd1 vccd1 net3404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2888 _03672_ vssd1 vssd1 vccd1 vccd1 net3415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2899 net7877 vssd1 vssd1 vccd1 vccd1 net3426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21826_ net268 net1187 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21757_ clknet_leaf_84_i_clk net4104 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_1
X_20375__129 clknet_1_0__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__inv_2
XFILLER_0_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20708_ net754 net5400 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ net4110 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21688_ clknet_leaf_114_i_clk net5829 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ rbzero.spi_registers.texadd2\[2\] _04506_ _04632_ vssd1 vssd1 vccd1 vccd1
+ _04633_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_184_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _07328_ _07330_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__and2b_1
X_11372_ _04561_ _04562_ _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13111_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
Xhold6160 net616 vssd1 vssd1 vccd1 vccd1 net6687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6171 rbzero.tex_b1\[24\] vssd1 vssd1 vccd1 vccd1 net6698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6182 net1876 vssd1 vssd1 vccd1 vccd1 net6709 sky130_fd_sc_hd__dlygate4sd3_1
X_14091_ net580 _07249_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__nand2_1
Xhold6193 _04207_ vssd1 vssd1 vccd1 vccd1 net6720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5470 _03348_ vssd1 vssd1 vccd1 vccd1 net5997 sky130_fd_sc_hd__dlygate4sd3_1
X_13042_ _06213_ net3811 _06217_ net3766 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__o22a_1
Xhold5481 _03351_ vssd1 vssd1 vccd1 vccd1 net6008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5492 net1480 vssd1 vssd1 vccd1 vccd1 net6019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4780 rbzero.spi_registers.texadd1\[18\] vssd1 vssd1 vccd1 vccd1 net5307 sky130_fd_sc_hd__dlygate4sd3_1
X_17850_ _02085_ _02087_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4791 net875 vssd1 vssd1 vccd1 vccd1 net5318 sky130_fd_sc_hd__dlygate4sd3_1
X_16801_ _09827_ _09828_ _09829_ vssd1 vssd1 vccd1 vccd1 _09830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_195_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17781_ _09040_ net8008 _02018_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__o21ai_1
X_14993_ _08093_ net4149 vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19520_ net1494 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
X_16732_ _09765_ _09766_ _09768_ _09769_ net5554 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__a32o_1
X_13944_ _07107_ _07113_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19451_ net1658 _03334_ net5514 _03299_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13875_ net77 _06708_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__nor2_1
X_16663_ net4246 _09737_ _09740_ _07917_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__a22o_1
X_18402_ net4725 net8074 _02583_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15614_ net7836 _08204_ _08205_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__and3_1
X_12826_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__and2_1
X_19382_ net6317 _03284_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__or2_1
X_16594_ _09671_ _09682_ _09683_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__nand3_1
XFILLER_0_146_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18333_ _02520_ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15545_ _08636_ _08637_ _08639_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__nand3_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12757_ _05905_ _05932_ _05933_ _05906_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__o211a_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _04894_ _04895_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a21oi_1
X_15476_ _08374_ net4877 _08494_ _08366_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__or4b_2
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18264_ _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__buf_4
X_12688_ net52 _05852_ _05865_ net53 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17215_ _10207_ _10234_ vssd1 vssd1 vccd1 vccd1 _10235_ sky130_fd_sc_hd__nand2_1
X_14427_ _07586_ _07596_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03853_ clknet_0__03853_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03853_
+ sky130_fd_sc_hd__clkbuf_16
X_18195_ _02407_ _02411_ _02414_ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17146_ _08383_ _09062_ _10040_ vssd1 vssd1 vccd1 vccd1 _10166_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ _07459_ _07460_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold706 net5491 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 net6435 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold728 net8143 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13309_ _06473_ _06474_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__and2_1
X_17077_ _09666_ _09667_ _08402_ vssd1 vssd1 vccd1 vccd1 _10098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14289_ _07388_ _07392_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__xnor2_2
Xhold739 net6320 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _08615_ _09063_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2107 _01308_ vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2118 _03410_ vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2129 _01064_ vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1406 _03037_ vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_20480__224 clknet_1_0__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__inv_2
XFILLER_0_97_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1417 net6970 vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 net6765 vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ _02191_ _02215_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__xor2_1
Xhold1439 _01390_ vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19718_ net5280 net7273 net2310 vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o21ai_1
X_20990_ clknet_leaf_110_i_clk net4109 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19649_ net6727 net3866 _03441_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21611_ clknet_leaf_133_i_clk net2871 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21542_ net176 net2834 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21473_ clknet_leaf_23_i_clk net1639 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4010 net3723 vssd1 vssd1 vccd1 vccd1 net4537 sky130_fd_sc_hd__clkbuf_2
Xhold4021 _00418_ vssd1 vssd1 vccd1 vccd1 net4548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4032 net672 vssd1 vssd1 vccd1 vccd1 net4559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4054 net3796 vssd1 vssd1 vccd1 vccd1 net4581 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20286_ net6552 net4028 _03814_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__mux2_1
Xhold3320 net3384 vssd1 vssd1 vccd1 vccd1 net3847 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_179_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4065 _01230_ vssd1 vssd1 vccd1 vccd1 net4592 sky130_fd_sc_hd__dlygate4sd3_1
X_22025_ net467 net2995 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
Xhold4076 net8259 vssd1 vssd1 vccd1 vccd1 net4603 sky130_fd_sc_hd__buf_2
Xhold3331 _04663_ vssd1 vssd1 vccd1 vccd1 net3858 sky130_fd_sc_hd__buf_1
Xhold3342 net7978 vssd1 vssd1 vccd1 vccd1 net3869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4087 rbzero.row_render.size\[7\] vssd1 vssd1 vccd1 vccd1 net4614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3364 net5891 vssd1 vssd1 vccd1 vccd1 net3891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2630 _01105_ vssd1 vssd1 vccd1 vccd1 net3157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3375 net5939 vssd1 vssd1 vccd1 vccd1 net3902 sky130_fd_sc_hd__clkbuf_2
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3386 net8006 vssd1 vssd1 vccd1 vccd1 net3913 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2641 _01128_ vssd1 vssd1 vccd1 vccd1 net3168 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3397 _01019_ vssd1 vssd1 vccd1 vccd1 net3924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2652 net7555 vssd1 vssd1 vccd1 vccd1 net3179 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2663 net5740 vssd1 vssd1 vccd1 vccd1 net3190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2674 _01162_ vssd1 vssd1 vccd1 vccd1 net3201 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1940 _01557_ vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2685 _01087_ vssd1 vssd1 vccd1 vccd1 net3212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 net4927 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1951 _01404_ vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net4939 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net4945 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2696 net3311 vssd1 vssd1 vccd1 vccd1 net3223 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net4176 _04460_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__xor2_1
Xhold1962 net7378 vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold99 net5585 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1973 _04054_ vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 _01317_ vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ net7071 net2300 _04287_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__mux2_1
Xhold1995 _04224_ vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13660_ _06771_ _06829_ _06830_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__o21a_1
X_10872_ net2686 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ net21 net20 _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__or3b_2
X_21809_ net251 net2696 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _06575_ _06702_ _06754_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _04511_ _06370_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__nand2_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12542_ _04494_ _05700_ _05698_ _04500_ _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15261_ _08168_ _08221_ _08246_ _08186_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12473_ net4133 net4089 _05633_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17000_ _09927_ _10019_ _10020_ vssd1 vssd1 vccd1 vccd1 _10021_ sky130_fd_sc_hd__a21oi_4
X_14212_ _07334_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ _04540_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and2_1
X_15192_ _08144_ _08286_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__and2_2
XFILLER_0_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 _05743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14143_ _07033_ net569 vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11355_ _04513_ _04543_ _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ _07183_ _07226_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__nand2_2
X_18951_ net2839 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11286_ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13025_ net4581 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__inv_2
X_17902_ _02138_ _02139_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__nor2_1
X_18882_ net1195 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17833_ _02026_ _02028_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17764_ _09272_ _02002_ _01922_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_2
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14976_ net4653 _08017_ _08079_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19503_ net1493 net6844 _03365_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16715_ net3999 _09102_ vssd1 vssd1 vccd1 vccd1 _09753_ sky130_fd_sc_hd__or2_1
X_13927_ _06911_ _06997_ _07094_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_199_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17695_ _01891_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19434_ net4960 _03323_ _03326_ _03316_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__a211o_1
X_16646_ net3517 net4124 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13858_ _07028_ _07027_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__or2b_4
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _05980_ _05983_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a21oi_2
X_19365_ net1474 _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or2_1
X_16577_ net3934 _06123_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__nand2_2
X_13789_ _06954_ _06958_ _06959_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ net6162 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__clkbuf_1
X_15528_ _08621_ _08622_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__nor2_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19296_ net5216 _03236_ _03244_ _03230_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__o211a_1
Xhold7608 net4207 vssd1 vssd1 vccd1 vccd1 net8135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7619 rbzero.row_render.texu\[3\] vssd1 vssd1 vccd1 vccd1 net8146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ _02238_ _02239_ _02461_ _02245_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
X_15459_ _08255_ _08323_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6907 _04286_ vssd1 vssd1 vccd1 vccd1 net7434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6918 net3183 vssd1 vssd1 vccd1 vccd1 net7445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6929 rbzero.tex_r1\[31\] vssd1 vssd1 vccd1 vccd1 net7456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ net3751 net4435 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold503 net8194 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_1
X_17129_ _09249_ net4909 vssd1 vssd1 vccd1 vccd1 _10149_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold514 net6141 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold525 net6155 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03867_ _03867_ vssd1 vssd1 vccd1 vccd1 clknet_0__03867_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold536 net4325 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _01513_ vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _01433_ vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ net3609 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold569 net6101 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ net3372 _03660_ net5751 _03628_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__o211a_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 net6672 vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _01360_ vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1225 net1706 vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1236 _01079_ vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 net6943 vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1258 net6600 vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _01470_ vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20973_ clknet_leaf_111_i_clk net4143 vssd1 vssd1 vccd1 vccd1 reg_rgb\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21525_ clknet_leaf_20_i_clk net2139 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21456_ clknet_leaf_19_i_clk net1884 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21387_ clknet_leaf_3_i_clk net5199 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11140_ net6746 net1819 _04390_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 o_gpout[0] sky130_fd_sc_hd__buf_1
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__clkbuf_4
X_11071_ net6128 net2239 _04353_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__mux2_1
X_20269_ net4098 net4179 _09725_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and3b_1
Xhold3150 rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 net3677 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22008_ net450 net2627 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold3161 _03730_ vssd1 vssd1 vccd1 vccd1 net3688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3172 net7841 vssd1 vssd1 vccd1 vccd1 net3699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3183 _01018_ vssd1 vssd1 vccd1 vccd1 net3710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3194 _03725_ vssd1 vssd1 vccd1 vccd1 net3721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2460 net7404 vssd1 vssd1 vccd1 vccd1 net2987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2471 _01429_ vssd1 vssd1 vccd1 vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
X_14830_ net7793 vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__clkbuf_2
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2482 net1567 vssd1 vssd1 vccd1 vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2493 _03002_ vssd1 vssd1 vccd1 vccd1 net3020 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03856_ clknet_0__03856_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03856_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1770 net6887 vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1781 _01292_ vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11973_ rbzero.debug_overlay.vplaneY\[0\] _05093_ _05095_ rbzero.debug_overlay.vplaneY\[-3\]
+ _05161_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
X_14761_ net7846 _07926_ _07927_ net7785 vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__o211a_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1792 _04168_ vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _09574_ _09462_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__or2b_1
XFILLER_0_168_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ net7190 net6072 _04276_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__inv_2
X_17480_ _01718_ _01720_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__and2_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _07732_ _07862_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16431_ _09500_ _09521_ vssd1 vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__xnor2_1
X_10855_ net5702 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__clkbuf_1
X_13643_ _06813_ net540 vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ net4384 _03145_ net2067 _03149_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ _06742_ _06743_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__xnor2_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _09452_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__and2b_1
X_10786_ net2472 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18101_ _02333_ net3932 _02320_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ net13 net12 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__or2_1
X_15313_ net3453 _08405_ _08407_ _08133_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__a211o_2
X_16293_ _09383_ _09384_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__xnor2_2
X_19081_ net3033 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__clkbuf_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18032_ _02172_ _02179_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15244_ _08338_ _08139_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__nor2_2
X_12456_ _05634_ _05636_ _05637_ net8 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _04494_ _04572_ _04585_ _04590_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__o32a_2
X_15175_ _08244_ _08245_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__nand2_1
X_12387_ _05517_ _05569_ _05571_ _05306_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _07294_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__xnor2_1
X_11338_ _04521_ _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__nand2_1
X_19983_ net7502 net7425 _08092_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_132_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14057_ _07135_ _07186_ _07227_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__nand3_1
X_18934_ net6733 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
X_11269_ net4057 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ _06179_ net3847 net4565 _06177_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a22o_1
X_18865_ net1574 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ _02054_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__clkbuf_1
X_18796_ _02940_ _02941_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__xnor2_1
X_17747_ _10186_ _09114_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nor2_1
X_14959_ net4776 _07962_ _08068_ vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__mux2_1
X_17678_ _01808_ _01811_ _01809_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19417_ net2321 net3902 _03141_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__and3_1
X_20592__325 clknet_1_0__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__inv_2
X_16629_ _04665_ net4121 _09717_ vssd1 vssd1 vccd1 vccd1 _09718_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19348_ net5193 _03269_ _03274_ _03275_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7427 net4525 vssd1 vssd1 vccd1 vccd1 net7954 sky130_fd_sc_hd__dlygate4sd3_1
X_19279_ net5089 _03200_ _03233_ _03230_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__o211a_1
Xhold7438 rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 net7965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6704 rbzero.tex_g0\[27\] vssd1 vssd1 vccd1 vccd1 net7231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7449 net4656 vssd1 vssd1 vccd1 vccd1 net7976 sky130_fd_sc_hd__dlygate4sd3_1
X_21310_ clknet_leaf_9_i_clk net5123 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6715 net2512 vssd1 vssd1 vccd1 vccd1 net7242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6726 rbzero.tex_g0\[9\] vssd1 vssd1 vccd1 vccd1 net7253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6737 net2821 vssd1 vssd1 vccd1 vccd1 net7264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6748 net2518 vssd1 vssd1 vccd1 vccd1 net7275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6759 rbzero.tex_r0\[62\] vssd1 vssd1 vccd1 vccd1 net7286 sky130_fd_sc_hd__dlygate4sd3_1
X_21241_ clknet_leaf_44_i_clk net3879 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold300 net5062 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 net4358 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 net5385 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold333 net5263 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 net5233 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
X_21172_ clknet_leaf_97_i_clk net1196 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold355 net5188 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 net4849 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 net6095 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold388 net5339 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
X_20123_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__buf_2
Xhold399 _01363_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20054_ _03320_ net4020 vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and2_1
Xhold1000 net6549 vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 net6491 vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 net5880 vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1033 _00701_ vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 net6517 vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 net5512 vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 net6049 vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _00590_ vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _00720_ vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _03358_ vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ clknet_leaf_78_i_clk _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _03312_ net1096 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net2044 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10571_ net6609 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ _05494_ _05495_ _04976_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21508_ clknet_leaf_45_i_clk net1418 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13290_ _06350_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__xnor2_4
X_12241_ rbzero.tex_g1\[47\] rbzero.tex_g1\[46\] _04836_ vssd1 vssd1 vccd1 vccd1 _05428_
+ sky130_fd_sc_hd__mux2_1
X_21439_ clknet_leaf_25_i_clk net1738 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _04915_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11123_ net2351 net5680 _04030_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
X_16980_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10002_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ net1955 net6524 _04342_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
X_15931_ _08401_ _08402_ _08410_ _09025_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_64_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ net3619 _02805_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__nand2_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _08948_ _08691_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2290 net1894 vssd1 vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
X_17601_ _01721_ _01728_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ net7793 _07943_ net3638 vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__a21o_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _09752_ _09762_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__xor2_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _08886_ _08887_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__or2_1
X_20541__279 clknet_1_1__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__inv_2
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_102 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_102/HI o_rgb[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17532_ _01771_ _01772_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_113 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_113/HI zeros[2] sky130_fd_sc_hd__conb_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ net7784 vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_124 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_124/HI zeros[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_197_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11956_ rbzero.debug_overlay.facingY\[-9\] _05106_ _05114_ rbzero.debug_overlay.facingY\[-4\]
+ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a221o_1
Xtop_ew_algofoogle_135 vssd1 vssd1 vccd1 vccd1 ones[8] top_ew_algofoogle_135/LO sky130_fd_sc_hd__conb_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10907_ net7167 net3070 _04265_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__mux2_1
X_17463_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11887_ _04667_ _05075_ net4116 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__o21ba_1
X_14675_ _07841_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__nand2_1
X_19202_ net5121 _03182_ _03188_ _03189_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__o211a_1
X_16414_ _09502_ _09504_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__nand2_1
X_10838_ net2739 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__clkbuf_1
X_13626_ _06693_ _06796_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17394_ _09915_ _09116_ _10411_ vssd1 vssd1 vccd1 vccd1 _10412_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ net1176 _03147_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__or2_1
X_16345_ _09307_ _09309_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__nor2_1
X_10769_ net2552 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__clkbuf_1
X_13557_ _06681_ _06725_ _06726_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _05689_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
X_19064_ _02947_ _02969_ net3395 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__and3_2
XFILLER_0_113_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16276_ _09349_ _09367_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__xor2_2
X_13488_ _06568_ _06567_ net559 vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20435__184 clknet_1_0__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__inv_2
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ net4622 _02249_ _09845_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12439_ _04909_ _05582_ _05616_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a31o_1
X_15227_ _08128_ _08320_ _08321_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__o21a_2
Xclkbuf_leaf_17_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4609 rbzero.spi_registers.texadd2\[9\] vssd1 vssd1 vccd1 vccd1 net5136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ _08252_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__clkbuf_4
Xhold3908 net3532 vssd1 vssd1 vccd1 vccd1 net4435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3919 rbzero.debug_overlay.facingX\[10\] vssd1 vssd1 vccd1 vccd1 net4446 sky130_fd_sc_hd__buf_2
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14109_ _07243_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__xnor2_4
X_19966_ net3238 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
X_15089_ net4392 _08123_ _08148_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18917_ net3342 net7583 _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__mux2_1
X_19897_ net3126 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18848_ net5800 net1251 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18779_ _02925_ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__nand2_1
X_20600__332 clknet_1_1__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__inv_2
X_20810_ net991 net5739 vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__and2_1
X_21790_ clknet_leaf_19_i_clk net1388 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20741_ _03914_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7202 rbzero.color_floor\[0\] vssd1 vssd1 vccd1 vccd1 net7729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7224 net8315 vssd1 vssd1 vccd1 vccd1 net7751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6501 rbzero.tex_g1\[54\] vssd1 vssd1 vccd1 vccd1 net7028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6512 net2509 vssd1 vssd1 vccd1 vccd1 net7039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7257 _06547_ vssd1 vssd1 vccd1 vccd1 net7784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6523 rbzero.tex_g0\[49\] vssd1 vssd1 vccd1 vccd1 net7050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7268 net8443 vssd1 vssd1 vccd1 vccd1 net7795 sky130_fd_sc_hd__clkbuf_2
Xhold6534 net2212 vssd1 vssd1 vccd1 vccd1 net7061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7279 net4703 vssd1 vssd1 vccd1 vccd1 net7806 sky130_fd_sc_hd__buf_1
Xhold6545 _04291_ vssd1 vssd1 vccd1 vccd1 net7072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5800 net1260 vssd1 vssd1 vccd1 vccd1 net6327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6556 net775 vssd1 vssd1 vccd1 vccd1 net7083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5811 rbzero.spi_registers.new_texadd\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net6338
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6567 rbzero.tex_r0\[15\] vssd1 vssd1 vccd1 vccd1 net7094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5822 net1326 vssd1 vssd1 vccd1 vccd1 net6349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5833 _04175_ vssd1 vssd1 vccd1 vccd1 net6360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6578 net2176 vssd1 vssd1 vccd1 vccd1 net7105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5844 rbzero.spi_registers.new_texadd\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net6371
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 net5643 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6589 rbzero.tex_g1\[62\] vssd1 vssd1 vccd1 vccd1 net7116 sky130_fd_sc_hd__dlygate4sd3_1
X_21224_ clknet_leaf_23_i_clk net2865 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5855 net1445 vssd1 vssd1 vccd1 vccd1 net6382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 net4991 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5866 net597 vssd1 vssd1 vccd1 vccd1 net6393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 net6042 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5877 rbzero.spi_registers.new_texadd\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net6404
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5888 net1317 vssd1 vssd1 vccd1 vccd1 net6415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 net5058 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5899 net839 vssd1 vssd1 vccd1 vccd1 net6426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 net5076 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold185 net5082 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
X_21155_ clknet_leaf_122_i_clk net5881 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold196 net5092 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
X_20106_ net4374 _03631_ _03695_ _03696_ _03659_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o221a_1
X_21086_ clknet_leaf_46_i_clk net1398 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20037_ _03642_ _03643_ _03610_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _04984_ _04997_ _04999_ _04988_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__o211a_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__nand2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ net430 net2763 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _04912_ vssd1 vssd1 vccd1 vccd1 _04931_
+ sky130_fd_sc_hd__mux2_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ clknet_leaf_76_i_clk net4693 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _07588_ _07594_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__xnor2_2
X_11672_ net3423 net3365 _04859_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__nor3_1
XFILLER_0_166_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ net5579 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13411_ _06579_ _06581_ _06516_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14391_ _07308_ _07194_ _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16130_ net8068 _08129_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13342_ _06467_ _06468_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__nand2_1
X_10554_ net5661 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16061_ _09027_ _09029_ _09026_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13273_ _06351_ _06404_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__nand2_1
Xhold7780 net4245 vssd1 vssd1 vccd1 vccd1 net8307 sky130_fd_sc_hd__dlygate4sd3_1
X_10485_ net3129 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__clkbuf_1
Xhold7791 rbzero.row_render.size\[4\] vssd1 vssd1 vccd1 vccd1 net8318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _04836_ vssd1 vssd1 vccd1 vccd1 _05411_
+ sky130_fd_sc_hd__mux2_1
X_15012_ _04566_ net4011 _08104_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__mux2_1
X_19820_ net1815 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _04915_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11106_ net7077 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12086_ _04977_ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__or2_1
X_16963_ _09981_ _09982_ _09983_ vssd1 vssd1 vccd1 vccd1 _09985_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18702_ _02840_ _02851_ _02852_ _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a31o_1
X_11037_ net7196 net7344 _04331_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__mux2_1
X_15914_ _09006_ _09007_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__and2_1
X_19682_ net6353 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16894_ _09503_ _09638_ vssd1 vssd1 vccd1 vccd1 _09916_ sky130_fd_sc_hd__or2b_1
XFILLER_0_155_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18633_ _02781_ _02782_ _02783_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _08909_ _08908_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__and2b_1
XFILLER_0_204_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ net3443 net3960 _02245_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
X_15776_ _08161_ net8414 _08279_ _08318_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__or4_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ net4569 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__inv_2
X_17515_ _01754_ _01755_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__nor2_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14727_ _07841_ _07865_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__nand2_1
X_18495_ net8257 _02667_ net4868 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11939_ _05123_ _05125_ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__or3_1
XFILLER_0_185_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ _10348_ _01682_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14658_ _07828_ _07816_ _07812_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13609_ _06575_ _06702_ _06692_ _06753_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__or4_1
X_17377_ _08167_ net4909 vssd1 vssd1 vccd1 vccd1 _10395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ _07758_ _07759_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19116_ net4306 _03125_ net1077 _03128_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ _09419_ _09296_ _08474_ vssd1 vssd1 vccd1 vccd1 _09420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5107 net1949 vssd1 vssd1 vccd1 vccd1 net5634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19047_ net3739 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__clkbuf_1
X_16259_ _06122_ _08612_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__nor2_2
Xhold5118 net2250 vssd1 vssd1 vccd1 vccd1 net5645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5129 rbzero.hsync vssd1 vssd1 vccd1 vccd1 net5656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4406 _01645_ vssd1 vssd1 vccd1 vccd1 net4933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4417 net614 vssd1 vssd1 vccd1 vccd1 net4944 sky130_fd_sc_hd__buf_1
Xhold4428 rbzero.color_floor\[5\] vssd1 vssd1 vccd1 vccd1 net4955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4439 net622 vssd1 vssd1 vccd1 vccd1 net4966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3705 net1367 vssd1 vssd1 vccd1 vccd1 net4232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3716 net7912 vssd1 vssd1 vccd1 vccd1 net4243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3727 net8013 vssd1 vssd1 vccd1 vccd1 net4254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3738 rbzero.wall_tracer.visualWallDist\[9\] vssd1 vssd1 vccd1 vccd1 net4265 sky130_fd_sc_hd__buf_1
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3749 net985 vssd1 vssd1 vccd1 vccd1 net4276 sky130_fd_sc_hd__dlygate4sd3_1
X_19949_ net7520 net7449 _03583_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21911_ net353 net1807 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21842_ net284 net1160 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21773_ clknet_leaf_48_i_clk net1265 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20724_ net5404 _03877_ _03874_ _03903_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7010 rbzero.pov.ready_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net7537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7021 net3289 vssd1 vssd1 vccd1 vccd1 net7548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7032 rbzero.pov.spi_buffer\[55\] vssd1 vssd1 vccd1 vccd1 net7559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7043 _04907_ vssd1 vssd1 vccd1 vccd1 net7570 sky130_fd_sc_hd__buf_2
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7054 net3482 vssd1 vssd1 vccd1 vccd1 net7581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6320 _04366_ vssd1 vssd1 vccd1 vccd1 net6847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7065 rbzero.pov.ready_buffer\[35\] vssd1 vssd1 vccd1 vccd1 net7592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7076 net3632 vssd1 vssd1 vccd1 vccd1 net7603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6331 net1133 vssd1 vssd1 vccd1 vccd1 net6858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6342 _04444_ vssd1 vssd1 vccd1 vccd1 net6869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7087 rbzero.spi_registers.spi_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net7614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6353 net2128 vssd1 vssd1 vccd1 vccd1 net6880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6364 _04380_ vssd1 vssd1 vccd1 vccd1 net6891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5630 _04415_ vssd1 vssd1 vccd1 vccd1 net6157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6375 net2348 vssd1 vssd1 vccd1 vccd1 net6902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6386 rbzero.tex_r0\[41\] vssd1 vssd1 vccd1 vccd1 net6913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5641 net1083 vssd1 vssd1 vccd1 vccd1 net6168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6397 net2035 vssd1 vssd1 vccd1 vccd1 net6924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5652 rbzero.spi_registers.new_texadd\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net6179
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5663 rbzero.spi_registers.new_texadd\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net6190
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21207_ clknet_leaf_116_i_clk net1908 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5674 net1110 vssd1 vssd1 vccd1 vccd1 net6201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5685 _04232_ vssd1 vssd1 vccd1 vccd1 net6212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4940 rbzero.map_overlay.i_mapdy\[5\] vssd1 vssd1 vccd1 vccd1 net5467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5696 net1179 vssd1 vssd1 vccd1 vccd1 net6223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4951 net1109 vssd1 vssd1 vccd1 vccd1 net5478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4962 _01613_ vssd1 vssd1 vccd1 vccd1 net5489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4973 net1634 vssd1 vssd1 vccd1 vccd1 net5500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4984 net1415 vssd1 vssd1 vccd1 vccd1 net5511 sky130_fd_sc_hd__dlygate4sd3_1
X_21138_ clknet_leaf_95_i_clk net3310 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20607__338 clknet_1_0__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__inv_2
Xhold4995 net1284 vssd1 vssd1 vccd1 vccd1 net5522 sky130_fd_sc_hd__dlygate4sd3_1
X_20682__3 clknet_1_0__leaf__03506_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
X_13960_ _07102_ _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__xnor2_2
X_21069_ clknet_leaf_80_i_clk _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12911_ _06080_ _06083_ _06085_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__or4b_1
XFILLER_0_88_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13891_ _07019_ _07018_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__nor2_1
X_15630_ _08715_ _08723_ _08724_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_159_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _05948_ _05976_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a21oi_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _08354_ _08655_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__xnor2_4
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12773_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__nor2_2
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17300_ _10163_ net8008 _10318_ vssd1 vssd1 vccd1 vccd1 _10319_ sky130_fd_sc_hd__or3_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _07672_ _07681_ _07682_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__a21o_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _04913_ vssd1 vssd1 vccd1 vccd1 _04914_
+ sky130_fd_sc_hd__mux2_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18280_ net6390 net2205 _02477_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
X_15492_ _08247_ _08267_ _08242_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__a21bo_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17231_ _10123_ _10125_ vssd1 vssd1 vccd1 vccd1 _10251_ sky130_fd_sc_hd__nor2_1
X_14443_ _07306_ _07193_ _07611_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__or3b_1
X_11655_ net4132 _04701_ net4145 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10606_ net7069 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__clkbuf_1
X_17162_ _10147_ _10181_ vssd1 vssd1 vccd1 vccd1 _10182_ sky130_fd_sc_hd__xnor2_2
X_20352__108 clknet_1_0__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__inv_2
X_11586_ _04771_ _04775_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__xnor2_1
X_14374_ _07544_ _07541_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16113_ _09204_ _09206_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__xnor2_4
X_10537_ net6754 net6985 _04075_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13325_ _06343_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__inv_2
X_17093_ _10082_ _10113_ vssd1 vssd1 vccd1 vccd1 _10114_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _08542_ _08616_ vssd1 vssd1 vccd1 vccd1 _09138_ sky130_fd_sc_hd__nor2_1
X_10468_ net2852 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13256_ _06307_ _06421_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _04930_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13187_ net4513 net6015 vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__nand2_1
X_12138_ _05324_ _05325_ _04910_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__mux2_1
X_17995_ _02230_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__xor2_1
X_20547__285 clknet_1_0__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__inv_2
XFILLER_0_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12069_ _04933_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__buf_4
X_16946_ _09964_ _09967_ vssd1 vssd1 vccd1 vccd1 _09968_ sky130_fd_sc_hd__xnor2_1
X_19734_ net3921 _03496_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19665_ net6313 net4028 _03457_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16877_ _09897_ _09898_ vssd1 vssd1 vccd1 vccd1 _09899_ sky130_fd_sc_hd__nand2_1
X_18616_ _02771_ _02774_ _04489_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15828_ _08915_ _08922_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__nand2_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19596_ net6065 _03139_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18547_ _02717_ net5933 _06242_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
X_15759_ _08808_ _08813_ _08853_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18478_ _02617_ net3494 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ _10324_ _10325_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22110_ net148 net2395 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
Xhold4203 _08049_ vssd1 vssd1 vccd1 vccd1 net4730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4214 net8356 vssd1 vssd1 vccd1 vccd1 net4741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4225 _08059_ vssd1 vssd1 vccd1 vccd1 net4752 sky130_fd_sc_hd__dlygate4sd3_1
X_22041_ net483 net2532 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4247 net3535 vssd1 vssd1 vccd1 vccd1 net4774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3502 _02479_ vssd1 vssd1 vccd1 vccd1 net4029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3513 net4016 vssd1 vssd1 vccd1 vccd1 net4040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4258 _02565_ vssd1 vssd1 vccd1 vccd1 net4785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3524 _00622_ vssd1 vssd1 vccd1 vccd1 net4051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3535 net3032 vssd1 vssd1 vccd1 vccd1 net4062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2801 rbzero.pov.spi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net3328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3546 rbzero.spi_registers.spi_buffer\[3\] vssd1 vssd1 vccd1 vccd1 net4073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 net5767 vssd1 vssd1 vccd1 vccd1 net3339 sky130_fd_sc_hd__clkbuf_2
Xhold3557 _03987_ vssd1 vssd1 vccd1 vccd1 net4084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2823 rbzero.pov.spi_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net3350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3568 _04672_ vssd1 vssd1 vccd1 vccd1 net4095 sky130_fd_sc_hd__clkbuf_4
Xhold2834 rbzero.pov.ready_buffer\[36\] vssd1 vssd1 vccd1 vccd1 net3361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3579 _04683_ vssd1 vssd1 vccd1 vccd1 net4106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2845 net7767 vssd1 vssd1 vccd1 vccd1 net3372 sky130_fd_sc_hd__buf_2
Xhold2856 net4544 vssd1 vssd1 vccd1 vccd1 net3383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2867 net3694 vssd1 vssd1 vccd1 vccd1 net3394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2878 net4338 vssd1 vssd1 vccd1 vccd1 net3405 sky130_fd_sc_hd__clkbuf_2
Xhold2889 net4345 vssd1 vssd1 vccd1 vccd1 net3416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21825_ net267 net1410 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21756_ clknet_leaf_29_i_clk net5210 vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20707_ _03884_ _03885_ _03886_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21687_ clknet_leaf_115_i_clk net4494 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ _04554_ _04555_ rbzero.spi_registers.texadd3\[2\] vssd1 vssd1 vccd1 vccd1
+ _04632_ sky130_fd_sc_hd__or3b_1
X_20638_ clknet_1_0__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__buf_1
XFILLER_0_0_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ rbzero.spi_registers.texadd3\[20\] rbzero.spi_registers.texadd1\[20\] rbzero.spi_registers.texadd0\[20\]
+ rbzero.spi_registers.texadd2\[20\] _04554_ _04555_ vssd1 vssd1 vccd1 vccd1 _04563_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6150 net1767 vssd1 vssd1 vccd1 vccd1 net6677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6161 rbzero.tex_r1\[55\] vssd1 vssd1 vccd1 vccd1 net6688 sky130_fd_sc_hd__dlygate4sd3_1
X_13110_ _06279_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__nor2_2
Xhold6172 net1660 vssd1 vssd1 vccd1 vccd1 net6699 sky130_fd_sc_hd__dlygate4sd3_1
X_14090_ _07259_ _07260_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__xnor2_1
Xhold6183 rbzero.tex_g0\[21\] vssd1 vssd1 vccd1 vccd1 net6710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6194 net2430 vssd1 vssd1 vccd1 vccd1 net6721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5460 rbzero.pov.spi_buffer\[68\] vssd1 vssd1 vccd1 vccd1 net5987 sky130_fd_sc_hd__dlygate4sd3_1
X_13041_ net4657 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__inv_2
Xhold5471 net2322 vssd1 vssd1 vccd1 vccd1 net5998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5482 rbzero.spi_registers.new_floor\[2\] vssd1 vssd1 vccd1 vccd1 net6009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5493 rbzero.spi_registers.new_floor\[5\] vssd1 vssd1 vccd1 vccd1 net6020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4770 _00838_ vssd1 vssd1 vccd1 vccd1 net5297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4781 net909 vssd1 vssd1 vccd1 vccd1 net5308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4792 rbzero.spi_registers.texadd1\[15\] vssd1 vssd1 vccd1 vccd1 net5319 sky130_fd_sc_hd__dlygate4sd3_1
X_16800_ _09818_ _09089_ vssd1 vssd1 vccd1 vccd1 _09829_ sky130_fd_sc_hd__nand2_1
X_17780_ _09040_ net8008 _02018_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__or3_1
X_14992_ net63 net7571 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16731_ net4648 vssd1 vssd1 vccd1 vccd1 _09769_ sky130_fd_sc_hd__buf_4
X_13943_ _07107_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19450_ net5513 _03335_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16662_ net4080 _09737_ _09740_ _08111_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
X_13874_ _07043_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__nand2_1
X_19794__72 clknet_1_1__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
XFILLER_0_202_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18401_ net4725 net8074 _02583_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a21o_1
X_15613_ _08704_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__xnor2_4
Xclkbuf_1_0__f__05688_ clknet_0__05688_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05688_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19381_ net5173 _03283_ _03293_ _03288_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__o211a_1
X_12825_ _05949_ _05956_ _05960_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__o21ai_1
X_16593_ _09678_ _09679_ _09681_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18332_ net3661 net4883 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nand2_1
X_15544_ _08638_ _08208_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__xnor2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12756_ _05203_ _05912_ _05916_ net41 net36 vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _04458_ _02475_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__nor2_4
X_11707_ net3014 _04467_ _04896_ net4115 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__o22ai_1
X_15475_ _08496_ _08497_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and2b_1
X_17214_ _10232_ _10233_ vssd1 vssd1 vccd1 vccd1 _10234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ _07586_ _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__xor2_2
Xclkbuf_1_1__f__03852_ clknet_0__03852_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03852_
+ sky130_fd_sc_hd__clkbuf_16
X_11638_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__buf_4
XFILLER_0_142_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18194_ net3811 net4430 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17145_ _08383_ _08614_ vssd1 vssd1 vccd1 vccd1 _10165_ sky130_fd_sc_hd__nor2_1
X_14357_ _07521_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__or2_1
X_11569_ net1138 net1122 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 net5493 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 net6437 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ _06438_ _06454_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__nor2_1
X_17076_ _09537_ _10096_ vssd1 vssd1 vccd1 vccd1 _10097_ sky130_fd_sc_hd__nor2_1
Xhold729 net5502 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ _06699_ _07391_ _07458_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__nor3_2
XFILLER_0_126_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16027_ _09119_ _09120_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__or2b_2
X_13239_ _06308_ _06310_ _06367_ _06381_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2108 net7219 vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2119 _00951_ vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1407 _00686_ vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 _01026_ vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ _02200_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__xnor2_1
Xhold1429 _04351_ vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16929_ _09940_ _09950_ vssd1 vssd1 vccd1 vccd1 _09951_ sky130_fd_sc_hd__xnor2_1
X_19717_ net2309 _04102_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19648_ net6864 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__clkbuf_1
X_19579_ net2599 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21610_ clknet_leaf_132_i_clk net3103 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21541_ net175 net3007 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21472_ clknet_leaf_21_i_clk net1781 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4000 net7699 vssd1 vssd1 vccd1 vccd1 net4527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4011 net8081 vssd1 vssd1 vccd1 vccd1 net4538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4022 net3385 vssd1 vssd1 vccd1 vccd1 net4549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4033 net8245 vssd1 vssd1 vccd1 vccd1 net4560 sky130_fd_sc_hd__buf_2
X_20285_ net1341 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
Xhold4044 _08044_ vssd1 vssd1 vccd1 vccd1 net4571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3310 rbzero.spi_registers.spi_buffer\[10\] vssd1 vssd1 vccd1 vccd1 net3837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4055 net8415 vssd1 vssd1 vccd1 vccd1 net4582 sky130_fd_sc_hd__dlygate4sd3_1
X_22024_ net466 net1850 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
Xhold4066 net1172 vssd1 vssd1 vccd1 vccd1 net4593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3321 net5932 vssd1 vssd1 vccd1 vccd1 net3848 sky130_fd_sc_hd__buf_2
Xhold4077 _03763_ vssd1 vssd1 vccd1 vccd1 net4604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3332 _09723_ vssd1 vssd1 vccd1 vccd1 net3859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3343 net5921 vssd1 vssd1 vccd1 vccd1 net3870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4088 net3365 vssd1 vssd1 vccd1 vccd1 net4615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4099 _03712_ vssd1 vssd1 vccd1 vccd1 net4626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3354 net7623 vssd1 vssd1 vccd1 vccd1 net3881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2620 _01096_ vssd1 vssd1 vccd1 vccd1 net3147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3365 net5893 vssd1 vssd1 vccd1 vccd1 net3892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 rbzero.pov.spi_buffer\[63\] vssd1 vssd1 vccd1 vccd1 net3158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3376 net5941 vssd1 vssd1 vccd1 vccd1 net3903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2642 net7372 vssd1 vssd1 vccd1 vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2653 net7545 vssd1 vssd1 vccd1 vccd1 net3180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03872_ clknet_0__03872_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03872_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3398 net7997 vssd1 vssd1 vccd1 vccd1 net3925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2664 net3236 vssd1 vssd1 vccd1 vccd1 net3191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1930 _04425_ vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 net7499 vssd1 vssd1 vccd1 vccd1 net3202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net4929 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1941 net7537 vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2686 rbzero.pov.spi_buffer\[40\] vssd1 vssd1 vccd1 vccd1 net3213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 net4941 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1952 net7296 vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2697 _03055_ vssd1 vssd1 vccd1 vccd1 net3224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1963 _01069_ vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold89 net6686 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1974 _01577_ vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1985 net7241 vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ net6725 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
Xhold1996 _01426_ vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ net7216 net6593 _04253_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ _05783_ _05785_ _05786_ _05745_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a221o_2
X_21808_ net250 net2559 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13590_ _06756_ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _04021_ _05701_ _05699_ _04495_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a22o_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21739_ clknet_leaf_99_i_clk net3497 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _08168_ _08211_ _08221_ _08241_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12472_ _04648_ _04461_ _04468_ _04023_ _05633_ net5 vssd1 vssd1 vccd1 vccd1 _05654_
+ sky130_fd_sc_hd__mux4_1
X_14211_ _07380_ _07381_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11423_ _04539_ _04517_ _04537_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nand3_1
X_15191_ _08132_ _08143_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _05795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14142_ _07240_ _07233_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nor2_1
X_11354_ rbzero.spi_registers.texadd2\[13\] _04544_ _04545_ rbzero.spi_registers.texadd0\[13\]
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14073_ _07200_ _07230_ _07228_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_46_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11285_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__clkbuf_4
X_18950_ net3138 net5704 _03036_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
Xhold5290 _03616_ vssd1 vssd1 vccd1 vccd1 net5817 sky130_fd_sc_hd__dlygate4sd3_1
X_17901_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__and2_1
X_13024_ net3803 _06198_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__o21ba_1
X_20464__209 clknet_1_0__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__inv_2
X_18881_ net2771 net4803 _03003_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17832_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _09272_ _01693_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14975_ _08085_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19502_ net1644 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
X_16714_ net4007 _09102_ vssd1 vssd1 vccd1 vccd1 _09752_ sky130_fd_sc_hd__xnor2_2
X_13926_ _06911_ _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__xnor2_2
X_17694_ _01932_ _01933_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19433_ net1593 net3519 _03141_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ net4108 net4124 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__nor2_1
X_13857_ _06952_ _06990_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__xor2_2
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20659__386 clknet_1_1__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__inv_2
X_12808_ net7746 net5955 vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__and2_1
X_19364_ _03270_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__clkbuf_4
X_16576_ _09548_ _09417_ _06123_ vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__a21o_2
XFILLER_0_128_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20358__114 clknet_1_1__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__inv_2
X_13788_ _06703_ _06698_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__nor2_1
X_18315_ net6160 net3583 _02476_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15527_ _08609_ _08610_ _08620_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__and3_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12739_ _05904_ net34 vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nor2_1
X_19295_ net6390 _03238_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7609 _00821_ vssd1 vssd1 vccd1 vccd1 net8136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18246_ _02459_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15458_ _08551_ _08552_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6908 net3090 vssd1 vssd1 vccd1 vccd1 net7435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6919 rbzero.tex_b0\[44\] vssd1 vssd1 vccd1 vccd1 net7446 sky130_fd_sc_hd__dlygate4sd3_1
X_14409_ _07568_ _07577_ _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__a21oi_2
X_18177_ _02400_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__clkbuf_1
X_15389_ _08467_ _08471_ _08478_ _08483_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17128_ _10081_ _10059_ vssd1 vssd1 vccd1 vccd1 _10148_ sky130_fd_sc_hd__or2b_1
Xhold504 _03423_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03866_ _03866_ vssd1 vssd1 vccd1 vccd1 clknet_0__03866_ sky130_fd_sc_hd__clkbuf_16
Xhold515 _01583_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold526 net6157 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold537 net6143 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold548 net7897 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkdlybuf4s25_1
X_17059_ _10060_ _10061_ _10078_ vssd1 vssd1 vccd1 vccd1 _10080_ sky130_fd_sc_hd__nand3_1
Xhold559 net7894 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20070_ net5750 _03485_ _03662_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a211o_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 net6674 vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 net6543 vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _03012_ vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1237 net5569 vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _01054_ vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 _03827_ vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20972_ clknet_leaf_111_i_clk net4151 vssd1 vssd1 vccd1 vccd1 reg_rgb\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19773__53 clknet_1_0__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21524_ clknet_leaf_3_i_clk net2416 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21455_ clknet_leaf_26_i_clk net3981 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vshift
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21386_ clknet_leaf_3_i_clk net5191 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__buf_1
X_11070_ net5594 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__clkbuf_4
X_20268_ net4128 net4097 net4178 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3140 _02397_ vssd1 vssd1 vccd1 vccd1 net3667 sky130_fd_sc_hd__dlygate4sd3_1
X_22007_ net449 net2093 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold3151 _02792_ vssd1 vssd1 vccd1 vccd1 net3678 sky130_fd_sc_hd__clkbuf_4
Xhold3162 _01208_ vssd1 vssd1 vccd1 vccd1 net3689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3173 _02316_ vssd1 vssd1 vccd1 vccd1 net3700 sky130_fd_sc_hd__buf_1
X_20199_ net4698 _03744_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__or2_1
Xhold3184 net7582 vssd1 vssd1 vccd1 vccd1 net3711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2450 rbzero.tex_b1\[13\] vssd1 vssd1 vccd1 vccd1 net2977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3195 _01205_ vssd1 vssd1 vccd1 vccd1 net3722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2461 _04399_ vssd1 vssd1 vccd1 vccd1 net2988 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2472 net7426 vssd1 vssd1 vccd1 vccd1 net2999 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 _03591_ vssd1 vssd1 vccd1 vccd1 net3010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03855_ clknet_0__03855_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03855_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2494 _00655_ vssd1 vssd1 vccd1 vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 _01337_ vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1771 _04038_ vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ net7787 _07864_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__or2_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ rbzero.debug_overlay.vplaneY\[-9\] _05106_ _05114_ net3575 _05160_ vssd1
+ vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a221o_1
Xhold1782 net7505 vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1793 _01476_ vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _06872_ _06880_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__o21ai_2
X_10923_ net2732 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _07695_ _07774_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16430_ _09519_ _09520_ vssd1 vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__nand2_1
X_13642_ net79 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ net3104 net5700 _04238_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _09450_ net8520 vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ _06634_ _06732_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__or2_4
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ net7210 net7399 _04205_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18100_ _06058_ _02332_ _09810_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__o21ai_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _04511_ net8500 _08114_ _08406_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__o211a_1
X_19080_ net4062 net7277 _09725_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
X_12524_ net12 _05704_ net13 vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__o21a_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _08389_ _09262_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20677__22 clknet_1_0__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
X_18031_ _02173_ _02178_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nor2_1
X_15243_ _08131_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12455_ net4149 net4141 net4164 net7727 _05633_ net7 vssd1 vssd1 vccd1 vccd1 _05637_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ _04496_ _04596_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a21o_1
X_15174_ _08213_ _08268_ vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12386_ _04922_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or2_1
X_14125_ _07257_ _07295_ _07262_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ rbzero.texu_hot\[2\] _04520_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or2_1
X_19982_ net2890 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
X_14056_ _07183_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__xor2_1
X_18933_ net6731 net3435 _03025_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
X_11268_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _06178_ _06180_ _06181_ _06182_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__or4_1
X_11199_ net6096 net1897 _04423_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
X_18864_ net6413 net6560 _02993_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17815_ _02053_ net4723 _10260_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
X_18795_ _02866_ net5955 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_206_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17746_ _01982_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14958_ _08076_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ _07076_ _07078_ _07074_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17677_ _01892_ _01916_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__xnor2_1
X_14889_ _04481_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ _04684_ _04648_ _05057_ vssd1 vssd1 vccd1 vccd1 _09717_ sky130_fd_sc_hd__and3_1
X_19416_ net3571 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16559_ _09639_ _09648_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__xnor2_1
X_19347_ _03205_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7406 _00499_ vssd1 vssd1 vccd1 vccd1 net7933 sky130_fd_sc_hd__dlygate4sd3_1
X_19278_ net1523 _03202_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7428 rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 net7955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7439 net3789 vssd1 vssd1 vccd1 vccd1 net7966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6705 net2722 vssd1 vssd1 vccd1 vccd1 net7232 sky130_fd_sc_hd__dlygate4sd3_1
X_18229_ _02444_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__nor2_1
Xhold6716 rbzero.tex_b0\[49\] vssd1 vssd1 vccd1 vccd1 net7243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6727 net2670 vssd1 vssd1 vccd1 vccd1 net7254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6738 rbzero.tex_r1\[8\] vssd1 vssd1 vccd1 vccd1 net7265 sky130_fd_sc_hd__dlygate4sd3_1
X_21240_ clknet_leaf_44_i_clk net3865 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6749 rbzero.spi_registers.ss_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net7276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold301 net5180 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 net6425 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 net8078 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold334 net5265 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03849_ _03849_ vssd1 vssd1 vccd1 vccd1 clknet_0__03849_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21171_ clknet_leaf_132_i_clk net2945 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_20412__163 clknet_1_1__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__inv_2
XFILLER_0_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold345 net5399 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold356 net5190 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 net5407 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 net6097 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20122_ _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold389 net5341 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20053_ net4019 _03651_ _03656_ _03606_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _01333_ vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _02489_ vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 net5517 vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1034 net6020 vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1045 _00985_ vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 _03390_ vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 _03356_ vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1078 net6580 vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 net5580 vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ clknet_leaf_81_i_clk _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ net4940 net6100 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ net2336 net6607 _04086_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7940 net4907 vssd1 vssd1 vccd1 vccd1 net8467 sky130_fd_sc_hd__clkbuf_2
X_21507_ clknet_leaf_45_i_clk net1348 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7973 _05995_ vssd1 vssd1 vccd1 vccd1 net8500 sky130_fd_sc_hd__dlygate4sd3_1
X_12240_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _04968_ vssd1 vssd1 vccd1 vccd1 _05427_
+ sky130_fd_sc_hd__mux2_1
X_21438_ clknet_leaf_25_i_clk net1642 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12171_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _04916_ vssd1 vssd1 vccd1 vccd1 _05359_
+ sky130_fd_sc_hd__mux2_1
X_21369_ clknet_leaf_14_i_clk net5043 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11122_ net5686 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
X_20387__140 clknet_1_1__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__inv_2
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold890 net6420 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ net6221 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
X_15930_ _08427_ _08428_ _08429_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__a21oi_4
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _08946_ _08950_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__or2_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _01839_ _01840_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__nand2_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2280 net3076 vssd1 vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
Xhold2291 _04125_ vssd1 vssd1 vccd1 vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _07926_ _07944_ _07959_ _07972_ net7787 net7785 vssd1 vssd1 vccd1 vccd1 _07973_
+ sky130_fd_sc_hd__mux4_2
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ net4000 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15792_ _08860_ _08884_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__xnor2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1590 net6875 vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
X_17531_ _10407_ _10418_ _10416_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a21oi_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_103 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_103/HI o_rgb[12]
+ sky130_fd_sc_hd__conb_1
X_14743_ net8354 _07910_ net7833 vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__o21a_1
Xtop_ew_algofoogle_114 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_114/HI zeros[3] sky130_fd_sc_hd__conb_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ rbzero.debug_overlay.facingY\[-5\] _05108_ _04657_ net4126 net4160 vssd1
+ vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a2111o_1
Xtop_ew_algofoogle_125 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_125/HI zeros[14]
+ sky130_fd_sc_hd__conb_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_136 vssd1 vssd1 vccd1 vccd1 ones[9] top_ew_algofoogle_136/LO sky130_fd_sc_hd__conb_1
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ net6166 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
X_17462_ _01700_ _01702_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14674_ _07818_ _07837_ net8491 vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__o21ai_1
X_11886_ _05066_ _05067_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and2b_1
X_16413_ _09374_ _09503_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19201_ _09721_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__buf_4
X_19752__34 clknet_1_0__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ _06724_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__xnor2_4
X_10837_ net7043 net7005 _04227_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__mux2_1
X_17393_ _10409_ _10410_ vssd1 vssd1 vccd1 vccd1 _10411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19132_ net4354 _03145_ net1290 _03149_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__o211a_1
X_16344_ _09390_ _09435_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ _06666_ _06668_ _06671_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__nand3_4
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10768_ net7091 net7137 _04194_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12507_ reg_gpout\[0\] clknet_1_1__leaf__05688_ _05054_ vssd1 vssd1 vccd1 vccd1 _05689_
+ sky130_fd_sc_hd__mux2_2
X_19063_ net7603 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16275_ _09365_ _09366_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13487_ _06656_ _06657_ _06606_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a21o_1
X_10699_ net1927 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__clkbuf_1
X_18014_ net4622 _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__nor2_1
X_15226_ _08162_ _08194_ _08295_ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__or3_1
X_12438_ _05617_ _05620_ _05622_ _05018_ _05203_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15157_ _08118_ _08250_ _08251_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__a21o_2
X_12369_ _04922_ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14108_ _07244_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__xnor2_4
Xhold3909 net8235 vssd1 vssd1 vccd1 vccd1 net4436 sky130_fd_sc_hd__clkbuf_4
X_19965_ net3237 net5764 net2312 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__mux2_1
X_15088_ _07957_ net8378 _08113_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ _07122_ _07170_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18916_ _02992_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__clkbuf_4
X_19896_ net3125 net6731 _03550_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__mux2_1
X_19815__90 clknet_1_1__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__inv_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18847_ net5799 _02983_ _02969_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_207_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18778_ _02866_ net4709 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20442__189 clknet_1_1__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__inv_2
XFILLER_0_171_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17729_ _01966_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20740_ _03915_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20671_ clknet_1_0__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__buf_1
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7203 net3656 vssd1 vssd1 vccd1 vccd1 net7730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7214 _03724_ vssd1 vssd1 vccd1 vccd1 net7741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7225 net8317 vssd1 vssd1 vccd1 vccd1 net7752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7236 net8361 vssd1 vssd1 vccd1 vccd1 net7763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6502 net2417 vssd1 vssd1 vccd1 vccd1 net7029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6513 _04345_ vssd1 vssd1 vccd1 vccd1 net7040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7258 _07912_ vssd1 vssd1 vccd1 vccd1 net7785 sky130_fd_sc_hd__buf_2
Xhold6524 net1964 vssd1 vssd1 vccd1 vccd1 net7051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7269 rbzero.wall_tracer.stepDistY\[10\] vssd1 vssd1 vccd1 vccd1 net7796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6535 rbzero.tex_r1\[41\] vssd1 vssd1 vccd1 vccd1 net7062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6546 net2218 vssd1 vssd1 vccd1 vccd1 net7073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5801 _03596_ vssd1 vssd1 vccd1 vccd1 net6328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5812 net1380 vssd1 vssd1 vccd1 vccd1 net6339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6557 rbzero.spi_registers.new_mapd\[8\] vssd1 vssd1 vccd1 vccd1 net7084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6568 net2187 vssd1 vssd1 vccd1 vccd1 net7095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5823 rbzero.spi_registers.new_texadd\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net6350
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6579 rbzero.tex_b0\[28\] vssd1 vssd1 vccd1 vccd1 net7106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5834 net1795 vssd1 vssd1 vccd1 vccd1 net6361 sky130_fd_sc_hd__dlygate4sd3_1
X_21223_ clknet_leaf_24_i_clk net1473 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 net7862 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5845 net1355 vssd1 vssd1 vccd1 vccd1 net6372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 net4983 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5856 rbzero.spi_registers.new_texadd\[2\]\[16\] vssd1 vssd1 vccd1 vccd1 net6383
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net4993 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5867 rbzero.spi_registers.new_mapd\[2\] vssd1 vssd1 vccd1 vccd1 net6394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _01658_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5878 net1508 vssd1 vssd1 vccd1 vccd1 net6405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 net5048 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
X_21154_ clknet_leaf_23_i_clk net3912 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5889 rbzero.spi_registers.new_texadd\[1\]\[10\] vssd1 vssd1 vccd1 vccd1 net6416
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 net5078 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 net5052 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 net5094 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20105_ net3473 _03690_ _03484_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21085_ clknet_leaf_46_i_clk net1288 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20036_ net3990 _03634_ net3389 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__o21ai_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21987_ net429 net2594 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04832_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__buf_4
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ clknet_leaf_77_i_clk net4697 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_131_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ net3365 _04859_ net3423 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_193_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20869_ _02510_ _02516_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__or2b_1
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13410_ _06472_ _06558_ _06580_ _06550_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__a211o_1
X_10622_ net5577 net2581 _04116_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14390_ _06771_ _07232_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20419__169 clknet_1_1__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__inv_2
XFILLER_0_14_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13341_ _06500_ _06507_ _06474_ _06498_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__and4b_1
XFILLER_0_162_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10553_ net2342 net5659 _04075_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16060_ _09019_ _09021_ _09018_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__a21bo_1
Xhold7770 net4193 vssd1 vssd1 vccd1 vccd1 net8297 sky130_fd_sc_hd__dlygate4sd3_1
X_13272_ _06335_ _06337_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and2_1
Xhold7781 net1361 vssd1 vssd1 vccd1 vccd1 net8308 sky130_fd_sc_hd__dlygate4sd3_1
X_10484_ net7268 net7359 _04042_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__mux2_1
Xhold7792 net4406 vssd1 vssd1 vccd1 vccd1 net8319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ net1004 net4010 net3985 vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__mux2_1
X_12223_ rbzero.tex_g1\[27\] rbzero.tex_g1\[26\] _04837_ vssd1 vssd1 vccd1 vccd1 _05410_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12154_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _04916_ vssd1 vssd1 vccd1 vccd1 _05342_
+ sky130_fd_sc_hd__mux2_1
X_11105_ net2601 net7075 _04375_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
X_12085_ rbzero.tex_r1\[61\] rbzero.tex_r1\[60\] _05220_ vssd1 vssd1 vccd1 vccd1 _05274_
+ sky130_fd_sc_hd__mux2_1
X_16962_ _09981_ _09982_ _09983_ vssd1 vssd1 vccd1 vccd1 _09984_ sky130_fd_sc_hd__nand3_1
XFILLER_0_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18701_ _04490_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__nand2_1
X_11036_ net6444 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
X_15913_ _09006_ _09007_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16893_ _08383_ vssd1 vssd1 vccd1 vccd1 _09915_ sky130_fd_sc_hd__clkbuf_4
X_19681_ net6351 net2953 _03457_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15844_ _08902_ _08911_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__xnor2_1
X_18632_ net4528 _02780_ _04480_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a21oi_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15775_ _08161_ _08280_ _08318_ _08402_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18563_ net7577 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _06162_ net4742 vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__and2_2
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17514_ _01752_ _01753_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__and2_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07841_ _07819_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__o21ai_1
X_18494_ _02666_ _02667_ net4868 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a21o_1
X_11938_ net3445 _05080_ _05093_ net3326 _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17445_ _01685_ _01686_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _07814_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__inv_2
X_11869_ _04461_ _04026_ _04601_ _05057_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and4_1
XFILLER_0_185_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ _06765_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ _10335_ _10313_ vssd1 vssd1 vccd1 vccd1 _10394_ sky130_fd_sc_hd__or2b_1
XFILLER_0_172_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14588_ _07751_ _07757_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16327_ net4537 _08491_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19115_ net1076 _03126_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or2_1
X_13539_ _06706_ _06695_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20630__359 clknet_1_1__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__inv_2
X_19046_ net3738 net7621 net3398 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
X_16258_ _09231_ _09234_ _09232_ vssd1 vssd1 vccd1 vccd1 _09350_ sky130_fd_sc_hd__a21bo_1
Xhold5108 _04352_ vssd1 vssd1 vccd1 vccd1 net5635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5119 _04066_ vssd1 vssd1 vccd1 vccd1 net5646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15209_ _08133_ _08302_ _08303_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4407 net596 vssd1 vssd1 vccd1 vccd1 net4934 sky130_fd_sc_hd__dlygate4sd3_1
X_16189_ _09274_ _09281_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__xnor2_1
Xhold4418 _01021_ vssd1 vssd1 vccd1 vccd1 net4945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4429 net612 vssd1 vssd1 vccd1 vccd1 net4956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3706 rbzero.wall_tracer.visualWallDist\[6\] vssd1 vssd1 vccd1 vccd1 net4233 sky130_fd_sc_hd__buf_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3717 net7914 vssd1 vssd1 vccd1 vccd1 net4244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3728 net1010 vssd1 vssd1 vccd1 vccd1 net4255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3739 _00519_ vssd1 vssd1 vccd1 vccd1 net4266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19948_ net6241 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19879_ net7556 net3342 _03539_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__mux2_1
X_21910_ net352 net2888 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
X_20524__264 clknet_1_0__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__inv_2
XFILLER_0_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21841_ net283 net2065 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21772_ clknet_leaf_45_i_clk net1467 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20723_ _03899_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7000 rbzero.pov.spi_buffer\[3\] vssd1 vssd1 vccd1 vccd1 net7527 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_63_i_clk clknet_4_14__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold7011 net2468 vssd1 vssd1 vccd1 vccd1 net7538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7022 rbzero.pov.ready_buffer\[31\] vssd1 vssd1 vccd1 vccd1 net7549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7033 net2829 vssd1 vssd1 vccd1 vccd1 net7560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7044 net4068 vssd1 vssd1 vccd1 vccd1 net7571 sky130_fd_sc_hd__clkbuf_4
Xhold6310 _04039_ vssd1 vssd1 vccd1 vccd1 net6837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7055 rbzero.pov.ready_buffer\[29\] vssd1 vssd1 vccd1 vccd1 net7582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6321 net2108 vssd1 vssd1 vccd1 vccd1 net6848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7066 net1113 vssd1 vssd1 vccd1 vccd1 net7593 sky130_fd_sc_hd__buf_1
Xhold6332 rbzero.tex_r0\[28\] vssd1 vssd1 vccd1 vccd1 net6859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7077 rbzero.pov.ready_buffer\[72\] vssd1 vssd1 vccd1 vccd1 net7604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6343 net1910 vssd1 vssd1 vccd1 vccd1 net6870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7088 net3674 vssd1 vssd1 vccd1 vccd1 net7615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6354 _04051_ vssd1 vssd1 vccd1 vccd1 net6881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7099 _03733_ vssd1 vssd1 vccd1 vccd1 net7626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6365 net2579 vssd1 vssd1 vccd1 vccd1 net6892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5620 rbzero.spi_registers.new_texadd\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net6147
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5631 net1053 vssd1 vssd1 vccd1 vccd1 net6158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6376 rbzero.tex_b0\[63\] vssd1 vssd1 vccd1 vccd1 net6903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6387 net2423 vssd1 vssd1 vccd1 vccd1 net6914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5642 _04217_ vssd1 vssd1 vccd1 vccd1 net6169 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_78_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold6398 _04268_ vssd1 vssd1 vccd1 vccd1 net6925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5653 net1219 vssd1 vssd1 vccd1 vccd1 net6180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5664 net1343 vssd1 vssd1 vccd1 vccd1 net6191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5675 rbzero.tex_g1\[48\] vssd1 vssd1 vccd1 vccd1 net6202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21206_ clknet_leaf_117_i_clk net3254 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4930 _00845_ vssd1 vssd1 vccd1 vccd1 net5457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5686 net1174 vssd1 vssd1 vccd1 vccd1 net6213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4941 net1163 vssd1 vssd1 vccd1 vccd1 net5468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4952 rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 net5479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5697 _04242_ vssd1 vssd1 vccd1 vccd1 net6224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4963 net1218 vssd1 vssd1 vccd1 vccd1 net5490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4974 _03307_ vssd1 vssd1 vccd1 vccd1 net5501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4985 rbzero.spi_registers.new_vshift\[1\] vssd1 vssd1 vccd1 vccd1 net5512 sky130_fd_sc_hd__dlygate4sd3_1
X_21137_ clknet_leaf_95_i_clk net4533 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4996 net8230 vssd1 vssd1 vccd1 vccd1 net5523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21068_ clknet_leaf_59_i_clk _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20019_ _03608_ net4491 vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or2_1
X_12910_ net3443 net3960 net3884 _06084_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__o22a_1
X_13890_ _07058_ _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nor2_1
X_20499__241 clknet_1_0__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__inv_2
X_12841_ _05978_ _05977_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__or2b_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _08624_ _08654_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__xnor2_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12772_ net4416 net3761 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__nand2_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _07673_ _07674_ _07680_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__and3_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__clkbuf_8
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _08568_ _08569_ _08585_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__a21o_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _10021_ _10249_ vssd1 vssd1 vccd1 vccd1 _10250_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _07284_ _07326_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ _04814_ _04816_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nor2_4
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10605_ net7067 net2384 _04105_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__mux2_1
X_17161_ _10179_ _10180_ vssd1 vssd1 vccd1 vccd1 _10181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14373_ _07492_ _07538_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__nand2_2
X_11585_ net2494 _04774_ _04772_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _08621_ _09075_ _09205_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_181_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ _06351_ _06434_ _06442_ _06454_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__or4_4
XFILLER_0_107_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17092_ _10111_ _10112_ vssd1 vssd1 vccd1 vccd1 _10113_ sky130_fd_sc_hd__xor2_2
X_10536_ net2466 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _09134_ _09136_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _06414_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__nand2_1
X_10467_ net6689 net7236 _04031_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ rbzero.tex_g1\[7\] rbzero.tex_g1\[6\] _04923_ vssd1 vssd1 vccd1 vccd1 _05393_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ net8269 _06265_ _06306_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__o21a_1
XFILLER_0_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _04950_ vssd1 vssd1 vccd1 vccd1 _05325_
+ sky130_fd_sc_hd__mux2_1
X_17994_ _02064_ _02140_ _02138_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19733_ net7648 _03496_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__and2_1
X_12068_ _05255_ _05256_ _04984_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__mux2_1
X_16945_ _09965_ _09966_ vssd1 vssd1 vccd1 vccd1 _09967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_205_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11019_ net2063 net6249 _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19664_ net1308 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
X_16876_ _09603_ _09896_ vssd1 vssd1 vccd1 vccd1 _09898_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18615_ _02771_ _02774_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15827_ _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__nor2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ net6576 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15758_ _08826_ _08851_ _08852_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18546_ net4436 _09818_ _02715_ _02716_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a22o_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14709_ net7843 _07877_ _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__or3_4
X_15689_ _08241_ _08328_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__nor2_1
X_18477_ _02640_ _02646_ _02653_ _04489_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _01668_ _01669_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17359_ _10266_ _10268_ _10377_ vssd1 vssd1 vccd1 vccd1 _10378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19029_ net3863 net3816 _03078_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4204 _00421_ vssd1 vssd1 vccd1 vccd1 net4731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4215 net3933 vssd1 vssd1 vccd1 vccd1 net4742 sky130_fd_sc_hd__clkbuf_2
X_22040_ net482 net2160 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold4226 _00429_ vssd1 vssd1 vccd1 vccd1 net4753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4237 _02820_ vssd1 vssd1 vccd1 vccd1 net4764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3503 net1396 vssd1 vssd1 vccd1 vccd1 net4030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4248 net8446 vssd1 vssd1 vccd1 vccd1 net4775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3514 _03084_ vssd1 vssd1 vccd1 vccd1 net4041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4259 net8050 vssd1 vssd1 vccd1 vccd1 net4786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3525 net4747 vssd1 vssd1 vccd1 vccd1 net4052 sky130_fd_sc_hd__clkbuf_2
Xhold3536 _02969_ vssd1 vssd1 vccd1 vccd1 net4063 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2802 net3210 vssd1 vssd1 vccd1 vccd1 net3329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3547 net1425 vssd1 vssd1 vccd1 vccd1 net4074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2813 net4444 vssd1 vssd1 vccd1 vccd1 net3340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3558 _03990_ vssd1 vssd1 vccd1 vccd1 net4085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 net3230 vssd1 vssd1 vccd1 vccd1 net3351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3569 _03118_ vssd1 vssd1 vccd1 vccd1 net4096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2835 net1026 vssd1 vssd1 vccd1 vccd1 net3362 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2846 net5752 vssd1 vssd1 vccd1 vccd1 net3373 sky130_fd_sc_hd__dlygate4sd3_1
X_20448__195 clknet_1_0__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__inv_2
Xhold2857 net7972 vssd1 vssd1 vccd1 vccd1 net3384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2868 _03075_ vssd1 vssd1 vccd1 vccd1 net3395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2879 net7906 vssd1 vssd1 vccd1 vccd1 net3406 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21824_ net266 net1957 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21755_ clknet_leaf_83_i_clk net5986 vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20706_ net5384 _03877_ _03874_ _03888_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a22o_1
X_21686_ clknet_leaf_115_i_clk net5853 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ rbzero.spi_registers.texadd3\[19\] rbzero.spi_registers.texadd1\[19\] rbzero.spi_registers.texadd0\[19\]
+ rbzero.spi_registers.texadd2\[19\] _04554_ _04555_ vssd1 vssd1 vccd1 vccd1 _04562_
+ sky130_fd_sc_hd__mux4_2
Xhold6140 net1870 vssd1 vssd1 vccd1 vccd1 net6667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6151 _03833_ vssd1 vssd1 vccd1 vccd1 net6678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6162 net2119 vssd1 vssd1 vccd1 vccd1 net6689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6173 _04362_ vssd1 vssd1 vccd1 vccd1 net6700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6184 net2110 vssd1 vssd1 vccd1 vccd1 net6711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5450 rbzero.spi_registers.got_new_leak vssd1 vssd1 vccd1 vccd1 net5977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6195 rbzero.tex_g0\[26\] vssd1 vssd1 vccd1 vccd1 net6722 sky130_fd_sc_hd__dlygate4sd3_1
X_13040_ _06205_ net3888 _06214_ _06215_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__a211o_1
Xhold5461 net587 vssd1 vssd1 vccd1 vccd1 net5988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5472 gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 net5999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5483 net1564 vssd1 vssd1 vccd1 vccd1 net6010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5494 net1561 vssd1 vssd1 vccd1 vccd1 net6021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4760 rbzero.spi_registers.texadd3\[9\] vssd1 vssd1 vccd1 vccd1 net5287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4771 net903 vssd1 vssd1 vccd1 vccd1 net5298 sky130_fd_sc_hd__dlygate4sd3_1
X_22169_ clknet_leaf_91_i_clk net1097 vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4782 _00825_ vssd1 vssd1 vccd1 vccd1 net5309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4793 net944 vssd1 vssd1 vccd1 vccd1 net5320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14991_ net4157 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
X_13942_ _07111_ _07112_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__xor2_1
X_16730_ _06058_ net4648 vssd1 vssd1 vccd1 vccd1 _09768_ sky130_fd_sc_hd__nor2_2
X_16661_ _09739_ vssd1 vssd1 vccd1 vccd1 _09740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13873_ _06715_ _06754_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15612_ _08705_ _08706_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__nor2_2
X_18400_ _02574_ _02575_ _02576_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a21bo_1
X_12824_ _05949_ _05956_ _05960_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__or3_4
X_16592_ _09678_ _09679_ _09681_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__nand3_1
X_19380_ net6677 _03284_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15543_ _08212_ _08187_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18331_ net3660 net4883 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__nor2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _04020_ _04495_ _04494_ _04500_ _05901_ net35 vssd1 vssd1 vccd1 vccd1 _05932_
+ sky130_fd_sc_hd__mux4_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ net1880 net4815 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__nand2_2
X_11706_ net3365 net3014 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__xnor2_1
X_15474_ _08505_ _08499_ _08504_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ net28 net29 vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17213_ _10094_ _10110_ _10108_ vssd1 vssd1 vccd1 vccd1 _10233_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_155_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14425_ _07588_ _07594_ _07595_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__a21oi_2
X_11637_ _04800_ _04814_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__or3_1
X_18193_ net3811 net4430 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__03851_ clknet_0__03851_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03851_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17144_ _10062_ _10163_ _09935_ vssd1 vssd1 vccd1 vccd1 _10164_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14356_ _07522_ _07525_ _07526_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__a21boi_4
X_11568_ net1138 net1122 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold708 net6258 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13307_ _06386_ _06388_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ net5639 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__clkbuf_1
X_17075_ _10095_ vssd1 vssd1 vccd1 vccd1 _10096_ sky130_fd_sc_hd__buf_4
Xhold719 _00680_ vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14287_ _06696_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11499_ net3682 _04022_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16026_ _08995_ _08999_ _09118_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ _06264_ _06408_ _06307_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_204_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13169_ _06339_ _06271_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__xnor2_1
Xhold2109 _04152_ vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1408 net6811 vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
X_17977_ _02212_ _02213_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__xor2_1
Xhold1419 net3185 vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19716_ net7272 net3220 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__nor2b_1
X_16928_ _09948_ _09949_ vssd1 vssd1 vccd1 vccd1 _09950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19647_ net6862 net3674 _03441_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16859_ _09881_ net4581 net4649 vssd1 vssd1 vccd1 vccd1 _09882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19578_ net7475 net3816 _03403_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18529_ _02627_ net5952 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21540_ net174 net2317 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
X_20636__365 clknet_1_0__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__inv_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ clknet_leaf_21_i_clk net1657 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4001 net3538 vssd1 vssd1 vccd1 vccd1 net4528 sky130_fd_sc_hd__buf_4
XFILLER_0_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4012 net3728 vssd1 vssd1 vccd1 vccd1 net4539 sky130_fd_sc_hd__clkbuf_2
Xhold4023 net4239 vssd1 vssd1 vccd1 vccd1 net4550 sky130_fd_sc_hd__clkbuf_2
X_20284_ net6275 net3897 _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__mux2_1
Xhold4034 _03778_ vssd1 vssd1 vccd1 vccd1 net4561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4045 _00417_ vssd1 vssd1 vccd1 vccd1 net4572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3311 net1477 vssd1 vssd1 vccd1 vccd1 net3838 sky130_fd_sc_hd__buf_2
X_22023_ net465 net2425 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4056 net3788 vssd1 vssd1 vccd1 vccd1 net4583 sky130_fd_sc_hd__clkbuf_2
Xhold3322 net5934 vssd1 vssd1 vccd1 vccd1 net3849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4078 _01228_ vssd1 vssd1 vccd1 vccd1 net4605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3333 _00473_ vssd1 vssd1 vccd1 vccd1 net3860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4089 net5703 vssd1 vssd1 vccd1 vccd1 net4616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3344 _04473_ vssd1 vssd1 vccd1 vccd1 net3871 sky130_fd_sc_hd__buf_2
Xhold2610 rbzero.pov.spi_buffer\[45\] vssd1 vssd1 vccd1 vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3355 _03738_ vssd1 vssd1 vccd1 vccd1 net3882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 net3194 vssd1 vssd1 vccd1 vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3366 net5973 vssd1 vssd1 vccd1 vccd1 net3893 sky130_fd_sc_hd__buf_2
Xhold2632 net1471 vssd1 vssd1 vccd1 vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3377 _00910_ vssd1 vssd1 vccd1 vccd1 net3904 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2643 _04215_ vssd1 vssd1 vccd1 vccd1 net3170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3388 _02834_ vssd1 vssd1 vccd1 vccd1 net3915 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03871_ clknet_0__03871_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03871_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2654 _00675_ vssd1 vssd1 vccd1 vccd1 net3181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3399 net3476 vssd1 vssd1 vccd1 vccd1 net3926 sky130_fd_sc_hd__clkbuf_2
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1920 net6937 vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2665 net5792 vssd1 vssd1 vccd1 vccd1 net3192 sky130_fd_sc_hd__dlygate4sd3_1
X_20381__135 clknet_1_0__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__inv_2
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1931 _01052_ vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2676 _04267_ vssd1 vssd1 vccd1 vccd1 net3203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 net5787 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1942 _03001_ vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 net4931 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net4951 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2687 net2584 vssd1 vssd1 vccd1 vccd1 net3214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 _04435_ vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 _00703_ vssd1 vssd1 vccd1 vccd1 net3225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1964 net7193 vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1975 rbzero.tex_g0\[63\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1986 _04397_ vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1997 net7265 vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _04104_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21807_ net249 net2369 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _05705_ _05710_ _05715_ _05720_ net15 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__o32a_2
XFILLER_0_186_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21738_ clknet_leaf_98_i_clk net4701 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ _05641_ _05648_ _05650_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a22o_2
XFILLER_0_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21669_ clknet_leaf_123_i_clk net3239 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
X_14210_ _07370_ _07379_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ _04537_ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and2_1
X_15190_ _08213_ _08268_ _08284_ vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__a21bo_2
X_14141_ _07284_ _07305_ _07310_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__o31a_1
XFILLER_0_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11353_ _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14072_ _07191_ _07231_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nor2_4
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11284_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13023_ _06194_ net4575 net3803 _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__a22o_1
X_17900_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__nor2_1
Xhold5291 _03617_ vssd1 vssd1 vccd1 vccd1 net5818 sky130_fd_sc_hd__dlygate4sd3_1
X_18880_ net7411 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
Xhold4590 net760 vssd1 vssd1 vccd1 vccd1 net5117 sky130_fd_sc_hd__dlygate4sd3_1
X_17831_ _01815_ _02006_ _02067_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nand3_1
XFILLER_0_207_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17762_ _01919_ _01922_ _01920_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14974_ net4522 _08010_ _08079_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__mux2_1
X_19501_ net1396 net6546 _03365_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16713_ net7631 _09102_ vssd1 vssd1 vccd1 vccd1 _09751_ sky130_fd_sc_hd__xor2_2
X_13925_ _07095_ _06997_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nand2_2
X_17693_ _01930_ _01931_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19432_ net3658 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__clkbuf_1
X_13856_ _07024_ _07025_ _07026_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__nand3b_2
X_16644_ net4059 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12807_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19363_ _03268_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__buf_4
X_16575_ _08916_ _09664_ vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13787_ _06955_ _06956_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__and3_1
X_10999_ net1299 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18314_ net6150 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__clkbuf_1
X_15526_ _08609_ _08610_ _08620_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__a21oi_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _05904_ net34 vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ net5201 _03236_ _03243_ _03230_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__o211a_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15457_ _08207_ _08294_ _08306_ _08229_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__o22ai_1
X_18245_ _02450_ _02453_ _02451_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a21bo_1
X_12669_ reg_gpout\[3\] clknet_1_1__leaf__05847_ net45 vssd1 vssd1 vccd1 vccd1 _05848_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6909 rbzero.tex_g0\[35\] vssd1 vssd1 vccd1 vccd1 net7436 sky130_fd_sc_hd__dlygate4sd3_1
X_14408_ _07459_ _07578_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388_ _08479_ _08481_ _08482_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__and3_1
X_18176_ _02399_ net4526 _02393_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17127_ _10038_ _10053_ _10051_ vssd1 vssd1 vccd1 vccd1 _10147_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0__03865_ _03865_ vssd1 vssd1 vccd1 vccd1 clknet_0__03865_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ _07454_ _07509_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__xor2_2
Xhold505 net4836 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold516 net4841 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _01061_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold538 net6145 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ _10060_ _10061_ _10078_ vssd1 vssd1 vccd1 vccd1 _10079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 net6485 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16009_ _09103_ net7777 _08111_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _01046_ vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1216 _03393_ vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _00664_ vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1238 _03384_ vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 net3905 vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
X_20971_ clknet_leaf_108_i_clk net4069 vssd1 vssd1 vccd1 vccd1 reg_rgb\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21523_ clknet_leaf_3_i_clk net2077 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21454_ clknet_leaf_39_i_clk net2225 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20405_ clknet_1_0__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__buf_1
XFILLER_0_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21385_ clknet_leaf_6_i_clk net5175 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__buf_1
XFILLER_0_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__clkbuf_4
X_20267_ net4178 net4128 net4097 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__and3_1
Xhold3130 _03324_ vssd1 vssd1 vccd1 vccd1 net3657 sky130_fd_sc_hd__dlygate4sd3_1
X_22006_ net448 net768 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold3141 net4896 vssd1 vssd1 vccd1 vccd1 net3668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3152 _03776_ vssd1 vssd1 vccd1 vccd1 net3679 sky130_fd_sc_hd__dlygate4sd3_1
X_20198_ net3511 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
Xhold3163 net7480 vssd1 vssd1 vccd1 vccd1 net3690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3174 _02325_ vssd1 vssd1 vccd1 vccd1 net3701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2440 _01414_ vssd1 vssd1 vccd1 vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3185 net7645 vssd1 vssd1 vccd1 vccd1 net3712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2451 net2883 vssd1 vssd1 vccd1 vccd1 net2978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3196 net8333 vssd1 vssd1 vccd1 vccd1 net3723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2462 _01075_ vssd1 vssd1 vccd1 vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2473 _04188_ vssd1 vssd1 vccd1 vccd1 net3000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03854_ clknet_0__03854_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03854_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2484 _01153_ vssd1 vssd1 vccd1 vccd1 net3011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1750 net5604 vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2495 net7442 vssd1 vssd1 vccd1 vccd1 net3022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1761 net7014 vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ net3618 _05108_ net4160 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a21bo_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1772 _01591_ vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1783 _03487_ vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__clkbuf_2
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1794 net5995 vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__clkdlybuf4s25_1
X_13710_ _06707_ _06711_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__xor2_1
X_10922_ net7234 net7190 _04276_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__mux2_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _07776_ _07778_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__xor2_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _06772_ _06773_ _06811_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ net5664 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16360_ _09450_ net8520 vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__and2_1
X_13572_ _06683_ _06737_ net80 vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10784_ net7182 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__clkbuf_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _04511_ _08150_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__nand2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _05703_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__inv_2
X_16291_ _09381_ _09382_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _08285_ _08336_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__xnor2_4
X_18030_ _02165_ _02265_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__xnor2_1
X_12454_ _05633_ net4068 net8 _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ net3954 vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__inv_2
X_15173_ _08248_ _08267_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__xnor2_4
X_12385_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _05258_ vssd1 vssd1 vccd1 vccd1 _05570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _07263_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__inv_2
X_11336_ _04525_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19981_ net55 net7425 _03109_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _07224_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__nor2_2
X_18932_ net3363 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11267_ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006_ net4762 _06167_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__and2_1
X_18863_ net1863 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
X_11198_ net2457 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17814_ _01960_ _01961_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18794_ _02935_ _02936_ _02934_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17745_ _01760_ _08612_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14957_ net4789 net7825 _08068_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__mux2_1
X_13908_ _07074_ _07076_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__or3_1
X_17676_ _01914_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__nand2_1
X_14888_ _06237_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19415_ _08093_ net3570 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ net7752 _08115_ _09715_ _09716_ _01633_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__o221a_1
X_13839_ _06715_ _06755_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19346_ net6374 _03271_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__or2_1
X_16558_ _09646_ _09647_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15509_ _08567_ _08594_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__nor2_1
Xhold7407 net4288 vssd1 vssd1 vccd1 vccd1 net7934 sky130_fd_sc_hd__dlygate4sd3_1
X_19277_ net5368 _03200_ _03232_ _03230_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__o211a_1
Xhold7418 _01209_ vssd1 vssd1 vccd1 vccd1 net7945 sky130_fd_sc_hd__dlygate4sd3_1
X_16489_ _09577_ net7772 vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__and2_1
Xhold7429 net4566 vssd1 vssd1 vccd1 vccd1 net7956 sky130_fd_sc_hd__dlygate4sd3_1
X_18228_ _02434_ _02437_ _02435_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__o21a_1
Xhold6706 rbzero.tex_g0\[34\] vssd1 vssd1 vccd1 vccd1 net7233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6717 net2572 vssd1 vssd1 vccd1 vccd1 net7244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6728 _04308_ vssd1 vssd1 vccd1 vccd1 net7255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6739 net2524 vssd1 vssd1 vccd1 vccd1 net7266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18159_ _02383_ _02384_ _09872_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__o21ai_1
Xhold302 net5182 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 _03262_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03848_ _03848_ vssd1 vssd1 vccd1 vccd1 clknet_0__03848_ sky130_fd_sc_hd__clkbuf_16
Xhold324 net4251 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
X_21170_ clknet_leaf_132_i_clk net3113 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold335 net5184 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 net5401 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 net5375 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 net5409 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
X_20121_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold379 _01051_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _03650_ _03655_ net5784 _03484_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__a2bb2o_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 rbzero.tex_r1\[2\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _00578_ vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 net5519 vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1035 net6022 vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 net6559 vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1057 _00937_ vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1068 _00912_ vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 net6582 vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20954_ clknet_leaf_58_i_clk _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20885_ net4940 net63 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20493__236 clknet_1_0__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__inv_2
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7930 rbzero.texu_hot\[1\] vssd1 vssd1 vccd1 vccd1 net8457 sky130_fd_sc_hd__dlygate4sd3_1
X_21506_ clknet_leaf_11_i_clk net1696 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7974 _08407_ vssd1 vssd1 vccd1 vccd1 net8501 sky130_fd_sc_hd__buf_1
XFILLER_0_161_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21437_ clknet_leaf_18_i_clk net3219 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_leak
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12170_ _05276_ _05355_ _05357_ _04928_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21368_ clknet_leaf_14_i_clk net5019 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11121_ net5680 net5684 _04375_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20319_ net6677 net3674 _03825_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold880 _00979_ vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
X_21299_ clknet_leaf_43_i_clk net5007 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold891 _00995_ vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ net1408 net6219 _04342_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _08939_ _08952_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__o21ai_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2270 net975 vssd1 vssd1 vccd1 vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2281 _03534_ vssd1 vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
X_14811_ _07821_ _07830_ _07971_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__a21o_1
Xhold2292 _01515_ vssd1 vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _08882_ _08879_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__or2b_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1580 net6845 vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _01759_ _01770_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__xnor2_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1591 _01345_ vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
X_11954_ net4446 _05135_ _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a21oi_1
X_14742_ _07877_ _07878_ net7813 net7843 vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_104 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_104/HI o_rgb[13]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_115 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_115/HI zeros[4] sky130_fd_sc_hd__conb_1
XFILLER_0_153_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_126 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_126/HI zeros[15]
+ sky130_fd_sc_hd__conb_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_137 vssd1 vssd1 vccd1 vccd1 ones[10] top_ew_algofoogle_137/LO sky130_fd_sc_hd__conb_1
X_10905_ net6164 net2282 _04265_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17461_ _01700_ _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__nor2_1
X_14673_ _07820_ _07842_ _07843_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__a21o_1
X_11885_ net4105 _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19200_ net6697 _03183_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16412_ _09135_ _08167_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13624_ _06436_ _06637_ _06638_ _06642_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__a31o_2
X_10836_ net7007 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17392_ _08413_ _08612_ vssd1 vssd1 vccd1 vccd1 _10410_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19131_ _09721_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__clkbuf_4
X_16343_ _09433_ _09434_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__and2b_1
XFILLER_0_184_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ _06724_ net576 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10767_ net7139 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _05639_ _05686_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__o21a_2
X_16274_ _09363_ _09364_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__and2_1
X_19062_ net7601 net3631 net3397 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13486_ _06564_ _06579_ _06581_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__nand3_1
X_10698_ net6834 net5688 _04160_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15225_ net7776 _08129_ _08299_ _08319_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__o31a_1
X_18013_ net4742 _02248_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__xor2_1
X_12437_ _05026_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15156_ net4403 _08124_ _06119_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__a21o_1
X_12368_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _05258_ vssd1 vssd1 vccd1 vccd1 _05553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14107_ _07245_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11319_ net4181 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__clkbuf_8
X_19964_ net588 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
X_15087_ net8377 _06321_ net4181 vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ _04911_ _05482_ _05484_ _04919_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__o211a_1
X_14038_ _07207_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__nand2_1
X_18915_ net7546 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
X_19895_ net3096 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18846_ net5799 _02983_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18777_ _02866_ net4709 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__or2_1
X_15989_ _08992_ _09083_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__xor2_4
XFILLER_0_59_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ _01888_ _01964_ _01965_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17659_ _01760_ net8008 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19329_ net1343 _03237_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7204 _04908_ vssd1 vssd1 vccd1 vccd1 net7731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7215 rbzero.spi_registers.got_new_texadd\[0\] vssd1 vssd1 vccd1 vccd1 net7742
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold7237 rbzero.debug_overlay.playerX\[-7\] vssd1 vssd1 vccd1 vccd1 net7764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6503 _04187_ vssd1 vssd1 vccd1 vccd1 net7030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7248 _06026_ vssd1 vssd1 vccd1 vccd1 net7775 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold6514 net2510 vssd1 vssd1 vccd1 vccd1 net7041 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__05898_ clknet_0__05898_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05898_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7259 _06529_ vssd1 vssd1 vccd1 vccd1 net7786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6525 _04263_ vssd1 vssd1 vccd1 vccd1 net7052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6536 net2259 vssd1 vssd1 vccd1 vccd1 net7063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6547 rbzero.tex_b1\[11\] vssd1 vssd1 vccd1 vccd1 net7074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5802 net1261 vssd1 vssd1 vccd1 vccd1 net6329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5813 rbzero.spi_registers.new_texadd\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net6340
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6558 net836 vssd1 vssd1 vccd1 vccd1 net7085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6569 rbzero.tex_b1\[10\] vssd1 vssd1 vccd1 vccd1 net7096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5824 net1511 vssd1 vssd1 vccd1 vccd1 net6351 sky130_fd_sc_hd__dlygate4sd3_1
X_21222_ clknet_leaf_24_i_clk net3271 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold110 net4452 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5835 rbzero.spi_registers.new_texadd\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net6362
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 net4971 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold132 net4985 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5846 rbzero.spi_registers.new_texadd\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net6373
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5857 net1371 vssd1 vssd1 vccd1 vccd1 net6384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 net4996 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5868 net1319 vssd1 vssd1 vccd1 vccd1 net6395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold154 net8099 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold5879 rbzero.spi_registers.new_texadd\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net6406
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 net5050 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
X_21153_ clknet_leaf_122_i_clk net5847 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold176 net5036 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold187 net5054 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__inv_2
Xhold198 net5072 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
X_21084_ clknet_leaf_69_i_clk _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20035_ net5915 net3990 _03634_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ net428 net592 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20501__243 clknet_1_0__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__inv_2
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20937_ clknet_leaf_77_i_clk net4587 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11670_ net3365 _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__xnor2_1
X_20868_ _09739_ _02514_ net4715 _02508_ net8105 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10621_ net5708 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20799_ _03964_ _03965_ _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13340_ _06463_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__nand2_4
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ net5732 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _06438_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__or2_2
X_10483_ net7330 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7771 net654 vssd1 vssd1 vccd1 vccd1 net8298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7782 rbzero.row_render.size\[3\] vssd1 vssd1 vccd1 vccd1 net8309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7793 rbzero.wall_tracer.stepDistX\[9\] vssd1 vssd1 vccd1 vccd1 net8320 sky130_fd_sc_hd__dlygate4sd3_1
X_15010_ net4009 _08099_ net951 _06102_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__a2bb2o_1
X_12222_ _05407_ _05408_ _04930_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12153_ _05276_ _05338_ _05340_ _04928_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__o211a_1
X_11104_ net6273 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
X_12084_ _05213_ _05268_ _05270_ _05272_ _04942_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a221o_1
X_16961_ _09671_ _09683_ _09682_ vssd1 vssd1 vccd1 vccd1 _09983_ sky130_fd_sc_hd__a21bo_1
X_18700_ _02840_ _02852_ _02851_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a21o_1
X_11035_ net2937 net6442 _04331_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
X_15912_ _08255_ _08323_ _08553_ _08551_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__o31a_1
XFILLER_0_21_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19680_ net1553 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16892_ _09912_ _09913_ vssd1 vssd1 vccd1 vccd1 _09914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ net4528 net4635 _05164_ net4423 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__or4_2
XFILLER_0_95_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _08923_ _08937_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__and2_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _02729_ net7575 _06240_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _08417_ _08329_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__or2_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ net4498 vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__inv_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _01752_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nor2_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _07841_ _07856_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__nand2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _02642_ _02643_ _02668_ net4867 net4820 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a311o_1
X_11937_ net3473 _05100_ _05109_ net4052 vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20476__220 clknet_1_1__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__inv_2
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17444_ _09272_ _10096_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__nor2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14656_ _07822_ _07826_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__xor2_4
X_11868_ _04023_ _04468_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10819_ net2639 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13607_ _06762_ _06764_ _06763_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a21o_1
X_17375_ _10291_ _10306_ _10304_ vssd1 vssd1 vccd1 vccd1 _10393_ sky130_fd_sc_hd__a21o_1
X_11799_ _04984_ _04985_ _04987_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o211a_1
X_14587_ _07306_ _07457_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19114_ net4324 _03125_ net1062 _03128_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__o211a_1
X_16326_ net8041 _06122_ _09413_ _09417_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13538_ _06708_ _06697_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19045_ net3563 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__clkbuf_1
X_16257_ _09346_ _09348_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__nor2_1
X_13469_ _06445_ _06498_ _06639_ _06459_ _06528_ _06491_ vssd1 vssd1 vccd1 vccd1 _06640_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5109 net1950 vssd1 vssd1 vccd1 vccd1 net5636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15208_ net8021 _08119_ _06120_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16188_ _09279_ _09280_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4408 gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4419 net615 vssd1 vssd1 vccd1 vccd1 net4946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15139_ net4280 _08233_ _08122_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__mux2_1
Xhold3707 net8003 vssd1 vssd1 vccd1 vccd1 net4234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3718 net8306 vssd1 vssd1 vccd1 vccd1 net4245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3729 rbzero.wall_tracer.visualWallDist\[-1\] vssd1 vssd1 vccd1 vccd1 net4256
+ sky130_fd_sc_hd__clkbuf_1
X_19947_ net6239 net3286 _03583_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19878_ net3149 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18829_ net3486 _02971_ net5864 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21840_ net282 net2669 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21771_ clknet_leaf_45_i_clk net1461 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20722_ _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__and2b_1
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7001 rbzero.pov.spi_buffer\[12\] vssd1 vssd1 vccd1 vccd1 net7528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7012 rbzero.pov.spi_buffer\[16\] vssd1 vssd1 vccd1 vccd1 net7539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7023 net3276 vssd1 vssd1 vccd1 vccd1 net7550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7034 gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 net7561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6300 _04134_ vssd1 vssd1 vccd1 vccd1 net6827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7045 rbzero.pov.ready_buffer\[48\] vssd1 vssd1 vccd1 vccd1 net7572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6311 net1977 vssd1 vssd1 vccd1 vccd1 net6838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7056 net3711 vssd1 vssd1 vccd1 vccd1 net7583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6322 rbzero.tex_b0\[24\] vssd1 vssd1 vccd1 vccd1 net6849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7067 rbzero.pov.ready_buffer\[34\] vssd1 vssd1 vccd1 vccd1 net7594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6333 net2140 vssd1 vssd1 vccd1 vccd1 net6860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7078 net3345 vssd1 vssd1 vccd1 vccd1 net7605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6344 rbzero.tex_r1\[17\] vssd1 vssd1 vccd1 vccd1 net6871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7089 _03098_ vssd1 vssd1 vccd1 vccd1 net7616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6355 net2129 vssd1 vssd1 vccd1 vccd1 net6882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5610 _03836_ vssd1 vssd1 vccd1 vccd1 net6137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6366 rbzero.tex_b1\[51\] vssd1 vssd1 vccd1 vccd1 net6893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5621 net1505 vssd1 vssd1 vccd1 vccd1 net6148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6377 net1967 vssd1 vssd1 vccd1 vccd1 net6904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5632 rbzero.spi_registers.new_texadd\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net6159
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6388 _04131_ vssd1 vssd1 vccd1 vccd1 net6915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5643 net1084 vssd1 vssd1 vccd1 vccd1 net6170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5654 _03838_ vssd1 vssd1 vccd1 vccd1 net6181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6399 net2036 vssd1 vssd1 vccd1 vccd1 net6926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4920 rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 net5447 sky130_fd_sc_hd__dlygate4sd3_1
X_21205_ clknet_leaf_117_i_clk net2840 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5665 _02504_ vssd1 vssd1 vccd1 vccd1 net6192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5676 net1127 vssd1 vssd1 vccd1 vccd1 net6203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4931 net1119 vssd1 vssd1 vccd1 vccd1 net5458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5687 rbzero.tex_b0\[10\] vssd1 vssd1 vccd1 vccd1 net6214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4942 _00778_ vssd1 vssd1 vccd1 vccd1 net5469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5698 net1180 vssd1 vssd1 vccd1 vccd1 net6225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4953 net1228 vssd1 vssd1 vccd1 vccd1 net5480 sky130_fd_sc_hd__buf_1
Xhold4964 rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 net5491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21136_ clknet_leaf_31_i_clk net3886 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4975 _00882_ vssd1 vssd1 vccd1 vccd1 net5502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4986 net1582 vssd1 vssd1 vccd1 vccd1 net5513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4997 net1285 vssd1 vssd1 vccd1 vccd1 net5524 sky130_fd_sc_hd__dlygate4sd3_1
X_21067_ clknet_leaf_59_i_clk _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20018_ net4490 _08292_ _03614_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12840_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__inv_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _05947_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
XFILLER_0_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21969_ net411 net2520 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _04835_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__buf_4
XFILLER_0_178_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14510_ _07673_ _07674_ _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__a21o_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _08578_ _08583_ _08584_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ net5518 _04818_ _04821_ net5509 _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__o221a_1
X_14441_ _06725_ _07191_ _07192_ _07611_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__a31o_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ net2202 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17160_ _10079_ _10148_ _10178_ vssd1 vssd1 vccd1 vccd1 _10180_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14372_ _07517_ _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__and2_2
X_11584_ _04772_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16111_ _09073_ _09074_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ net7810 vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__clkbuf_1
X_10535_ net6985 net7192 _04075_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17091_ _09963_ _09985_ _09984_ vssd1 vssd1 vccd1 vccd1 _10112_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_80_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16042_ _08996_ _08864_ _09133_ _09135_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__a22o_1
X_13254_ _06383_ _06410_ _06418_ _06422_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__and4b_1
Xhold7590 rbzero.spi_registers.texadd2\[1\] vssd1 vssd1 vccd1 vccd1 net8117 sky130_fd_sc_hd__dlygate4sd3_1
X_10466_ net6838 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12205_ _05390_ _05391_ _04938_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13185_ _06018_ _06019_ _06266_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12136_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _04950_ vssd1 vssd1 vccd1 vccd1 _05324_
+ sky130_fd_sc_hd__mux2_1
X_17993_ _02228_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__nand2_1
X_19732_ net7676 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__clkbuf_1
X_20508__249 clknet_1_1__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__inv_2
X_12067_ rbzero.tex_r1\[45\] rbzero.tex_r1\[44\] _05249_ vssd1 vssd1 vccd1 vccd1 _05256_
+ sky130_fd_sc_hd__mux2_1
X_16944_ _09540_ _09541_ _08916_ vssd1 vssd1 vccd1 vccd1 _09966_ sky130_fd_sc_hd__a21oi_1
X_11018_ _04193_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19663_ net6474 net3897 _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
X_16875_ _09603_ _09896_ vssd1 vssd1 vccd1 vccd1 _09897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18614_ _02772_ _02773_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__or2b_1
X_15826_ _08919_ _08917_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__and2b_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ net6574 net3592 net1779 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18545_ _06057_ _06045_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__nor2_1
X_15757_ _08827_ _08850_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__nand2_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ net3893 _06133_ _06144_ _06098_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14708_ net7795 _07837_ _07838_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__and3_4
X_18476_ _02640_ _02646_ _02653_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15688_ _08220_ _08317_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17427_ _01666_ _01667_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14639_ _07795_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17358_ _10375_ _10376_ vssd1 vssd1 vccd1 vccd1 _10377_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ _09391_ _09400_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _10204_ _10277_ _10307_ vssd1 vssd1 vccd1 vccd1 _10308_ sky130_fd_sc_hd__a21o_1
X_19028_ net3864 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4205 net3429 vssd1 vssd1 vccd1 vccd1 net4732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4227 net3360 vssd1 vssd1 vccd1 vccd1 net4754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4238 _02823_ vssd1 vssd1 vccd1 vccd1 net4765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3504 _03081_ vssd1 vssd1 vccd1 vccd1 net4031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4249 net3626 vssd1 vssd1 vccd1 vccd1 net4776 sky130_fd_sc_hd__buf_2
XFILLER_0_167_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3515 _00726_ vssd1 vssd1 vccd1 vccd1 net4042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3526 _06067_ vssd1 vssd1 vccd1 vccd1 net4053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3537 _03076_ vssd1 vssd1 vccd1 vccd1 net4064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2803 _02994_ vssd1 vssd1 vccd1 vccd1 net3330 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_130_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold3548 _02483_ vssd1 vssd1 vccd1 vccd1 net4075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 rbzero.pov.spi_buffer\[29\] vssd1 vssd1 vccd1 vccd1 net3341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3559 _03991_ vssd1 vssd1 vccd1 vccd1 net4086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2825 _02995_ vssd1 vssd1 vccd1 vccd1 net3352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2836 _03033_ vssd1 vssd1 vccd1 vccd1 net3363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2847 net7728 vssd1 vssd1 vccd1 vccd1 net3374 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2858 net4548 vssd1 vssd1 vccd1 vccd1 net3385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2869 net4064 vssd1 vssd1 vccd1 vccd1 net3396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21823_ net265 net1951 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21754_ clknet_leaf_124_i_clk net3953 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20705_ _03884_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__xnor2_1
X_21685_ clknet_leaf_115_i_clk net4445 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20613__344 clknet_1_1__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__inv_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6130 net1797 vssd1 vssd1 vccd1 vccd1 net6657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6141 rbzero.tex_r0\[42\] vssd1 vssd1 vccd1 vccd1 net6668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6152 net1768 vssd1 vssd1 vccd1 vccd1 net6679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6163 _04041_ vssd1 vssd1 vccd1 vccd1 net6690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6174 net1661 vssd1 vssd1 vccd1 vccd1 net6701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6185 _04295_ vssd1 vssd1 vccd1 vccd1 net6712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5440 rbzero.row_render.side vssd1 vssd1 vccd1 vccd1 net5967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6196 net1782 vssd1 vssd1 vccd1 vccd1 net6723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5451 net3217 vssd1 vssd1 vccd1 vccd1 net5978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5462 _03593_ vssd1 vssd1 vccd1 vccd1 net5989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5473 net4101 vssd1 vssd1 vccd1 vccd1 net6000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5484 _03357_ vssd1 vssd1 vccd1 vccd1 net6011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5495 _03360_ vssd1 vssd1 vccd1 vccd1 net6022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4750 _00848_ vssd1 vssd1 vccd1 vccd1 net5277 sky130_fd_sc_hd__dlygate4sd3_1
X_22168_ clknet_leaf_91_i_clk net4942 vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4761 net993 vssd1 vssd1 vccd1 vccd1 net5288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4772 rbzero.spi_registers.texadd2\[12\] vssd1 vssd1 vccd1 vccd1 net5299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4783 net910 vssd1 vssd1 vccd1 vccd1 net5310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4794 _00822_ vssd1 vssd1 vccd1 vccd1 net5321 sky130_fd_sc_hd__dlygate4sd3_1
X_21119_ clknet_leaf_92_i_clk net4823 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_206_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22099_ net161 net2782 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
X_14990_ _08093_ net4156 vssd1 vssd1 vccd1 vccd1 _08094_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _06721_ _06693_ _06683_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _09738_ vssd1 vssd1 vccd1 vccd1 _09739_ sky130_fd_sc_hd__buf_4
X_13872_ _06702_ _06813_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__or2_1
X_15611_ _08694_ _08700_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12823_ _05976_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16591_ _08446_ _09680_ _09549_ _09550_ _09542_ vssd1 vssd1 vccd1 vccd1 _09681_ sky130_fd_sc_hd__a32o_1
XFILLER_0_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18330_ _02509_ _02517_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15542_ _08576_ _08629_ _08635_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__a21o_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12754_ net37 _05926_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__o21ai_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ net3940 net4814 net3906 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__and3b_1
X_11705_ net3014 _04467_ _04684_ net3151 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_182_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15473_ _08505_ _08499_ _08504_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__nand3_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ net31 _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__nor2_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17212_ _10218_ _10231_ vssd1 vssd1 vccd1 vccd1 _10232_ sky130_fd_sc_hd__xor2_1
X_11636_ _04799_ _04787_ _04796_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__nor3_1
X_14424_ _07589_ _07593_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03850_ clknet_0__03850_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03850_
+ sky130_fd_sc_hd__clkbuf_16
X_18192_ _02413_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17143_ _08413_ vssd1 vssd1 vccd1 vccd1 _10163_ sky130_fd_sc_hd__clkbuf_4
X_11567_ _04753_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nand2_1
X_14355_ _07242_ _07327_ _07523_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20588__321 clknet_1_1__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__inv_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10518_ net2373 net5637 _04064_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
X_13306_ _06466_ _06469_ _06471_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a31o_1
Xhold709 net6260 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
X_17074_ _09540_ _09541_ vssd1 vssd1 vccd1 vccd1 _10095_ sky130_fd_sc_hd__and2_1
X_14286_ _07145_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ _04682_ net3473 net3389 _04684_ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16025_ _08995_ _08999_ _09118_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__and3_1
X_13237_ net8002 _06266_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__or2_1
X_10449_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__nand2_1
X_12119_ _05300_ _05302_ _05305_ _05306_ _05263_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a221o_1
X_17976_ _02113_ _02123_ _02121_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a21oi_1
X_13099_ net4462 net3604 vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__nor2_1
Xhold1409 net6813 vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19715_ net3950 net4997 _08093_ _03485_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__o211a_1
X_16927_ _09941_ _09942_ _09947_ vssd1 vssd1 vccd1 vccd1 _09949_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_62_i_clk clknet_4_14__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19646_ net6303 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__clkbuf_1
X_16858_ _09809_ _09878_ _09879_ _09880_ vssd1 vssd1 vccd1 vccd1 _09881_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_205_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15809_ _08863_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19577_ net2645 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16789_ _09813_ _09816_ _09818_ vssd1 vssd1 vccd1 vccd1 _09819_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_77_i_clk clknet_4_13__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18528_ _02697_ _02698_ _02696_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18459_ rbzero.wall_tracer.rayAddendX\[4\] _02638_ _02537_ vssd1 vssd1 vccd1 vccd1
+ _02639_ sky130_fd_sc_hd__mux2_1
X_21470_ clknet_leaf_23_i_clk net1543 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4002 _02760_ vssd1 vssd1 vccd1 vccd1 net4529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4013 net7949 vssd1 vssd1 vccd1 vccd1 net4540 sky130_fd_sc_hd__dlygate4sd3_1
X_20283_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__buf_4
Xhold4024 _08051_ vssd1 vssd1 vccd1 vccd1 net4551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4035 _01238_ vssd1 vssd1 vccd1 vccd1 net4562 sky130_fd_sc_hd__dlygate4sd3_1
X_22022_ net464 net2045 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
Xhold4046 net2878 vssd1 vssd1 vccd1 vccd1 net4573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3301 net5883 vssd1 vssd1 vccd1 vccd1 net3828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4057 net4274 vssd1 vssd1 vccd1 vccd1 net4584 sky130_fd_sc_hd__clkbuf_2
Xhold3312 _03090_ vssd1 vssd1 vccd1 vccd1 net3839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4068 net8212 vssd1 vssd1 vccd1 vccd1 net4595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3323 _00614_ vssd1 vssd1 vccd1 vccd1 net3850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3334 net7980 vssd1 vssd1 vccd1 vccd1 net3861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4079 net792 vssd1 vssd1 vccd1 vccd1 net4606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2600 _01123_ vssd1 vssd1 vccd1 vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3345 _03994_ vssd1 vssd1 vccd1 vccd1 net3872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2611 net2838 vssd1 vssd1 vccd1 vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3356 _01212_ vssd1 vssd1 vccd1 vccd1 net3883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 _03548_ vssd1 vssd1 vccd1 vccd1 net3149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3367 _02710_ vssd1 vssd1 vccd1 vccd1 net3894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3378 rbzero.spi_registers.spi_done vssd1 vssd1 vccd1 vccd1 net3905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 _03588_ vssd1 vssd1 vccd1 vccd1 net3160 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2644 _01434_ vssd1 vssd1 vccd1 vccd1 net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03870_ clknet_0__03870_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03870_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3389 net4766 vssd1 vssd1 vccd1 vccd1 net3916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1910 _00751_ vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2655 rbzero.pov.ready_buffer\[22\] vssd1 vssd1 vccd1 vccd1 net3182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold58 net5789 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1921 _03366_ vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2666 _00716_ vssd1 vssd1 vccd1 vccd1 net3193 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2677 _01388_ vssd1 vssd1 vccd1 vccd1 net3204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 net7209 vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 net4933 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 _00654_ vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2688 _03563_ vssd1 vssd1 vccd1 vccd1 net3215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 _01043_ vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2699 rbzero.pov.spi_buffer\[49\] vssd1 vssd1 vccd1 vccd1 net3226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 _04303_ vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1976 net2476 vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1987 _01077_ vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1998 _04093_ vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21806_ net248 net1071 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21737_ clknet_leaf_98_i_clk net3512 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12470_ net54 _05643_ _05644_ net55 _05651_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21668_ clknet_leaf_123_i_clk net589 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _04536_ _04519_ _04534_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21599_ clknet_leaf_130_i_clk net1816 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14140_ _07307_ _07309_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11352_ _04506_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14071_ _06914_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__clkbuf_4
X_11283_ net3337 net92 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nand2_2
X_13022_ net4659 vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__inv_2
Xhold5270 _00629_ vssd1 vssd1 vccd1 vccd1 net5797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5281 _02788_ vssd1 vssd1 vccd1 vccd1 net5808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5292 _01168_ vssd1 vssd1 vccd1 vccd1 net5819 sky130_fd_sc_hd__dlygate4sd3_1
X_17830_ _01815_ _02006_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a21o_1
Xhold4580 net796 vssd1 vssd1 vccd1 vccd1 net5107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4591 _00837_ vssd1 vssd1 vccd1 vccd1 net5118 sky130_fd_sc_hd__dlygate4sd3_1
X_17761_ _01969_ _01999_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__xnor2_2
Xhold3890 _03745_ vssd1 vssd1 vccd1 vccd1 net4417 sky130_fd_sc_hd__dlygate4sd3_1
X_14973_ _08084_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19500_ net2448 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ net5554 _09102_ vssd1 vssd1 vccd1 vccd1 _09750_ sky130_fd_sc_hd__xor2_1
X_13924_ _06993_ _06995_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__nand2_1
X_17692_ _01930_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19431_ _03320_ net3657 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16643_ _04666_ net4058 _09727_ vssd1 vssd1 vccd1 vccd1 _09728_ sky130_fd_sc_hd__and3_1
X_13855_ _06960_ _06988_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ net7746 net4838 vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nand2_1
X_19362_ net5288 _03269_ _03282_ _03275_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16574_ _09411_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__clkbuf_4
X_10998_ net5653 net6345 _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__mux2_1
X_13786_ _06703_ _06914_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18313_ net6148 net3481 _02476_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
X_15525_ _08618_ _08619_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__or2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ net6058 _05912_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a21oi_2
X_19293_ net6299 _03238_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _02457_ net3588 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__nand2_1
X_15456_ _08207_ _08229_ _08294_ _08305_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__or4_1
X_12668_ net7571 _05800_ _05808_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_26_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ _06699_ _07391_ _07458_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__o21a_1
X_11619_ _04761_ _04763_ _04807_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a21oi_1
X_18175_ _02245_ net3667 _02398_ _10010_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a31o_1
X_15387_ _08467_ _08471_ _08478_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12599_ net20 _05755_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ _10144_ _10145_ vssd1 vssd1 vccd1 vccd1 _10146_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03864_ _03864_ vssd1 vssd1 vccd1 vccd1 clknet_0__03864_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14338_ _07506_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__and2_1
Xhold506 net6612 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold517 net4843 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold528 net7543 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _10067_ _10077_ vssd1 vssd1 vccd1 vccd1 _10078_ sky130_fd_sc_hd__xnor2_1
Xhold539 _01543_ vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14269_ _07438_ _07439_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_5__f_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16008_ _09102_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 net5993 vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 _00940_ vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 net6606 vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ _02194_ _02195_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__xnor2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1239 _00934_ vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
X_20642__370 clknet_1_0__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__inv_2
XFILLER_0_174_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20970_ clknet_leaf_111_i_clk net4158 vssd1 vssd1 vccd1 vccd1 reg_rgb\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19629_ net1279 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21522_ clknet_leaf_0_i_clk net1667 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21453_ clknet_leaf_36_i_clk net1744 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21384_ clknet_leaf_6_i_clk net5155 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20266_ _03352_ net4129 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__nor2_1
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__buf_1
Xhold3120 _00895_ vssd1 vssd1 vccd1 vccd1 net3647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22005_ net447 net2296 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold3131 _03325_ vssd1 vssd1 vccd1 vccd1 net3658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3142 net1680 vssd1 vssd1 vccd1 vccd1 net3669 sky130_fd_sc_hd__clkbuf_2
Xhold3153 _03777_ vssd1 vssd1 vccd1 vccd1 net3680 sky130_fd_sc_hd__dlygate4sd3_1
X_20197_ _03728_ net3510 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or2_1
Xhold3164 net7662 vssd1 vssd1 vccd1 vccd1 net3691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2430 _03004_ vssd1 vssd1 vccd1 vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3175 net8353 vssd1 vssd1 vccd1 vccd1 net3702 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2441 net5721 vssd1 vssd1 vccd1 vccd1 net2968 sky130_fd_sc_hd__buf_1
Xhold3186 _03742_ vssd1 vssd1 vccd1 vccd1 net3713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2452 _04374_ vssd1 vssd1 vccd1 vccd1 net2979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3197 net8335 vssd1 vssd1 vccd1 vccd1 net3724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2463 net5717 vssd1 vssd1 vccd1 vccd1 net2990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03853_ clknet_0__03853_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03853_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2474 _01458_ vssd1 vssd1 vccd1 vccd1 net3001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1740 _01361_ vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 net4906 vssd1 vssd1 vccd1 vccd1 net3012 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1751 net5606 vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2496 _03543_ vssd1 vssd1 vccd1 vccd1 net3023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1762 _04196_ vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
X_11970_ rbzero.debug_overlay.vplaneX\[10\] _05135_ _05154_ _05158_ vssd1 vssd1 vccd1
+ vccd1 _05159_ sky130_fd_sc_hd__a211o_1
Xhold1773 net7315 vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _03515_ vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ net3177 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
Xhold1795 net5997 vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10852_ net5662 net2462 _04238_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__mux2_1
X_13640_ _06727_ _06793_ _06774_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__and3_1
XFILLER_0_211_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ net2471 net7180 _04205_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
X_13571_ net79 _06734_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__nor2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _07991_ _08404_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__xnor2_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _05203_ _05698_ _05699_ net40 _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__a221o_1
X_16290_ _08308_ _08418_ _09380_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20470__215 clknet_1_1__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__inv_2
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15241_ _08287_ _08335_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__xor2_4
X_12453_ net7 vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _04503_ _04558_ _04592_ _04593_ _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o32a_1
X_15172_ _08255_ _08266_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__nor2_2
X_12384_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _05369_ vssd1 vssd1 vccd1 vccd1 _05569_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14123_ _07286_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__xnor2_1
X_11335_ _04523_ _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19980_ net3049 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18931_ net3125 net3362 _03025_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14054_ _07177_ _07201_ _07223_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__and3_1
X_11266_ net5946 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13005_ net4508 _06170_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18862_ net3045 net6681 _02993_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__mux2_1
X_11197_ net6987 net6096 _04423_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17813_ _02049_ _02050_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a21o_1
XFILLER_0_206_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18793_ net4838 _02537_ _09747_ _02937_ net8247 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__o221a_1
X_17744_ _01876_ _01877_ _01982_ _01762_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__o2bb2ai_2
X_14956_ _08075_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
X_13907_ _07048_ _07077_ _07000_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__a21oi_1
X_17675_ _01893_ _01894_ _01913_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__nand3_1
XFILLER_0_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _08035_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19414_ net1532 net3569 _03310_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__mux2_1
X_16626_ _09586_ _09714_ _08115_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__o21ai_1
X_13838_ _06964_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__xnor2_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19345_ net5041 _03269_ _03273_ _03259_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__o211a_1
X_16557_ _09644_ _09645_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _06927_ _06939_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15508_ _08597_ _08602_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19276_ net6132 _03202_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16488_ _09577_ net7772 vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__nor2_1
Xhold7408 rbzero.wall_tracer.trackDistY\[-10\] vssd1 vssd1 vccd1 vccd1 net7935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7419 net4410 vssd1 vssd1 vccd1 vccd1 net7946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18227_ _02442_ _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__or2b_1
X_15439_ _06122_ net8008 vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__or2_1
Xhold6707 net2731 vssd1 vssd1 vccd1 vccd1 net7234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6718 _04405_ vssd1 vssd1 vccd1 vccd1 net7245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6729 net2671 vssd1 vssd1 vccd1 vccd1 net7256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18158_ _02382_ _02380_ _02381_ _06057_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold303 net5403 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17109_ _10128_ _10129_ vssd1 vssd1 vccd1 vccd1 _10130_ sky130_fd_sc_hd__or2_2
Xhold314 net4196 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03847_ _03847_ vssd1 vssd1 vccd1 vccd1 clknet_0__03847_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 net5227 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ net4518 net4351 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold336 net5186 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold347 net5315 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 net5377 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
X_20120_ net4997 _03122_ _03484_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold369 net8122 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20051_ net4019 _03484_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__or2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 net5551 vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 net3595 vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 net6398 vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _00916_ vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 _02998_ vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 net8359 vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 net6292 vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ clknet_leaf_58_i_clk _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ net4848 _02508_ _02559_ _04015_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a22o_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21505_ clknet_leaf_12_i_clk net1339 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7920 net4775 vssd1 vssd1 vccd1 vccd1 net8447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21436_ clknet_leaf_40_i_clk net2148 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7964 net5902 vssd1 vssd1 vccd1 vccd1 net8491 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21367_ clknet_leaf_18_i_clk net5346 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ net2931 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20318_ net6498 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
Xhold870 _02480_ vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
X_21298_ clknet_leaf_43_i_clk net5238 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold881 net6523 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net2358 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
Xhold892 net6389 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
X_20249_ _04464_ _04684_ _04749_ net5207 net900 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a41o_1
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2260 net7288 vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2271 _04068_ vssd1 vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
X_14810_ _07821_ _07874_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2282 _01101_ vssd1 vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _08860_ _08884_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__or2_1
Xhold2293 net7261 vssd1 vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1570 rbzero.spi_registers.new_vshift\[3\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1581 net6847 vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ net7850 _07905_ _07906_ _07908_ net7839 vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__a311o_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1592 net6688 vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ rbzero.debug_overlay.facingX\[-2\] _05080_ _05136_ _05141_ vssd1 vssd1 vccd1
+ vccd1 _05142_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_105 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_105/HI o_rgb[16]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_116 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_116/HI zeros[5] sky130_fd_sc_hd__conb_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_127 vssd1 vssd1 vccd1 vccd1 ones[0] top_ew_algofoogle_127/LO sky130_fd_sc_hd__conb_1
X_10904_ net2454 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__clkbuf_1
X_17460_ _10345_ _10354_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a21oi_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_138 vssd1 vssd1 vccd1 vccd1 ones[11] top_ew_algofoogle_138/LO sky130_fd_sc_hd__conb_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ net7850 vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ _04666_ net4058 _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and3_1
X_16411_ _08996_ _08167_ _09373_ _09135_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__a22o_1
X_13623_ _06729_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ net7005 net2848 _04227_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_1
X_17391_ _10408_ _09062_ vssd1 vssd1 vccd1 vccd1 _10409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19130_ net1289 _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__or2_1
X_16342_ _09430_ _09432_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _06722_ _06723_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__o21ai_4
X_10766_ net7137 net2376 _04194_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19061_ net7599 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__clkbuf_1
X_12505_ net4149 _05641_ _05640_ _05646_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__nand4b_1
X_16273_ _09363_ _09364_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10697_ net3357 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__clkbuf_1
X_13485_ _06564_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18012_ _02241_ _02243_ _02240_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a21bo_1
X_15224_ net8269 _08129_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ net4321 _04848_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _07929_ net8418 _08113_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__mux2_1
X_12367_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _05369_ vssd1 vssd1 vccd1 vccd1 _05552_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14106_ _07275_ _07276_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__nand2_2
X_11318_ net4180 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__clkbuf_2
X_12298_ _04938_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__or2_1
X_15086_ _08162_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__clkbuf_8
X_19963_ net5988 net3237 _03583_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ net7023 net6969 _04445_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__mux2_1
X_14037_ _07160_ _07206_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__or2_1
X_18914_ net3179 net7544 _03014_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19894_ net3298 net3125 _03550_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18845_ net5864 net3486 _02985_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18776_ _02915_ _02916_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or2b_1
X_15988_ _09081_ _09082_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__and2_4
XFILLER_0_136_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17727_ _01888_ _01964_ _01965_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a21oi_2
X_14939_ _08037_ net1792 net4332 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17658_ _01896_ _01897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__and2_1
X_16609_ _09696_ _09697_ vssd1 vssd1 vccd1 vccd1 _09699_ sky130_fd_sc_hd__and2_1
X_17589_ _01828_ _01829_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19328_ net8116 _03250_ net840 _03259_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7205 rbzero.color_sky\[3\] vssd1 vssd1 vccd1 vccd1 net7732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7216 gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 net7743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19259_ net986 _03217_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7238 net3348 vssd1 vssd1 vccd1 vccd1 net7765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6504 net2418 vssd1 vssd1 vccd1 vccd1 net7031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7249 _06027_ vssd1 vssd1 vccd1 vccd1 net7776 sky130_fd_sc_hd__buf_2
Xhold6515 rbzero.tex_g1\[9\] vssd1 vssd1 vccd1 vccd1 net7042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6526 net1965 vssd1 vssd1 vccd1 vccd1 net7053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6537 _04056_ vssd1 vssd1 vccd1 vccd1 net7064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5803 rbzero.spi_registers.new_texadd\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net6330
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6548 net2664 vssd1 vssd1 vccd1 vccd1 net7075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6559 rbzero.tex_r1\[26\] vssd1 vssd1 vccd1 vccd1 net7086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 net4720 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
X_21221_ clknet_leaf_24_i_clk net3413 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5814 net1337 vssd1 vssd1 vccd1 vccd1 net6341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5825 _03467_ vssd1 vssd1 vccd1 vccd1 net6352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold111 net8102 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5836 net1514 vssd1 vssd1 vccd1 vccd1 net6363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 net4973 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5847 net1368 vssd1 vssd1 vccd1 vccd1 net6374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 net6051 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5858 _02500_ vssd1 vssd1 vccd1 vccd1 net6385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 net4998 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
X_21152_ clknet_leaf_106_i_clk net3613 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5869 _03406_ vssd1 vssd1 vccd1 vccd1 net6396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 net4601 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 net8104 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 net5038 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ net3473 _03690_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__or2_1
Xhold188 net4987 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 net5074 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
X_21083_ clknet_leaf_69_i_clk _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20034_ net3993 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ net427 net1750 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ clknet_leaf_76_i_clk net4579 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _02511_ net4714 _02512_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a21bo_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ net5706 net5577 _04116_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
X_20798_ net1015 net5522 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10551_ net5659 net5730 _04075_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ net3128 net7328 _04042_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__mux2_1
X_13270_ _06439_ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7783 net4302 vssd1 vssd1 vccd1 vccd1 net8310 sky130_fd_sc_hd__dlygate4sd3_1
X_12221_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _04950_ vssd1 vssd1 vccd1 vccd1 _05408_
+ sky130_fd_sc_hd__mux2_1
Xhold7794 net4387 vssd1 vssd1 vccd1 vccd1 net8321 sky130_fd_sc_hd__dlygate4sd3_1
X_21419_ clknet_leaf_40_i_clk net2323 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ _04976_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20582__316 clknet_1_1__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__inv_2
X_11103_ net2664 net6271 _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16960_ _09979_ _09980_ _09968_ vssd1 vssd1 vccd1 vccd1 _09982_ sky130_fd_sc_hd__a21o_1
X_12083_ _04911_ _05271_ _04988_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11034_ net2001 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
X_15911_ _09004_ _09005_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__xnor2_1
X_16891_ _08226_ _09116_ vssd1 vssd1 vccd1 vccd1 _09913_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18630_ net5809 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _08915_ _08922_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__or2_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2090 _04282_ vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ net3469 _02728_ _02245_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _08862_ _08867_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__xor2_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ net4646 _06124_ net4781 vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__o21a_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17512_ _10398_ _10399_ _10397_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a21oi_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14724_ _07893_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__clkbuf_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] _02617_
+ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__o21a_1
X_11936_ net4188 _05103_ _05115_ net3469 _05124_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a221o_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _01683_ _01684_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nand2_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14655_ _07808_ _07824_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__a21o_2
XFILLER_0_68_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11867_ net4147 net4066 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__or2_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13606_ _06721_ _06730_ _06728_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__and3_1
X_17374_ _10390_ _10391_ vssd1 vssd1 vccd1 vccd1 _10392_ sky130_fd_sc_hd__nor2_1
X_10818_ net6478 net7293 _04216_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14586_ _07489_ _07391_ _07752_ _07756_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__o31a_1
X_11798_ net87 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19113_ net1061 _03126_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16325_ _09415_ _09416_ _08441_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__o21ai_4
X_13537_ _06634_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__clkbuf_4
X_10749_ net7264 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ net3562 net3738 net3398 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
X_16256_ _09226_ _09347_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__nor2_1
X_13468_ _06461_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15207_ _08301_ net4188 _06027_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__mux2_2
X_12419_ rbzero.tex_b1\[57\] rbzero.tex_b1\[56\] _05258_ vssd1 vssd1 vccd1 vccd1 _05604_
+ sky130_fd_sc_hd__mux2_1
X_16187_ _09277_ _09278_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__nor2_1
X_13399_ _06430_ _06551_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4409 net600 vssd1 vssd1 vccd1 vccd1 net4936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _08232_ net3317 _06027_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3708 net1016 vssd1 vssd1 vccd1 vccd1 net4235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3719 net8308 vssd1 vssd1 vccd1 vccd1 net4246 sky130_fd_sc_hd__dlygate4sd3_1
X_19946_ net2904 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
X_15069_ _07962_ net8372 _08113_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__mux2_2
X_19877_ net3195 net7556 _03539_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18828_ net5863 net2182 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__or2b_1
X_18759_ _02881_ _02882_ _02906_ net4856 net4807 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21770_ clknet_leaf_11_i_clk net1306 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20721_ net1048 net5404 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7002 rbzero.tex_b1\[20\] vssd1 vssd1 vccd1 vccd1 net7529 sky130_fd_sc_hd__dlygate4sd3_1
X_20583_ clknet_1_1__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__buf_1
Xhold7013 net3063 vssd1 vssd1 vccd1 vccd1 net7540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7024 rbzero.pov.ready_buffer\[27\] vssd1 vssd1 vccd1 vccd1 net7551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7035 net4057 vssd1 vssd1 vccd1 vccd1 net7562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6301 net1518 vssd1 vssd1 vccd1 vccd1 net6828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7046 net3414 vssd1 vssd1 vccd1 vccd1 net7573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6312 rbzero.tex_r0\[27\] vssd1 vssd1 vccd1 vccd1 net6839 sky130_fd_sc_hd__dlygate4sd3_1
X_20334__92 clknet_1_0__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__inv_2
Xhold7057 rbzero.spi_registers.spi_buffer\[19\] vssd1 vssd1 vccd1 vccd1 net7584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6323 net1758 vssd1 vssd1 vccd1 vccd1 net6850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7068 net2242 vssd1 vssd1 vccd1 vccd1 net7595 sky130_fd_sc_hd__buf_1
Xhold6334 rbzero.spi_registers.new_texadd\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 net6861
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold7079 _03654_ vssd1 vssd1 vccd1 vccd1 net7606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5600 rbzero.tex_b1\[26\] vssd1 vssd1 vccd1 vccd1 net6127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6345 net2020 vssd1 vssd1 vccd1 vccd1 net6872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6356 rbzero.tex_g0\[50\] vssd1 vssd1 vccd1 vccd1 net6883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5611 net1400 vssd1 vssd1 vccd1 vccd1 net6138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5622 _02505_ vssd1 vssd1 vccd1 vccd1 net6149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6367 net2063 vssd1 vssd1 vccd1 vccd1 net6894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6378 rbzero.tex_r0\[58\] vssd1 vssd1 vccd1 vccd1 net6905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5633 net1599 vssd1 vssd1 vccd1 vccd1 net6160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5644 rbzero.tex_r0\[44\] vssd1 vssd1 vccd1 vccd1 net6171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6389 net2424 vssd1 vssd1 vccd1 vccd1 net6916 sky130_fd_sc_hd__dlygate4sd3_1
X_21204_ clknet_leaf_116_i_clk net2760 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4910 _00805_ vssd1 vssd1 vccd1 vccd1 net5437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5655 net1220 vssd1 vssd1 vccd1 vccd1 net6182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4921 net1046 vssd1 vssd1 vccd1 vccd1 net5448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5666 net1344 vssd1 vssd1 vccd1 vccd1 net6193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5677 _04195_ vssd1 vssd1 vccd1 vccd1 net6204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4932 rbzero.floor_leak\[1\] vssd1 vssd1 vccd1 vccd1 net5459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4943 net1164 vssd1 vssd1 vccd1 vccd1 net5470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5688 net1148 vssd1 vssd1 vccd1 vccd1 net6215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5699 rbzero.tex_g1\[58\] vssd1 vssd1 vccd1 vccd1 net6226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4954 _01620_ vssd1 vssd1 vccd1 vccd1 net5481 sky130_fd_sc_hd__dlygate4sd3_1
X_21135_ clknet_leaf_29_i_clk net4051 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4965 net1233 vssd1 vssd1 vccd1 vccd1 net5492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4976 net1256 vssd1 vssd1 vccd1 vccd1 net5503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4987 _03337_ vssd1 vssd1 vccd1 vccd1 net5514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4998 rbzero.spi_registers.new_other\[0\] vssd1 vssd1 vccd1 vccd1 net5525 sky130_fd_sc_hd__dlygate4sd3_1
X_21066_ clknet_leaf_61_i_clk _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20017_ net3457 _03607_ net5851 _03628_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__o211a_1
X_20425__175 clknet_1_0__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__inv_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ reg_gpout\[5\] clknet_1_1__leaf__05946_ net45 vssd1 vssd1 vccd1 vccd1 _05947_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ net410 net1452 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__clkbuf_8
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ clknet_leaf_77_i_clk _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21899_ net341 net2591 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14440_ _07308_ _07197_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__nor2_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ net1255 _04825_ _04817_ net1550 _04841_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a221o_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ net7135 net7067 _04105_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__mux2_1
X_14371_ _07514_ _07515_ _07516_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ net1086 net1851 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16110_ _09070_ _09203_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__buf_4
X_17090_ _10094_ _10110_ vssd1 vssd1 vccd1 vccd1 _10111_ sky130_fd_sc_hd__xnor2_2
X_10534_ _04030_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16041_ _06123_ net8072 vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__nor2_2
X_10465_ net2851 net6836 _04031_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13253_ _06415_ _06417_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__mux2_1
Xhold7591 net4198 vssd1 vssd1 vccd1 vccd1 net8118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _04916_ vssd1 vssd1 vccd1 vccd1 _05391_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6890 net2654 vssd1 vssd1 vccd1 vccd1 net7417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13184_ _04491_ _06314_ _06316_ _06319_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_209_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ _05317_ _05319_ _05322_ _04928_ _04942_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17992_ _02222_ _02227_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__or2_1
X_16943_ _09666_ _09667_ _08401_ vssd1 vssd1 vccd1 vccd1 _09965_ sky130_fd_sc_hd__a21oi_1
X_19731_ net7674 _03493_ net3708 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ rbzero.tex_r1\[47\] rbzero.tex_r1\[46\] _05249_ vssd1 vssd1 vccd1 vccd1 _05255_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11017_ net2546 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
X_16874_ _08542_ _09345_ vssd1 vssd1 vccd1 vccd1 _09896_ sky130_fd_sc_hd__nor2_1
X_19662_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__buf_4
X_15825_ _08917_ _08919_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__and2b_1
X_18613_ net3575 net5925 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nand2_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ net1780 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _08827_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__xor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _06038_ _06042_ _06044_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__or3_1
X_12968_ _06104_ net4034 _06134_ _06143_ _06129_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a311o_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14707_ net7795 _07837_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__nor2_2
XFILLER_0_206_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18475_ _02617_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _02653_
+ sky130_fd_sc_hd__xnor2_2
X_11919_ _05107_ _05077_ _05099_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_2
X_15687_ _08266_ _08341_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__or2_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ net3683 net4049 _06063_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__a211o_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _01666_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14638_ net8355 _07806_ _07807_ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__o31a_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17357_ _10269_ _10270_ _10374_ vssd1 vssd1 vccd1 vccd1 _10376_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14569_ _07712_ _07715_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _09398_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__nand2_1
X_17288_ _10291_ _10306_ vssd1 vssd1 vccd1 vccd1 _10307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19027_ net2205 net3863 _03078_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
X_16239_ _09330_ _09331_ vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4206 net8253 vssd1 vssd1 vccd1 vccd1 net4733 sky130_fd_sc_hd__buf_2
XFILLER_0_207_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4217 net8205 vssd1 vssd1 vccd1 vccd1 net4744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20565__300 clknet_1_0__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__inv_2
Xhold4228 net7814 vssd1 vssd1 vccd1 vccd1 net4755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4239 net8095 vssd1 vssd1 vccd1 vccd1 net4766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3505 _00723_ vssd1 vssd1 vccd1 vccd1 net4032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3516 net8272 vssd1 vssd1 vccd1 vccd1 net4043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3527 _02713_ vssd1 vssd1 vccd1 vccd1 net4054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3538 net5964 vssd1 vssd1 vccd1 vccd1 net4065 sky130_fd_sc_hd__buf_1
Xhold2804 _00647_ vssd1 vssd1 vccd1 vccd1 net3331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3549 net1426 vssd1 vssd1 vccd1 vccd1 net4076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 net3292 vssd1 vssd1 vccd1 vccd1 net3342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2826 _00648_ vssd1 vssd1 vccd1 vccd1 net3353 sky130_fd_sc_hd__dlygate4sd3_1
X_19929_ net3053 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
Xhold2837 _00683_ vssd1 vssd1 vccd1 vccd1 net3364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2848 _03138_ vssd1 vssd1 vccd1 vccd1 net3375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2859 net8251 vssd1 vssd1 vccd1 vccd1 net3386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21822_ net264 net2216 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21753_ clknet_leaf_101_i_clk net5047 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20704_ _03885_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21684_ clknet_leaf_114_i_clk net3546 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6120 net1923 vssd1 vssd1 vccd1 vccd1 net6647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6131 _04361_ vssd1 vssd1 vccd1 vccd1 net6658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6142 net1848 vssd1 vssd1 vccd1 vccd1 net6669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6153 rbzero.pov.ready_buffer\[3\] vssd1 vssd1 vccd1 vccd1 net6680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6164 net2120 vssd1 vssd1 vccd1 vccd1 net6691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6175 rbzero.tex_r0\[25\] vssd1 vssd1 vccd1 vccd1 net6702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5430 net3612 vssd1 vssd1 vccd1 vccd1 net5957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5441 net4079 vssd1 vssd1 vccd1 vccd1 net5968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6186 net2111 vssd1 vssd1 vccd1 vccd1 net6713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6197 _04290_ vssd1 vssd1 vccd1 vccd1 net6724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5452 _03372_ vssd1 vssd1 vccd1 vccd1 net5979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5463 rbzero.tex_r0\[4\] vssd1 vssd1 vccd1 vccd1 net5990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5474 _03795_ vssd1 vssd1 vccd1 vccd1 net6001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5485 net1565 vssd1 vssd1 vccd1 vccd1 net6012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4740 rbzero.spi_registers.texadd2\[3\] vssd1 vssd1 vccd1 vccd1 net5267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5496 rbzero.spi_registers.new_floor\[4\] vssd1 vssd1 vccd1 vccd1 net6023 sky130_fd_sc_hd__dlygate4sd3_1
X_22167_ clknet_leaf_96_i_clk net4850 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4751 net899 vssd1 vssd1 vccd1 vccd1 net5278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4762 _00864_ vssd1 vssd1 vccd1 vccd1 net5289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4773 net856 vssd1 vssd1 vccd1 vccd1 net5300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4784 rbzero.spi_registers.texadd3\[7\] vssd1 vssd1 vccd1 vccd1 net5311 sky130_fd_sc_hd__dlygate4sd3_1
X_21118_ clknet_leaf_92_i_clk net3814 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4795 net945 vssd1 vssd1 vccd1 vccd1 net5322 sky130_fd_sc_hd__dlygate4sd3_1
X_22098_ net160 net2690 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13940_ _07108_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__xor2_1
X_21049_ clknet_leaf_78_i_clk _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13871_ _07010_ _07041_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__xnor2_1
X_15610_ _08699_ _08697_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__and2b_1
X_12822_ _05975_ _05969_ _05973_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nand3_1
X_16590_ _09676_ _09546_ _06124_ vssd1 vssd1 vccd1 vccd1 _09680_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15541_ _08576_ _08629_ _08635_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__nand3_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12753_ net35 _05927_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21ai_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ net1879 _02472_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__nor2_1
X_11704_ net3151 _04684_ _04465_ net3488 _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
X_15472_ _08565_ _08566_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__or2_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ net30 vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__inv_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _10229_ _10230_ vssd1 vssd1 vccd1 vccd1 _10231_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _07589_ _07593_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__xnor2_2
X_11635_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__buf_4
X_18191_ _02412_ net3766 _02393_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17142_ _09617_ _10042_ _10043_ _10044_ vssd1 vssd1 vccd1 vccd1 _10162_ sky130_fd_sc_hd__o2bb2ai_1
X_14354_ _07523_ _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_182_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11566_ net1079 net1228 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13305_ _06467_ net574 _06468_ _06475_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17073_ _10083_ _10093_ vssd1 vssd1 vccd1 vccd1 _10094_ sky130_fd_sc_hd__xnor2_2
X_10517_ net5647 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__clkbuf_1
X_14285_ _07410_ _07426_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__xnor2_1
X_11497_ net4091 net3553 _04686_ _04460_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__o22a_1
X_16024_ _09113_ _09117_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13236_ _06399_ _06401_ _06403_ _06406_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or4_4
XFILLER_0_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10448_ _04021_ _04027_ net92 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and3_2
XFILLER_0_23_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ rbzero.wall_tracer.visualWallDist\[-8\] _06009_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ _04955_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17975_ _02201_ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__xnor2_2
X_13098_ net4513 net6015 vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__or2_2
X_19714_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16926_ _09941_ _09942_ _09947_ vssd1 vssd1 vccd1 vccd1 _09948_ sky130_fd_sc_hd__a21oi_1
X_12049_ rbzero.tex_r1\[25\] rbzero.tex_r1\[24\] _05237_ vssd1 vssd1 vccd1 vccd1 _05238_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19645_ net6301 net3556 _03441_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__mux2_1
X_16857_ _09818_ _09711_ vssd1 vssd1 vccd1 vccd1 _09880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20560__296 clknet_1_1__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__inv_2
XFILLER_0_137_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19785__64 clknet_1_1__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
XFILLER_0_205_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15808_ _08866_ _08865_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__or2b_1
XFILLER_0_153_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19576_ net7522 net3863 _03403_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
X_16788_ net4865 vssd1 vssd1 vccd1 vccd1 _09818_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15739_ _08229_ _08458_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__nor2_1
X_18527_ net4828 _02537_ _09747_ _02699_ _02701_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18458_ _02629_ _02637_ _02526_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17409_ _10425_ _10426_ vssd1 vssd1 vccd1 vccd1 _10427_ sky130_fd_sc_hd__nand2_1
X_18389_ _02570_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4003 _02761_ vssd1 vssd1 vccd1 vccd1 net4530 sky130_fd_sc_hd__dlygate4sd3_1
X_20282_ _04102_ net4816 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__nor2_4
Xhold4014 net3764 vssd1 vssd1 vccd1 vccd1 net4541 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4025 _00422_ vssd1 vssd1 vccd1 vccd1 net4552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22021_ net463 net2103 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
Xhold4036 net646 vssd1 vssd1 vccd1 vccd1 net4563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3302 net5885 vssd1 vssd1 vccd1 vccd1 net3829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4047 net7959 vssd1 vssd1 vccd1 vccd1 net4574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3313 _00731_ vssd1 vssd1 vccd1 vccd1 net3840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4058 _08054_ vssd1 vssd1 vccd1 vccd1 net4585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4069 _01204_ vssd1 vssd1 vccd1 vccd1 net4596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3324 net3939 vssd1 vssd1 vccd1 vccd1 net3851 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3335 net3876 vssd1 vssd1 vccd1 vccd1 net3862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2601 net7358 vssd1 vssd1 vccd1 vccd1 net3128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3346 _01625_ vssd1 vssd1 vccd1 vccd1 net3873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2612 _03568_ vssd1 vssd1 vccd1 vccd1 net3139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3357 net7630 vssd1 vssd1 vccd1 vccd1 net3884 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2623 _01114_ vssd1 vssd1 vccd1 vccd1 net3150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3368 _00612_ vssd1 vssd1 vccd1 vccd1 net3895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3379 net1776 vssd1 vssd1 vccd1 vccd1 net3906 sky130_fd_sc_hd__buf_1
Xhold2634 _01150_ vssd1 vssd1 vccd1 vccd1 net3161 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2645 rbzero.pov.spi_buffer\[24\] vssd1 vssd1 vccd1 vccd1 net3172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1900 _03052_ vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1911 net7327 vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2656 net7444 vssd1 vssd1 vccd1 vccd1 net3183 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1922 _00918_ vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2667 rbzero.pov.spi_buffer\[27\] vssd1 vssd1 vccd1 vccd1 net3194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 _01573_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1933 _04210_ vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 net7966 vssd1 vssd1 vccd1 vccd1 net3205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1944 net7398 vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 _01127_ vssd1 vssd1 vccd1 vccd1 net3216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1955 net7360 vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1966 _01355_ vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1977 _04247_ vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1988 net7152 vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1999 _01541_ vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21805_ net247 net2308 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21736_ clknet_leaf_95_i_clk net3664 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20537__276 clknet_1_0__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__inv_2
XFILLER_0_152_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21667_ clknet_leaf_121_i_clk net1569 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11420_ _04021_ _04607_ _04609_ _04611_ _04494_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a221o_2
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21598_ net232 net1969 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11351_ _04515_ _04540_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a21oi_1
X_20549_ clknet_1_0__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__buf_1
XFILLER_0_160_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14070_ _07240_ _07194_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11282_ net4186 vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5260 rbzero.tex_r1\[40\] vssd1 vssd1 vccd1 vccd1 net5787 sky130_fd_sc_hd__dlygate4sd3_1
X_13021_ _06191_ net3820 _06193_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5271 rbzero.spi_registers.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 net5798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5282 net3527 vssd1 vssd1 vccd1 vccd1 net5809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5293 net3537 vssd1 vssd1 vccd1 vccd1 net5820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4570 net733 vssd1 vssd1 vccd1 vccd1 net5097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4581 rbzero.spi_registers.texadd1\[17\] vssd1 vssd1 vccd1 vccd1 net5108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4592 net761 vssd1 vssd1 vccd1 vccd1 net5119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3880 net3488 vssd1 vssd1 vccd1 vccd1 net4407 sky130_fd_sc_hd__dlygate4sd3_1
X_17760_ _01997_ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__nand2_1
X_14972_ net4405 _08004_ _08079_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__mux2_1
Xhold3891 _01216_ vssd1 vssd1 vccd1 vccd1 net4418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13923_ net3503 _07029_ _07091_ _07093_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ net7611 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
X_17691_ _01805_ _01825_ _01823_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19430_ net1480 net3656 _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__mux2_1
X_16642_ _04458_ net4122 vssd1 vssd1 vccd1 vccd1 _09727_ sky130_fd_sc_hd__nor2_4
XFILLER_0_201_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13854_ _06982_ _06984_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__xor2_2
XFILLER_0_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12805_ net7746 net5955 vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__nor2_1
X_16573_ _09655_ _09662_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__xor2_1
X_19361_ net6309 _03271_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _06706_ net3634 vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__nor2_1
X_10997_ _04193_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15524_ _08615_ _08617_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__and2_1
X_18312_ net6193 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19292_ net5268 _03236_ _03242_ _03230_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__o211a_1
X_12736_ net144 net35 _05901_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ net3926 net4608 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__or2_1
X_15455_ _08548_ _08549_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _05828_ _05845_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14406_ _07570_ _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11618_ _04807_ _04761_ _04763_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand3_1
X_18174_ net3666 _02390_ _02395_ _02396_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15386_ _08388_ _08480_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ _05776_ _05777_ net19 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _10055_ _10141_ _10143_ vssd1 vssd1 vccd1 vccd1 _10145_ sky130_fd_sc_hd__and3_1
Xclkbuf_0__03863_ _03863_ vssd1 vssd1 vccd1 vccd1 clknet_0__03863_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ _07434_ _07507_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__nor2_2
XFILLER_0_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11549_ net3983 _04022_ _04600_ _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a22o_1
Xhold507 _03336_ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 net4845 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17056_ _10075_ _10076_ vssd1 vssd1 vccd1 vccd1 _10077_ sky130_fd_sc_hd__and2b_1
Xhold529 net4488 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ _07240_ _07242_ _07305_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__or3_2
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16007_ _08194_ vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__buf_4
X_13219_ _06356_ _06357_ _06361_ net8217 vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__a22o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _07368_ _07369_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__nand2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1207 _03346_ vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _09413_ _10163_ net7837 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__or3b_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 net6628 vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 net6608 vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16909_ _09639_ _09647_ _09646_ vssd1 vssd1 vccd1 vccd1 _09931_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17889_ _02124_ _02125_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__and2_1
X_19628_ net6281 net3402 _03430_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19559_ net3375 _03141_ net1881 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21521_ clknet_leaf_0_i_clk net1747 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21452_ clknet_leaf_39_i_clk net2100 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21383_ clknet_leaf_6_i_clk net5226 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20265_ net4128 net4097 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3110 net7929 vssd1 vssd1 vccd1 vccd1 net3637 sky130_fd_sc_hd__clkbuf_2
Xhold3121 net7608 vssd1 vssd1 vccd1 vccd1 net3648 sky130_fd_sc_hd__dlymetal6s2s_1
X_22004_ net446 net2637 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold3132 _00891_ vssd1 vssd1 vccd1 vccd1 net3659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20196_ net3509 net2125 _03709_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
Xhold3143 net7732 vssd1 vssd1 vccd1 vccd1 net3670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3154 _01237_ vssd1 vssd1 vccd1 vccd1 net3681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2420 net2303 vssd1 vssd1 vccd1 vccd1 net2947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3165 _03719_ vssd1 vssd1 vccd1 vccd1 net3692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2431 _00656_ vssd1 vssd1 vccd1 vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3176 net7684 vssd1 vssd1 vccd1 vccd1 net3703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2442 net5723 vssd1 vssd1 vccd1 vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3187 _01215_ vssd1 vssd1 vccd1 vccd1 net3714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2453 _01290_ vssd1 vssd1 vccd1 vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3198 net7858 vssd1 vssd1 vccd1 vccd1 net3725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2464 net5719 vssd1 vssd1 vccd1 vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03852_ clknet_0__03852_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03852_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1730 _03368_ vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2475 net7394 vssd1 vssd1 vccd1 vccd1 net3002 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2486 net4684 vssd1 vssd1 vccd1 vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1741 net6861 vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1752 net6972 vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19749__31 clknet_1_0__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2497 _01109_ vssd1 vssd1 vccd1 vccd1 net3024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1763 _01452_ vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1774 net7317 vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ net7437 net7234 _04276_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__mux2_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1785 _03516_ vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__buf_4
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1796 _00906_ vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ net7353 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__clkbuf_1
X_19764__45 clknet_1_1__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XFILLER_0_195_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ _06731_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__and2b_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ net6721 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ net41 _05700_ _05701_ net51 vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a22o_1
X_21719_ clknet_leaf_109_i_clk net4516 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _08325_ _08334_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__xor2_4
XFILLER_0_125_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ _05633_ net4156 vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_61_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ _04503_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__nand2_1
X_15171_ _06120_ _08260_ _08265_ vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__o21ai_4
X_12383_ _05517_ _05565_ _05567_ _05465_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ _07287_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__xnor2_1
X_11334_ rbzero.texu_hot\[1\] _04522_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14053_ _07177_ _07201_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a21oi_1
X_18930_ net1647 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_76_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11265_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__buf_4
Xhold5090 rbzero.wall_tracer.mapY\[9\] vssd1 vssd1 vccd1 vccd1 net5617 sky130_fd_sc_hd__dlygate4sd3_1
X_13004_ _06179_ net3847 vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nor2_1
X_18861_ net7421 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
X_11196_ net2745 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17812_ _02049_ _02050_ _08103_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_206_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _02925_ _02929_ net8246 _04482_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17743_ _08465_ _09354_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__nand2_1
X_14955_ net4383 _07947_ _08068_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _07045_ _07046_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__or2_1
X_17674_ _01893_ _01894_ _01913_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a21o_1
X_14886_ _06163_ _06235_ _06237_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_187_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19413_ net5356 _03310_ _03311_ _03312_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__a211o_1
X_13837_ _06966_ _06965_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__or2b_1
X_16625_ _09586_ _09714_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__and2_1
XFILLER_0_203_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap91 _09787_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16556_ _09644_ _09645_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19344_ net6552 _03271_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13768_ _06937_ _06938_ _06935_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15507_ _08599_ _08601_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__xor2_2
X_12719_ _05849_ _05871_ _05880_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a211o_2
X_19275_ net5037 _03200_ _03231_ _03230_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__o211a_1
X_16487_ net8225 net7771 _08111_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__mux2_1
X_13699_ _06868_ _06867_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_183_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7409 net4517 vssd1 vssd1 vccd1 vccd1 net7936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20668__14 clknet_1_0__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
X_15438_ net8267 _08129_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__nand2_1
X_18226_ net3820 net4537 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_i_clk clknet_4_11__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6708 rbzero.tex_r1\[56\] vssd1 vssd1 vccd1 vccd1 net7235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6719 net2573 vssd1 vssd1 vccd1 vccd1 net7246 sky130_fd_sc_hd__dlygate4sd3_1
X_15369_ _08463_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__buf_2
X_18157_ _02380_ _02381_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17108_ _10017_ _10018_ _10127_ vssd1 vssd1 vccd1 vccd1 _10129_ sky130_fd_sc_hd__and3_1
Xclkbuf_0__03846_ _03846_ vssd1 vssd1 vccd1 vccd1 clknet_0__03846_ sky130_fd_sc_hd__clkbuf_16
Xhold304 net5405 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18088_ net4518 net4351 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__or2_1
Xhold315 net5088 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold326 net5229 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 net8195 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold348 net5317 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
X_17039_ _09956_ _09961_ vssd1 vssd1 vccd1 vccd1 _10060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold359 net6064 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20050_ _03352_ net7607 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__nor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _01535_ vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _03416_ vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1026 _03466_ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1037 net6009 vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 _00651_ vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 net4272 vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ clknet_leaf_58_i_clk _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _02759_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21504_ clknet_leaf_14_i_clk net1312 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21435_ clknet_leaf_40_i_clk net1673 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21366_ clknet_leaf_20_i_clk net5306 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_20685__6 clknet_1_0__leaf__03506_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_0_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20317_ net6496 net3556 _03825_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 net6177 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_21297_ clknet_leaf_16_i_clk net5055 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold871 _00573_ vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 net6525 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net6219 net7099 _04342_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__mux2_1
X_20348__105 clknet_1_1__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__inv_2
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold893 net6391 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
X_20248_ net5206 _04648_ _04027_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__and3_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20179_ _03728_ net3928 vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or2_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 net7217 vssd1 vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2261 _01531_ vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2272 _01564_ vssd1 vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2283 net2906 vssd1 vssd1 vccd1 vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 net7263 vssd1 vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1560 _01421_ vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1571 net1365 vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ net7843 _07881_ _07882_ _07907_ net7812 vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__o311a_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ rbzero.debug_overlay.facingX\[-8\] _05113_ _05137_ _05140_ vssd1 vssd1 vccd1
+ vccd1 _05141_ sky130_fd_sc_hd__a211o_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1582 _01298_ vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 net6690 vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_106 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_106/HI o_rgb[17]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_117 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_117/HI zeros[6] sky130_fd_sc_hd__conb_1
X_10903_ net7033 net6164 _04265_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__mux2_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_128 vssd1 vssd1 vccd1 vccd1 ones[1] top_ew_algofoogle_128/LO sky130_fd_sc_hd__conb_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _07821_ _07830_ _07839_ _07841_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__a211o_1
Xtop_ew_algofoogle_139 vssd1 vssd1 vccd1 vccd1 ones[12] top_ew_algofoogle_139/LO sky130_fd_sc_hd__conb_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11883_ _05071_ net3919 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__and2b_1
X_16410_ _09400_ _09391_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ _06769_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__inv_2
X_10834_ net7494 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17390_ _08115_ _08369_ _08371_ vssd1 vssd1 vccd1 vccd1 _10408_ sky130_fd_sc_hd__o21a_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16341_ _09430_ _09432_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13553_ _06618_ _06634_ net80 vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__a21o_4
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10765_ net7081 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__clkbuf_1
X_19060_ net7597 net3583 net3397 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
X_12504_ _05640_ _05653_ _05662_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a211o_2
X_16272_ _09228_ _09238_ _09236_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__o21a_1
X_13484_ _06547_ _06546_ _06644_ _06651_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_180_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10696_ net7518 net6834 _04160_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15223_ _08317_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18011_ _02247_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__clkbuf_1
X_12435_ _05618_ _05619_ _05035_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ _06007_ _06334_ _04510_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__mux2_1
X_12366_ _05549_ _05550_ _04949_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14105_ _07224_ _07274_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _04505_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__or2b_1
X_19962_ net1568 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15085_ _08172_ _08173_ net8422 _08179_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__o2bb2a_4
X_12297_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _04978_ vssd1 vssd1 vccd1 vccd1 _05483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ _07160_ _07206_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__nand2_1
X_18913_ net3196 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
X_11248_ net3006 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__clkbuf_1
X_19893_ net3299 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18844_ _02983_ net4063 _02984_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__and3b_1
X_11179_ net6158 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18775_ _02904_ _02910_ _02921_ _04489_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a31o_1
X_15987_ _09079_ _09080_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ _01869_ _01870_ _01867_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14938_ net8034 _08037_ _01633_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17657_ _01784_ _09040_ _01895_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__o21ai_1
X_14869_ _08022_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16608_ _09696_ _09697_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19327_ net839 _03251_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__or2_1
X_16539_ _09614_ _09628_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7206 net3670 vssd1 vssd1 vccd1 vccd1 net7733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7217 net3927 vssd1 vssd1 vccd1 vccd1 net7744 sky130_fd_sc_hd__dlymetal6s2s_1
X_19258_ net5169 _03216_ _03222_ _03219_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__o211a_1
Xhold7239 _09090_ vssd1 vssd1 vccd1 vccd1 net7766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6505 rbzero.tex_g0\[43\] vssd1 vssd1 vccd1 vccd1 net7032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18209_ net3803 net4440 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nand2_1
Xhold6516 net2965 vssd1 vssd1 vccd1 vccd1 net7043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6527 rbzero.tex_r1\[18\] vssd1 vssd1 vccd1 vccd1 net7054 sky130_fd_sc_hd__dlygate4sd3_1
X_19189_ net5324 _03168_ _03181_ _03176_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__o211a_1
Xhold6538 net2658 vssd1 vssd1 vccd1 vccd1 net7065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6549 _04377_ vssd1 vssd1 vccd1 vccd1 net7076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5804 net1389 vssd1 vssd1 vccd1 vccd1 net6331 sky130_fd_sc_hd__dlygate4sd3_1
X_21220_ clknet_leaf_119_i_clk net1537 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5815 _03460_ vssd1 vssd1 vccd1 vccd1 net6342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 net2078 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5826 net1512 vssd1 vssd1 vccd1 vccd1 net6353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 net4735 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 net4979 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5837 _02492_ vssd1 vssd1 vccd1 vccd1 net6364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5848 _03817_ vssd1 vssd1 vccd1 vccd1 net6375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 net6053 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5859 net1372 vssd1 vssd1 vccd1 vccd1 net6386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 net8341 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21151_ clknet_leaf_106_i_clk net4840 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold156 net7418 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold167 net4716 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
X_20102_ net4436 _03660_ net664 _03679_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__o211a_1
Xhold178 net4975 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 net4989 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
X_21082_ clknet_leaf_68_i_clk _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20033_ _03109_ net5908 net3992 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__or3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21984_ net426 net2795 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20935_ clknet_leaf_78_i_clk net4553 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20866_ _09739_ _02512_ _04004_ _02508_ net5033 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20797_ net1015 net5522 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ net2021 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7740 net8012 vssd1 vssd1 vccd1 vccd1 net8267 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ net6142 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__clkbuf_1
X_12220_ rbzero.tex_g1\[31\] rbzero.tex_g1\[30\] _04950_ vssd1 vssd1 vccd1 vccd1 _05407_
+ sky130_fd_sc_hd__mux2_1
Xhold7784 net2910 vssd1 vssd1 vccd1 vccd1 net8311 sky130_fd_sc_hd__dlygate4sd3_1
X_21418_ clknet_leaf_42_i_clk net1534 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7795 net3466 vssd1 vssd1 vccd1 vccd1 net8322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _05239_ vssd1 vssd1 vccd1 vccd1 _05339_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21349_ clknet_leaf_45_i_clk net5218 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11102_ _04029_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__clkbuf_4
X_12082_ rbzero.tex_r1\[53\] rbzero.tex_r1\[52\] _04913_ vssd1 vssd1 vccd1 vccd1 _05271_
+ sky130_fd_sc_hd__mux2_1
Xhold690 net5487 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_102_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11033_ net6442 net6764 _04331_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__mux2_1
X_15910_ _08229_ _08322_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16890_ _09910_ _09911_ vssd1 vssd1 vccd1 vccd1 _09912_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15841_ _08888_ _08935_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__nand2_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 net7201 vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2091 _01374_ vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _06031_ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__xnor2_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _08863_ _08865_ _08866_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__a21o_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12984_ _06056_ net4645 net4780 _04479_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__o31a_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1390 _00673_ vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
X_17511_ _01750_ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xnor2_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ net4351 _07892_ _07872_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ net3417 _05106_ _05114_ net3317 vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18491_ _02653_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__inv_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20402__154 clknet_1_0__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__inv_2
XFILLER_0_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17442_ _10211_ _10220_ _10346_ _08918_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__o22ai_1
X_14654_ _07808_ _07824_ _07809_ _07795_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _05055_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _06767_ _06775_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__xnor2_1
X_10817_ net6810 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__clkbuf_1
X_17373_ _10308_ _10388_ _10389_ vssd1 vssd1 vccd1 vccd1 _10391_ sky130_fd_sc_hd__and3_1
X_14585_ _07753_ _07755_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__nand2_1
X_11797_ _04976_ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19112_ net2038 _03125_ net5541 _03128_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__o211a_1
X_13536_ _06703_ _06706_ _06697_ _06695_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__or4_4
XFILLER_0_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16324_ _08024_ _09414_ net75 _08115_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__a31o_1
XFILLER_0_166_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10748_ net2518 net7262 _04182_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16255_ _08127_ _09345_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19043_ net3597 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__clkbuf_1
X_13467_ _06493_ _06608_ _06610_ _06568_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__a211o_1
X_10679_ net7129 net6989 _04149_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _08299_ _08300_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__and2_1
X_12418_ rbzero.tex_b1\[59\] rbzero.tex_b1\[58\] _05369_ vssd1 vssd1 vccd1 vccd1 _05603_
+ sky130_fd_sc_hd__mux2_1
X_16186_ _09277_ _09278_ vssd1 vssd1 vccd1 vccd1 _09279_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13398_ _06564_ _06567_ _06568_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__o21a_1
X_15137_ _08230_ _08231_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _04849_ _05499_ _05516_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3709 rbzero.wall_tracer.visualWallDist\[-5\] vssd1 vssd1 vccd1 vccd1 net4236
+ sky130_fd_sc_hd__buf_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03514_ clknet_0__03514_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03514_
+ sky130_fd_sc_hd__clkbuf_16
X_19945_ net7455 net6239 _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
X_15068_ _05997_ _06317_ net4180 vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14019_ _07188_ _07189_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__xor2_1
X_19876_ net1231 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
X_18827_ net5877 net5845 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__nand2_1
X_18758_ rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\] _02856_
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17709_ _01947_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__nand2_2
XFILLER_0_210_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18689_ _02837_ _02842_ _02526_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720_ net1048 net5404 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20377__131 clknet_1_1__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__inv_2
XFILLER_0_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7003 net3243 vssd1 vssd1 vccd1 vccd1 net7530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7014 rbzero.pov.spi_buffer\[11\] vssd1 vssd1 vccd1 vccd1 net7541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7025 net1059 vssd1 vssd1 vccd1 vccd1 net7552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7036 _05087_ vssd1 vssd1 vccd1 vccd1 net7563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6302 rbzero.tex_b0\[29\] vssd1 vssd1 vccd1 vccd1 net6829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7047 rbzero.wall_tracer.mapY\[5\] vssd1 vssd1 vccd1 vccd1 net7574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6313 net1845 vssd1 vssd1 vccd1 vccd1 net6840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7058 net1447 vssd1 vssd1 vccd1 vccd1 net7585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6324 _04432_ vssd1 vssd1 vccd1 vccd1 net6851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7069 rbzero.spi_registers.spi_buffer\[21\] vssd1 vssd1 vccd1 vccd1 net7596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6335 net2268 vssd1 vssd1 vccd1 vccd1 net6862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5601 net1017 vssd1 vssd1 vccd1 vccd1 net6128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6346 rbzero.tex_g0\[4\] vssd1 vssd1 vccd1 vccd1 net6873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6357 net2014 vssd1 vssd1 vccd1 vccd1 net6884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5612 rbzero.tex_r1\[50\] vssd1 vssd1 vccd1 vccd1 net6139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6368 _04333_ vssd1 vssd1 vccd1 vccd1 net6895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5623 net1506 vssd1 vssd1 vccd1 vccd1 net6150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6379 net2158 vssd1 vssd1 vccd1 vccd1 net6906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5634 _02506_ vssd1 vssd1 vccd1 vccd1 net6161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5645 net1072 vssd1 vssd1 vccd1 vccd1 net6172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4900 rbzero.wall_tracer.mapY\[8\] vssd1 vssd1 vccd1 vccd1 net5427 sky130_fd_sc_hd__dlygate4sd3_1
X_21203_ clknet_leaf_109_i_clk net2090 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4911 net1088 vssd1 vssd1 vccd1 vccd1 net5438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5656 rbzero.tex_b1\[16\] vssd1 vssd1 vccd1 vccd1 net6183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4922 net8182 vssd1 vssd1 vccd1 vccd1 net5449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5667 rbzero.tex_r1\[11\] vssd1 vssd1 vccd1 vccd1 net6194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5678 net1128 vssd1 vssd1 vccd1 vccd1 net6205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4933 net1136 vssd1 vssd1 vccd1 vccd1 net5460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5689 _04448_ vssd1 vssd1 vccd1 vccd1 net6216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4944 rbzero.wall_tracer.mapX\[8\] vssd1 vssd1 vccd1 vccd1 net5471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4955 net1229 vssd1 vssd1 vccd1 vccd1 net5482 sky130_fd_sc_hd__dlygate4sd3_1
X_21134_ clknet_leaf_31_i_clk net4001 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_1
Xhold4966 _01612_ vssd1 vssd1 vccd1 vccd1 net5493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4977 rbzero.map_overlay.i_mapdx\[4\] vssd1 vssd1 vccd1 vccd1 net5504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4988 _00898_ vssd1 vssd1 vccd1 vccd1 net5515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4999 net1640 vssd1 vssd1 vccd1 vccd1 net5526 sky130_fd_sc_hd__dlygate4sd3_1
X_21065_ clknet_leaf_60_i_clk _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_20016_ _03205_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__clkbuf_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ net409 net2010 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ net88 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__buf_4
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ clknet_leaf_73_i_clk _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ net340 net2237 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ net1209 _04829_ _04824_ net1255 _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o221a_1
XFILLER_0_194_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20849_ net4192 _09745_ _09746_ _09091_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a22o_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ net6908 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14370_ _07539_ _07540_ _07491_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__a21bo_2
X_11582_ net1086 net1851 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _06491_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__buf_6
XFILLER_0_80_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ net2720 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16040_ _08131_ _08142_ _08226_ _09133_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__or4b_1
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7570 net652 vssd1 vssd1 vccd1 vccd1 net8097 sky130_fd_sc_hd__dlygate4sd3_1
X_13252_ _06410_ _06418_ _06422_ _06385_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__a31o_1
X_10464_ net2298 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7581 _02606_ vssd1 vssd1 vccd1 vccd1 net8108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7592 rbzero.traced_texa\[1\] vssd1 vssd1 vccd1 vccd1 net8119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12203_ rbzero.tex_g1\[3\] rbzero.tex_g1\[2\] _04916_ vssd1 vssd1 vccd1 vccd1 _05390_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6880 net2367 vssd1 vssd1 vccd1 vccd1 net7407 sky130_fd_sc_hd__dlygate4sd3_1
X_13183_ _04491_ _06321_ _06323_ _06327_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a2111o_1
Xhold6891 rbzero.pov.ready_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net7418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _05320_ _05321_ _04915_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17991_ _02222_ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__nand2_1
X_19730_ net1253 _03489_ net3707 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a21o_1
X_16942_ _09537_ _09664_ vssd1 vssd1 vccd1 vccd1 _09964_ sky130_fd_sc_hd__nor2_1
X_12065_ _05204_ _05251_ _05253_ _05213_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ net6249 net7338 _04320_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19661_ _04102_ net4835 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__nor2_4
X_16873_ _09652_ _09634_ vssd1 vssd1 vccd1 vccd1 _09895_ sky130_fd_sc_hd__or2b_1
XFILLER_0_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18612_ net3575 net5925 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ _08918_ _08691_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__nor2_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ net6858 net3738 net1779 vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__mux2_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ net4055 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__clkbuf_1
X_19800__77 clknet_1_1__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
X_15755_ _08829_ _08848_ _08849_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__a21o_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ net3965 net3848 _06136_ _06142_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a31o_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net4058 _05067_ net4107 net3516 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__o22a_1
X_14706_ _07860_ _07830_ _07875_ net7811 vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18474_ _02559_ net4821 net8086 net3947 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a31o_1
X_15686_ _08767_ _08769_ _08772_ _08778_ _08780_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _06066_ _06070_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or3_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _09262_ _09170_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11849_ net7570 net7731 _05012_ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__o22a_2
X_14637_ _07440_ _07794_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _10269_ _10270_ _10374_ vssd1 vssd1 vccd1 vccd1 _10375_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14568_ _07737_ _07738_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16307_ _09397_ _09396_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__or2b_1
XFILLER_0_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13519_ _06640_ _06689_ _06547_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__mux2_1
X_17287_ _10304_ _10305_ vssd1 vssd1 vccd1 vccd1 _10306_ sky130_fd_sc_hd__nor2_1
X_14499_ _07641_ _07640_ _07633_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19026_ net4041 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
X_16238_ _09209_ net3420 _09212_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4207 _03753_ vssd1 vssd1 vccd1 vccd1 net4734 sky130_fd_sc_hd__dlygate4sd3_1
X_16169_ _08323_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__clkbuf_4
Xhold4218 _00416_ vssd1 vssd1 vccd1 vccd1 net4745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4229 net3934 vssd1 vssd1 vccd1 vccd1 net4756 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3506 net7711 vssd1 vssd1 vccd1 vccd1 net4033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3517 _06035_ vssd1 vssd1 vccd1 vccd1 net4044 sky130_fd_sc_hd__clkbuf_4
Xhold3528 net5938 vssd1 vssd1 vccd1 vccd1 net4055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3539 _05051_ vssd1 vssd1 vccd1 vccd1 net4066 sky130_fd_sc_hd__buf_4
Xhold2805 rbzero.spi_registers.new_other\[7\] vssd1 vssd1 vccd1 vccd1 net3332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2816 _03549_ vssd1 vssd1 vccd1 vccd1 net3343 sky130_fd_sc_hd__dlygate4sd3_1
X_19928_ net7367 net3052 _03572_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2827 net4926 vssd1 vssd1 vccd1 vccd1 net3354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2838 net4614 vssd1 vssd1 vccd1 vccd1 net3365 sky130_fd_sc_hd__buf_2
Xhold2849 _03400_ vssd1 vssd1 vccd1 vccd1 net3376 sky130_fd_sc_hd__dlygate4sd3_1
X_19859_ net3156 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21821_ net263 net2634 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21752_ clknet_leaf_99_i_clk net4712 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_20703_ net967 net5384 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21683_ clknet_leaf_114_i_clk net5889 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6110 net1827 vssd1 vssd1 vccd1 vccd1 net6637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6121 rbzero.pov.spi_buffer\[25\] vssd1 vssd1 vccd1 vccd1 net6648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6132 net1798 vssd1 vssd1 vccd1 vccd1 net6659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6143 _04130_ vssd1 vssd1 vccd1 vccd1 net6670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6154 net1862 vssd1 vssd1 vccd1 vccd1 net6681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6165 rbzero.pov.ready_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net6692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5420 _04462_ vssd1 vssd1 vccd1 vccd1 net5947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6176 net2091 vssd1 vssd1 vccd1 vccd1 net6703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5431 rbzero.trace_state\[0\] vssd1 vssd1 vccd1 vccd1 net5958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6187 rbzero.tex_r1\[19\] vssd1 vssd1 vccd1 vccd1 net6714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5442 _05013_ vssd1 vssd1 vccd1 vccd1 net5969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6198 net1783 vssd1 vssd1 vccd1 vccd1 net6725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5453 gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 net5980 sky130_fd_sc_hd__dlygate4sd3_1
X_20431__180 clknet_1_1__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__inv_2
Xhold5464 net590 vssd1 vssd1 vccd1 vccd1 net5991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4730 _00790_ vssd1 vssd1 vccd1 vccd1 net5257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5475 rbzero.spi_registers.new_sky\[3\] vssd1 vssd1 vccd1 vccd1 net6002 sky130_fd_sc_hd__dlygate4sd3_1
X_22166_ clknet_leaf_96_i_clk net4881 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4741 net801 vssd1 vssd1 vccd1 vccd1 net5268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5486 rbzero.spi_registers.new_sky\[1\] vssd1 vssd1 vccd1 vccd1 net6013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5497 net2232 vssd1 vssd1 vccd1 vccd1 net6024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4752 rbzero.pov.spi_counter\[0\] vssd1 vssd1 vccd1 vccd1 net5279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4763 net994 vssd1 vssd1 vccd1 vccd1 net5290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4774 _00843_ vssd1 vssd1 vccd1 vccd1 net5301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4785 net931 vssd1 vssd1 vccd1 vccd1 net5312 sky130_fd_sc_hd__dlygate4sd3_1
X_21117_ clknet_leaf_92_i_clk net4795 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22097_ net159 net2498 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4796 rbzero.spi_registers.texadd0\[9\] vssd1 vssd1 vccd1 vccd1 net5323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21048_ clknet_leaf_78_i_clk _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13870_ _07012_ _07011_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__and2_1
XFILLER_0_199_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12821_ _05963_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15540_ _08631_ _08634_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__nand2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _05904_ _05928_ net37 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__o21a_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ net2910 _04464_ _04465_ net3488 _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15471_ _08519_ _08507_ _08518_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__a21oi_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ net33 _05860_ _05850_ net30 vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__and4b_1
XFILLER_0_210_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _10226_ _10227_ _10228_ vssd1 vssd1 vccd1 vccd1 _10230_ sky130_fd_sc_hd__a21o_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _07590_ _07591_ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__a21bo_4
X_11634_ _04823_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__clkbuf_8
X_18190_ _02245_ _02410_ _02411_ _10258_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17141_ _10159_ _10160_ vssd1 vssd1 vccd1 vccd1 _10161_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14353_ _07242_ _07326_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__nor2_1
X_11565_ _04753_ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13304_ _06472_ _06450_ _06473_ _06474_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and4_1
X_17072_ _10091_ _10092_ vssd1 vssd1 vccd1 vccd1 _10093_ sky130_fd_sc_hd__or2b_1
X_20514__255 clknet_1_0__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__inv_2
XFILLER_0_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10516_ net5637 net5645 _04064_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_1
X_14284_ _07431_ _07429_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__xor2_1
XFILLER_0_165_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11496_ net5915 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__inv_2
X_16023_ _08611_ _09116_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__nor2_1
X_13235_ _06365_ _06405_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__xor2_2
X_10447_ net47 net48 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__xor2_4
XFILLER_0_62_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ _06265_ _06007_ _06336_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1
+ vccd1 _06337_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12117_ _05303_ _05304_ _05276_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__mux2_1
X_17974_ _02209_ _02210_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__and2_1
X_13097_ net4446 net4828 vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__or2_1
X_19713_ _03122_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__nand2_2
X_12048_ _04916_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__clkbuf_8
X_16925_ _09945_ _09946_ vssd1 vssd1 vccd1 vccd1 _09947_ sky130_fd_sc_hd__xnor2_1
X_19644_ net6522 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__clkbuf_1
X_16856_ _09877_ _09876_ _09875_ _09868_ vssd1 vssd1 vccd1 vccd1 _09879_ sky130_fd_sc_hd__o211a_1
X_15807_ _08900_ _08901_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19575_ net2206 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
X_16787_ _09813_ _09816_ vssd1 vssd1 vccd1 vccd1 _09817_ sky130_fd_sc_hd__nor2_1
X_20595__327 clknet_1_0__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__inv_2
XFILLER_0_137_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13999_ _07168_ _07169_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__and2_1
X_18526_ _02687_ _02691_ net8260 _04482_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15738_ _08814_ _08817_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _02635_ _02636_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__or2_1
X_15669_ _08745_ _08746_ _08748_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17408_ _10333_ _10394_ _10424_ vssd1 vssd1 vccd1 vccd1 _10426_ sky130_fd_sc_hd__nand3_1
X_18388_ net3661 _02549_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17339_ _10355_ _10356_ vssd1 vssd1 vccd1 vccd1 _10358_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20350_ clknet_1_0__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__buf_1
XFILLER_0_109_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20489__232 clknet_1_1__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__inv_2
XFILLER_0_144_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19009_ net5786 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4004 _02766_ vssd1 vssd1 vccd1 vccd1 net4531 sky130_fd_sc_hd__dlygate4sd3_1
X_20281_ net3996 _03810_ _03812_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a21boi_1
X_22020_ net462 net1519 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
Xhold4026 net3393 vssd1 vssd1 vccd1 vccd1 net4553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4037 net7951 vssd1 vssd1 vccd1 vccd1 net4564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4048 net3791 vssd1 vssd1 vccd1 vccd1 net4575 sky130_fd_sc_hd__clkbuf_2
Xhold3303 net8337 vssd1 vssd1 vccd1 vccd1 net3830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3314 net8405 vssd1 vssd1 vccd1 vccd1 net3841 sky130_fd_sc_hd__buf_1
Xhold4059 _00424_ vssd1 vssd1 vccd1 vccd1 net4586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3325 net5896 vssd1 vssd1 vccd1 vccd1 net3852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3336 net2644 vssd1 vssd1 vccd1 vccd1 net3863 sky130_fd_sc_hd__buf_2
Xhold2602 _04049_ vssd1 vssd1 vccd1 vccd1 net3129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3347 net5584 vssd1 vssd1 vccd1 vccd1 net3874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 _01132_ vssd1 vssd1 vccd1 vccd1 net3140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3358 net7632 vssd1 vssd1 vccd1 vccd1 net3885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3369 rbzero.spi_registers.spi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net3896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2624 net4304 vssd1 vssd1 vccd1 vccd1 net3151 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2635 rbzero.tex_b1\[58\] vssd1 vssd1 vccd1 vccd1 net3162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1901 _00700_ vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
X_20663__9 clknet_1_1__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
Xhold2646 net2179 vssd1 vssd1 vccd1 vccd1 net3173 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1912 net7329 vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 _00669_ vssd1 vssd1 vccd1 vccd1 net3184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1923 net7207 vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 net3148 vssd1 vssd1 vccd1 vccd1 net3195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 _01439_ vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 net4578 vssd1 vssd1 vccd1 vccd1 net3206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1945 _04209_ vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1956 _04293_ vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1967 net5691 vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__buf_1
Xhold1978 _01405_ vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 _04219_ vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21804_ net246 net2885 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21735_ clknet_leaf_96_i_clk net4504 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21666_ clknet_leaf_122_i_clk net3011 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21597_ net231 net2084 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11350_ _04513_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ net4863 vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__clkbuf_2
X_13020_ _06194_ net4575 _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__o21ba_1
Xhold5250 net3464 vssd1 vssd1 vccd1 vccd1 net5777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5261 net584 vssd1 vssd1 vccd1 vccd1 net5788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5272 net1250 vssd1 vssd1 vccd1 vccd1 net5799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5283 _00626_ vssd1 vssd1 vccd1 vccd1 net5810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4560 net696 vssd1 vssd1 vccd1 vccd1 net5087 sky130_fd_sc_hd__dlygate4sd3_1
X_22149_ clknet_leaf_51_i_clk _01636_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4571 _00811_ vssd1 vssd1 vccd1 vccd1 net5098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4582 net797 vssd1 vssd1 vccd1 vccd1 net5109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4593 rbzero.spi_registers.texadd0\[14\] vssd1 vssd1 vccd1 vccd1 net5120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3870 net3467 vssd1 vssd1 vccd1 vccd1 net4397 sky130_fd_sc_hd__dlymetal6s2s_1
X_14971_ _08083_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__clkbuf_1
Xhold3892 net877 vssd1 vssd1 vccd1 vccd1 net4419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16710_ _04566_ net7609 _09747_ vssd1 vssd1 vccd1 vccd1 _09749_ sky130_fd_sc_hd__mux2_1
X_13922_ _06996_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__xor2_2
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17690_ _01917_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ net3919 net4124 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__nor2_1
X_13853_ _07004_ _07022_ _07023_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ _05948_ _05976_ _05977_ _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__a311o_4
X_19360_ net5105 _03269_ _03281_ _03275_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__o211a_1
X_16572_ _09656_ _09661_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__xor2_1
X_10996_ net2683 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
X_13784_ _06720_ _06953_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18311_ net6191 net3478 _02476_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15523_ _08615_ _08617_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__nor2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19291_ net1281 _03238_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__or2_1
X_12735_ net35 net34 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and2_2
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ net3926 net4608 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__nand2_1
X_15454_ _08127_ _08535_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nor2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12666_ _05830_ _05836_ _05844_ _05796_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a22o_2
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11617_ net3189 _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14405_ _07242_ _07391_ _07571_ _07575_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__o31a_1
X_18173_ _02395_ _02396_ net3666 _02390_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a211o_1
X_15385_ _08377_ _08387_ _08385_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__a21bo_1
X_12597_ _04020_ _04495_ net7678 _04500_ net16 _05747_ vssd1 vssd1 vccd1 vccd1 _05777_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17124_ _10055_ _10141_ _10143_ vssd1 vssd1 vccd1 vccd1 _10144_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03862_ _03862_ vssd1 vssd1 vccd1 vccd1 clknet_0__03862_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14336_ _07383_ _07433_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ net4369 vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold508 net4313 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _10072_ _10074_ vssd1 vssd1 vccd1 vccd1 _10076_ sky130_fd_sc_hd__nand2_1
Xhold519 net5447 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ _07347_ _07363_ _07361_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ net4138 _04661_ _04662_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _09099_ _09100_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__nand2_1
X_13218_ _06386_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _07355_ _07367_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__or2_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _06278_ _06291_ _06289_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_209_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17957_ _02192_ _02193_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__or2b_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _00904_ vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 net6630 vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
X_16908_ _09894_ _09929_ vssd1 vssd1 vccd1 vccd1 _09930_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17888_ _02124_ _02125_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19627_ net1669 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
X_16839_ _09818_ _09450_ vssd1 vssd1 vccd1 vccd1 _09864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19558_ net1883 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18509_ _02666_ _02672_ _02683_ _04489_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a31o_1
X_19489_ net4016 net6024 _03354_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21520_ clknet_leaf_0_i_clk net1699 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21451_ clknet_leaf_36_i_clk net1404 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21382_ clknet_leaf_9_i_clk net5103 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20264_ _05673_ net3970 _03801_ _03765_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3100 net5959 vssd1 vssd1 vccd1 vccd1 net3627 sky130_fd_sc_hd__dlygate4sd3_1
X_22003_ net445 net2034 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold3122 net7610 vssd1 vssd1 vccd1 vccd1 net3649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3133 net8254 vssd1 vssd1 vccd1 vccd1 net3660 sky130_fd_sc_hd__dlygate4sd3_1
X_20195_ net3663 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
Xhold3144 _03317_ vssd1 vssd1 vccd1 vccd1 net3671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2410 net7343 vssd1 vssd1 vccd1 vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3155 net7704 vssd1 vssd1 vccd1 vccd1 net3682 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2421 _04106_ vssd1 vssd1 vccd1 vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3166 _01202_ vssd1 vssd1 vccd1 vccd1 net3693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 net7402 vssd1 vssd1 vccd1 vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3177 _03490_ vssd1 vssd1 vccd1 vccd1 net3704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2443 net7000 vssd1 vssd1 vccd1 vccd1 net2970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03851_ clknet_0__03851_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03851_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2454 net7086 vssd1 vssd1 vccd1 vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1720 net7008 vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3199 net7875 vssd1 vssd1 vccd1 vccd1 net3726 sky130_fd_sc_hd__buf_1
Xhold2465 _01326_ vssd1 vssd1 vccd1 vccd1 net2992 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1731 _00920_ vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2476 _03407_ vssd1 vssd1 vccd1 vccd1 net3003 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1742 net6863 vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2487 net4511 vssd1 vssd1 vccd1 vccd1 net3014 sky130_fd_sc_hd__buf_2
Xhold1753 _04394_ vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2498 rbzero.pov.spi_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net3025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1764 net7144 vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20543__281 clknet_1_1__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__inv_2
XFILLER_0_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1775 _01365_ vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1786 _03595_ vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1797 net6966 vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ net7351 net2595 _04238_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10781_ net2569 net6719 _04205_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ net11 _05691_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21718_ clknet_leaf_109_i_clk net3722 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ net4 vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__clkbuf_4
X_21649_ clknet_leaf_126_i_clk net3229 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ _04558_ _04559_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__nand2_1
X_15170_ net3457 _08194_ _08264_ _08137_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__a211o_1
X_12382_ _04922_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_90 net4293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14121_ _07290_ _07291_ _07258_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ rbzero.texu_hot\[0\] _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _07221_ _07222_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__xnor2_1
X_11264_ net5911 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5080 net2278 vssd1 vssd1 vccd1 vccd1 net5607 sky130_fd_sc_hd__dlygate4sd3_1
X_13003_ net4547 vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5091 net2058 vssd1 vssd1 vccd1 vccd1 net5618 sky130_fd_sc_hd__dlygate4sd3_1
X_18860_ net2764 net7419 _02993_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__mux2_1
X_11195_ net7270 net6987 _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17811_ _01949_ _01951_ _01947_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__o21a_1
Xhold4390 net4694 vssd1 vssd1 vccd1 vccd1 net4917 sky130_fd_sc_hd__clkbuf_4
X_20626__356 clknet_1_0__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__inv_2
XFILLER_0_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ net4709 net4560 _02929_ _02866_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _01979_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__xor2_1
X_14954_ _08074_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _07047_ _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__or2_1
X_17673_ _01902_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__xnor2_1
X_14885_ _06239_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19412_ _04459_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__buf_6
X_16624_ _09711_ net4190 vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__xnor2_1
X_13836_ _06968_ _06969_ _06973_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap81 _06539_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap92 _04028_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_4
X_19343_ net5017 _03269_ _03272_ _03259_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__o211a_1
X_16555_ _09511_ _09512_ _09509_ vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__a21boi_1
X_10979_ net7013 net6655 _04309_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__mux2_1
X_13767_ _06719_ _06715_ _06725_ _06793_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_169_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15506_ _08539_ _08600_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19274_ net2414 _03202_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__or2_1
X_12718_ _05883_ _05885_ _05889_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a31o_1
X_16486_ _09460_ _09576_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__xnor2_4
X_13698_ _06727_ _06725_ _06726_ _06768_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__a22o_1
X_18225_ net3820 net4537 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__nor2_1
X_15437_ _08530_ _08531_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__or2b_1
XFILLER_0_183_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ _05810_ _05816_ _05821_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6709 net2851 vssd1 vssd1 vccd1 vccd1 net7236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20371__126 clknet_1_0__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__inv_2
XFILLER_0_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _02372_ _02373_ _02374_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__o21ai_2
X_15368_ _06119_ net4877 vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17107_ _10017_ _10018_ _10127_ vssd1 vssd1 vccd1 vccd1 _10128_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03845_ _03845_ vssd1 vssd1 vccd1 vccd1 clknet_0__03845_ sky130_fd_sc_hd__clkbuf_16
Xhold305 net5327 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ _07489_ _07305_ _07342_ _06931_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18087_ _02321_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__clkbuf_1
Xhold316 net5090 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ _08390_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold327 net5379 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold338 net8001 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17038_ _09940_ _09950_ _09948_ vssd1 vssd1 vccd1 vccd1 _10059_ sky130_fd_sc_hd__a21o_1
Xhold349 net7564 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ net1472 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 net6013 vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _00957_ vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _00998_ vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 net6011 vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 net6495 vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20951_ clknet_leaf_58_i_clk _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20882_ _02751_ net4529 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__and2b_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21503_ clknet_leaf_13_i_clk net1309 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21434_ clknet_leaf_40_i_clk net1636 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21365_ clknet_leaf_20_i_clk net5071 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20316_ net6572 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21296_ clknet_leaf_16_i_clk net5095 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold850 net6284 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _01277_ vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 net6135 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold883 _01312_ vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_20247_ _04648_ _04026_ _05184_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__nand3_1
Xhold894 _00577_ vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ net7744 net3276 _03723_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__mux2_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2240 net2879 vssd1 vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2251 _04344_ vssd1 vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2262 rbzero.tex_r1\[37\] vssd1 vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2273 rbzero.pov.spi_buffer\[48\] vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2284 _04177_ vssd1 vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2295 _01457_ vssd1 vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 _01010_ vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1561 net2973 vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1572 _03392_ vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
X_11951_ rbzero.debug_overlay.facingX\[-3\] _05095_ _05138_ _05139_ vssd1 vssd1 vccd1
+ vccd1 _05140_ sky130_fd_sc_hd__a211o_1
Xhold1583 net6710 vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1594 _01588_ vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_107 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_107/HI o_rgb[18]
+ sky130_fd_sc_hd__conb_1
X_10902_ net2236 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_118 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_118/HI zeros[7] sky130_fd_sc_hd__conb_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _04668_ net4121 _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__or3_1
X_14670_ net7843 vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__buf_2
Xtop_ew_algofoogle_129 vssd1 vssd1 vccd1 vccd1 ones[2] top_ew_algofoogle_129/LO sky130_fd_sc_hd__conb_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10833_ net2848 net7492 _04227_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13621_ _06759_ _06756_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _09285_ _09306_ _09431_ vssd1 vssd1 vccd1 vccd1 _09432_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10764_ net2376 net7079 _04194_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
X_13552_ net80 _06634_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12503_ _05664_ _05667_ _05671_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a31o_1
X_16271_ _09350_ _09362_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13483_ _06568_ _06653_ net559 vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__o21a_1
X_10695_ net6154 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18010_ _02246_ net4762 _10260_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_2
XFILLER_0_180_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ _05031_ _05026_ net4080 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__o21a_1
X_15222_ net4353 _08162_ _08315_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_125_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12365_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _05250_ vssd1 vssd1 vccd1 vccd1 _05550_
+ sky130_fd_sc_hd__mux2_1
X_15153_ _08242_ _08247_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__nand2_2
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14104_ _07224_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__nand2_1
X_11316_ rbzero.spi_registers.texadd3\[13\] rbzero.spi_registers.texadd1\[13\] _04504_
+ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__mux2_1
X_19961_ net3009 net5988 _03583_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15084_ net3315 _06033_ _08123_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__o211a_1
X_12296_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _05220_ vssd1 vssd1 vccd1 vccd1 _05482_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ _07204_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__and2_1
X_18912_ net3195 net7552 _03014_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__mux2_1
X_11247_ net7413 net7023 _04445_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19892_ net3273 net3298 _03550_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__mux2_1
X_18843_ _02947_ _02979_ net3485 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a21o_1
X_11178_ net6156 net1929 _04412_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__mux2_1
X_18774_ _02904_ _02910_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a21oi_1
X_15986_ _09079_ _09080_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17725_ _01890_ _01858_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__or2b_1
X_14937_ _04481_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17656_ _01784_ _09040_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__or3_1
X_14868_ net4428 _08021_ _07976_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16607_ _09522_ _09563_ _09562_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13819_ net3526 net566 _06989_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__a21boi_4
X_17587_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14799_ _07844_ _07847_ _07931_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__a31o_2
X_19326_ net5133 _03250_ _03261_ _03259_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__o211a_1
X_16538_ _09626_ _09627_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7207 _05381_ vssd1 vssd1 vccd1 vccd1 net7734 sky130_fd_sc_hd__dlygate4sd3_1
X_19257_ net6484 _03217_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ _09426_ _09428_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__and2b_1
Xhold7218 rbzero.spi_registers.got_new_vshift vssd1 vssd1 vccd1 vccd1 net7745 sky130_fd_sc_hd__dlygate4sd3_1
X_18208_ net3803 net4440 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6506 net2453 vssd1 vssd1 vccd1 vccd1 net7033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6517 rbzero.pov.ready_buffer\[16\] vssd1 vssd1 vccd1 vccd1 net7044 sky130_fd_sc_hd__dlygate4sd3_1
X_19188_ net6566 _03170_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__or2_1
Xhold6528 net2641 vssd1 vssd1 vccd1 vccd1 net7055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6539 rbzero.tex_r0\[56\] vssd1 vssd1 vccd1 vccd1 net7066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5805 _02507_ vssd1 vssd1 vccd1 vccd1 net6332 sky130_fd_sc_hd__dlygate4sd3_1
X_18139_ net3768 net4392 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__nand2_1
Xhold5816 net1338 vssd1 vssd1 vccd1 vccd1 net6343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold102 net4503 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5827 rbzero.spi_registers.new_texadd\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net6354
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 net4967 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5838 net1515 vssd1 vssd1 vccd1 vccd1 net6365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net4981 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5849 net1369 vssd1 vssd1 vccd1 vccd1 net6376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _01283_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ clknet_leaf_104_i_clk net3603 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold146 net4322 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 net4637 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ net663 _03610_ _03661_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a211o_1
Xhold168 net5084 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold179 net4977 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21081_ clknet_leaf_68_i_clk _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20609__340 clknet_1_0__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__inv_2
XFILLER_0_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20032_ _03606_ _03635_ net3991 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19806__83 clknet_1_0__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__inv_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21983_ net425 net1796 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ clknet_leaf_78_i_clk net4732 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20865_ net3565 net5033 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__or2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_75_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20796_ _03959_ _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20655__382 clknet_1_1__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__inv_2
XFILLER_0_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20354__110 clknet_1_1__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__inv_2
Xhold7730 _02666_ vssd1 vssd1 vccd1 vccd1 net8257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ net2438 net6140 _04042_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__mux2_1
Xhold7741 rbzero.debug_overlay.vplaneX\[-6\] vssd1 vssd1 vccd1 vccd1 net8268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7774 rbzero.traced_texVinit\[9\] vssd1 vssd1 vccd1 vccd1 net8301 sky130_fd_sc_hd__dlygate4sd3_1
X_21417_ clknet_leaf_41_i_clk net1735 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7785 rbzero.row_render.size\[9\] vssd1 vssd1 vccd1 vccd1 net8312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7796 rbzero.wall_tracer.stepDistY\[-7\] vssd1 vssd1 vccd1 vccd1 net8323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _04913_ vssd1 vssd1 vccd1 vccd1 _05338_
+ sky130_fd_sc_hd__mux2_1
X_21348_ clknet_leaf_45_i_clk net5203 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11101_ net2979 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_13_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12081_ _04984_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 net6278 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
X_21279_ clknet_leaf_25_i_clk net4453 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold691 net5489 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net6120 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15840_ _08925_ _08930_ _08929_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__a21bo_1
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 _01409_ vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2081 _04430_ vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 net6988 vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _08864_ _08253_ _08464_ _08573_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__and4_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net4779 _06146_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a21oi_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _09612_ _09373_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__and2b_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1380 _03045_ vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1391 net5608 vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ net7833 _07880_ _07891_ _07869_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__a31o_2
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _02626_ net3614 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__or2_1
X_11934_ net3489 _05113_ _05090_ net3315 _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _08918_ _10211_ _10220_ _10346_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__or4_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ net8355 _07823_ _07439_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ reg_rgb\[6\] _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__mux2_4
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13604_ _06770_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17372_ _10308_ _10388_ _10389_ vssd1 vssd1 vccd1 vccd1 _10390_ sky130_fd_sc_hd__a21oi_2
X_10816_ net2638 net6808 _04216_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _04978_ vssd1 vssd1 vccd1 vccd1 _04986_
+ sky130_fd_sc_hd__mux2_1
X_14584_ _07752_ _07754_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19111_ net5540 _03126_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16323_ _08024_ net75 _09414_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10747_ net3000 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19042_ net3596 net3562 net3398 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
X_16254_ _08127_ _09225_ _09345_ _08611_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ net2636 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__clkbuf_1
X_13466_ _06635_ _06636_ _06606_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15205_ net3445 _08256_ net4284 vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _05517_ _05599_ _05601_ _05233_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16185_ _08509_ _08418_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13397_ _06516_ _06539_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nand2_2
XFILLER_0_51_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15136_ net4344 _08188_ net3317 vssd1 vssd1 vccd1 vccd1 _08231_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ _05263_ _05521_ _05525_ _05533_ _04818_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03513_ clknet_0__03513_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03513_
+ sky130_fd_sc_hd__clkbuf_16
X_12279_ _04947_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__clkbuf_8
X_15067_ _08137_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__buf_4
X_19944_ net2311 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14018_ _07137_ _07139_ _07141_ _07098_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__a22o_1
X_19875_ net6357 net3195 _03539_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__mux2_1
X_18826_ net5845 _02968_ net4063 net2199 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__o211a_1
X_18757_ _02892_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__inv_2
X_15969_ _08127_ _08614_ _09062_ _08611_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17708_ _01944_ _01946_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18688_ _02826_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17639_ _01873_ _01788_ _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19309_ net5260 _03250_ _03252_ _03246_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7004 rbzero.tex_g0\[30\] vssd1 vssd1 vccd1 vccd1 net7531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7015 net2869 vssd1 vssd1 vccd1 vccd1 net7542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7026 rbzero.pov.spi_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net7553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7037 rbzero.pov.ready_buffer\[30\] vssd1 vssd1 vccd1 vccd1 net7564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6303 net1897 vssd1 vssd1 vccd1 vccd1 net6830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7048 net3447 vssd1 vssd1 vccd1 vccd1 net7575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6314 _04146_ vssd1 vssd1 vccd1 vccd1 net6841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7059 rbzero.pov.ready_buffer\[63\] vssd1 vssd1 vccd1 vccd1 net7586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6325 net1759 vssd1 vssd1 vccd1 vccd1 net6852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6336 _03449_ vssd1 vssd1 vccd1 vccd1 net6863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5602 _04360_ vssd1 vssd1 vccd1 vccd1 net6129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6347 net2116 vssd1 vssd1 vccd1 vccd1 net6874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5613 net1040 vssd1 vssd1 vccd1 vccd1 net6140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6358 _04262_ vssd1 vssd1 vccd1 vccd1 net6885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6369 net2064 vssd1 vssd1 vccd1 vccd1 net6896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5624 rbzero.tex_r0\[14\] vssd1 vssd1 vccd1 vccd1 net6151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21202_ clknet_leaf_109_i_clk net2332 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5635 net1600 vssd1 vssd1 vccd1 vccd1 net6162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5646 _04128_ vssd1 vssd1 vccd1 vccd1 net6173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4901 net1006 vssd1 vssd1 vccd1 vccd1 net5428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5657 net1069 vssd1 vssd1 vccd1 vccd1 net6184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4912 rbzero.floor_leak\[0\] vssd1 vssd1 vccd1 vccd1 net5439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4923 net1047 vssd1 vssd1 vccd1 vccd1 net5450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5668 net1115 vssd1 vssd1 vccd1 vccd1 net6195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4934 _00880_ vssd1 vssd1 vccd1 vccd1 net5461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5679 rbzero.spi_registers.new_texadd\[1\]\[23\] vssd1 vssd1 vccd1 vccd1 net6206
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21133_ clknet_leaf_29_i_clk net5920 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_1
Xhold4945 net1161 vssd1 vssd1 vccd1 vccd1 net5472 sky130_fd_sc_hd__buf_1
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4956 rbzero.floor_leak\[2\] vssd1 vssd1 vccd1 vccd1 net5483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4967 net1234 vssd1 vssd1 vccd1 vccd1 net5494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4978 net3982 vssd1 vssd1 vccd1 vccd1 net5505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4989 net1659 vssd1 vssd1 vccd1 vccd1 net5516 sky130_fd_sc_hd__dlygate4sd3_1
X_21064_ clknet_leaf_64_i_clk _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20015_ _03608_ net5850 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21966_ net408 net1129 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ clknet_leaf_74_i_clk _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ net339 net2455 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ net1050 _04833_ _04838_ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a31o_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ net5657 net63 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__nor2_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ net6906 net2201 _04105_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__mux2_1
X_11581_ _04768_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nand2_1
X_20779_ _03943_ _03947_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ net7192 net2719 _04064_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__buf_6
XFILLER_0_165_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7560 _00606_ vssd1 vssd1 vccd1 vccd1 net8087 sky130_fd_sc_hd__dlygate4sd3_1
X_10463_ net6836 net6888 _04031_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__mux2_1
Xhold7571 _01651_ vssd1 vssd1 vccd1 vccd1 net8098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13251_ _06420_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nor2_1
Xhold7582 net1609 vssd1 vssd1 vccd1 vccd1 net8109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7593 net948 vssd1 vssd1 vccd1 vccd1 net8120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12202_ _04943_ _05386_ _05388_ _04947_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6870 net3070 vssd1 vssd1 vccd1 vccd1 net7397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13182_ _04491_ _06329_ _06332_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__o211ai_2
X_20340__97 clknet_1_0__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__inv_2
Xhold6881 rbzero.pov.ready_buffer\[11\] vssd1 vssd1 vccd1 vccd1 net7408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6892 net683 vssd1 vssd1 vccd1 vccd1 net7419 sky130_fd_sc_hd__dlygate4sd3_1
X_12133_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _04933_ vssd1 vssd1 vccd1 vccd1 _05321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _02225_ _02226_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16941_ _09954_ _09962_ vssd1 vssd1 vccd1 vccd1 _09963_ sky130_fd_sc_hd__xor2_1
X_12064_ _04984_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
X_11015_ net7159 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19660_ net6323 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
X_16872_ _09614_ _09628_ _09626_ vssd1 vssd1 vccd1 vccd1 _09894_ sky130_fd_sc_hd__a21o_1
X_18611_ net4530 _02763_ _02764_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o21a_1
X_15823_ _08880_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__buf_4
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__05898_ clknet_0__05898_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05898_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19591_ net1656 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18542_ net4054 _06039_ _06242_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
X_15754_ _08830_ _08847_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__nor2_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _06137_ _06141_ net3999 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__a21oi_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _07818_ _07874_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__nor2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _02650_ _02651_ rbzero.wall_tracer.rayAddendX\[5\] _09735_ vssd1 vssd1 vccd1
+ vccd1 _02652_ sky130_fd_sc_hd__a2bb2o_1
X_11917_ _05088_ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__nor2_2
XFILLER_0_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15685_ _08779_ _08772_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__xnor2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ net3991 net4034 net3807 net3553 _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a221o_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _01664_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__xnor2_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _07240_ _07360_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__nor2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _05017_ _05037_ net7570 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a21bo_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _10144_ _10373_ vssd1 vssd1 vccd1 vccd1 _10374_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14567_ _07734_ _07736_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__or2_1
X_11779_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _04968_ vssd1 vssd1 vccd1 vccd1 _04969_
+ sky130_fd_sc_hd__mux2_1
X_16306_ _09396_ _09397_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ _06438_ _06447_ _06453_ _06450_ _06493_ _06571_ vssd1 vssd1 vccd1 vccd1 _06689_
+ sky130_fd_sc_hd__mux4_1
X_17286_ _10302_ _10303_ vssd1 vssd1 vccd1 vccd1 _10305_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498_ _07641_ _07633_ _07640_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ net4040 net2205 _03078_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__mux2_1
X_16237_ _09328_ _09329_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__nand2_1
X_13449_ _06551_ _06597_ _06598_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16168_ _09259_ _09260_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4208 _01221_ vssd1 vssd1 vccd1 vccd1 net4735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4219 net3355 vssd1 vssd1 vccd1 vccd1 net4746 sky130_fd_sc_hd__dlygate4sd3_1
X_15119_ net4344 _08188_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3507 _06071_ vssd1 vssd1 vccd1 vccd1 net4034 sky130_fd_sc_hd__clkbuf_4
X_16099_ _09189_ _09191_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__nand2_1
Xhold3518 net7637 vssd1 vssd1 vccd1 vccd1 net4045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3529 _00613_ vssd1 vssd1 vccd1 vccd1 net4056 sky130_fd_sc_hd__dlygate4sd3_1
X_19927_ net2412 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
Xhold2806 net3035 vssd1 vssd1 vccd1 vccd1 net3333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2817 _01115_ vssd1 vssd1 vccd1 vccd1 net3344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2828 net4745 vssd1 vssd1 vccd1 vccd1 net3355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2839 rbzero.spi_registers.new_other\[6\] vssd1 vssd1 vccd1 vccd1 net3366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19858_ net7498 net6125 _03528_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_1
X_18809_ net3770 net4832 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21820_ net262 net1890 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21751_ clknet_leaf_132_i_clk net4563 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20702_ net967 net5384 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21682_ clknet_leaf_113_i_clk net5839 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6100 net2613 vssd1 vssd1 vccd1 vccd1 net6627 sky130_fd_sc_hd__buf_1
Xhold6111 _04379_ vssd1 vssd1 vccd1 vccd1 net6638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6122 net1688 vssd1 vssd1 vccd1 vccd1 net6649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6133 rbzero.pov.spi_buffer\[5\] vssd1 vssd1 vccd1 vccd1 net6660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6144 net1849 vssd1 vssd1 vccd1 vccd1 net6671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6155 rbzero.spi_registers.new_texadd\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net6682
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5410 net4641 vssd1 vssd1 vccd1 vccd1 net5937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6166 net746 vssd1 vssd1 vccd1 vccd1 net6693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5421 _05185_ vssd1 vssd1 vccd1 vccd1 net5948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5432 net4861 vssd1 vssd1 vccd1 vccd1 net5959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6177 rbzero.tex_g0\[13\] vssd1 vssd1 vccd1 vccd1 net6704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6188 net1839 vssd1 vssd1 vccd1 vccd1 net6715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6199 rbzero.spi_registers.new_texadd\[0\]\[18\] vssd1 vssd1 vccd1 vccd1 net6726
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5454 net4023 vssd1 vssd1 vccd1 vccd1 net5981 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold5465 _04172_ vssd1 vssd1 vccd1 vccd1 net5992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4720 rbzero.spi_registers.texadd3\[21\] vssd1 vssd1 vccd1 vccd1 net5247 sky130_fd_sc_hd__dlygate4sd3_1
X_22165_ clknet_leaf_96_i_clk net4602 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4731 net923 vssd1 vssd1 vccd1 vccd1 net5258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5476 net1724 vssd1 vssd1 vccd1 vccd1 net6003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4742 _00834_ vssd1 vssd1 vccd1 vccd1 net5269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5487 net1532 vssd1 vssd1 vccd1 vccd1 net6014 sky130_fd_sc_hd__dlygate4sd3_1
X_20466__211 clknet_1_0__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__inv_2
XFILLER_0_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4753 net973 vssd1 vssd1 vccd1 vccd1 net5280 sky130_fd_sc_hd__buf_1
Xhold5498 rbzero.tex_b0\[60\] vssd1 vssd1 vccd1 vccd1 net6025 sky130_fd_sc_hd__dlygate4sd3_1
X_21116_ clknet_leaf_93_i_clk net3606 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4764 rbzero.spi_registers.texadd0\[11\] vssd1 vssd1 vccd1 vccd1 net5291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4775 net857 vssd1 vssd1 vccd1 vccd1 net5302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22096_ net158 net1042 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
Xhold4786 _00862_ vssd1 vssd1 vccd1 vccd1 net5313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4797 net962 vssd1 vssd1 vccd1 vccd1 net5324 sky130_fd_sc_hd__dlygate4sd3_1
X_21047_ clknet_leaf_58_i_clk _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ _05949_ _05956_ _05960_ _05967_ _05970_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__o41a_1
XFILLER_0_199_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _05680_ _05043_ _05730_ net3996 _05901_ net36 vssd1 vssd1 vccd1 vccd1 _05928_
+ sky130_fd_sc_hd__mux4_1
X_21949_ net391 net2568 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ net2910 _04463_ net3955 net3405 _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a221o_1
X_15470_ _08519_ _08507_ _08518_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__and3_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05856_ _05858_ _05859_ net32 vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _07072_ _06754_ _07304_ _07280_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__or4_4
X_11633_ _04802_ _04814_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__or3_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _08542_ net7818 vssd1 vssd1 vccd1 vccd1 _10160_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14352_ _07033_ _07197_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__or2_1
X_11564_ net941 net1918 vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ net570 _06406_ _06441_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__nor3_1
X_17071_ _10084_ _10085_ _10090_ vssd1 vssd1 vccd1 vccd1 _10092_ sky130_fd_sc_hd__or3_1
X_10515_ net2775 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__clkbuf_1
X_11495_ net3552 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__inv_2
X_14283_ _07434_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__xor2_2
X_16022_ _09115_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7390 net3475 vssd1 vssd1 vccd1 vccd1 net7917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13234_ _06404_ _06355_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__and2_1
X_10446_ _04023_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13165_ net4277 net8051 vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12116_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _05258_ vssd1 vssd1 vccd1 vccd1 _05304_
+ sky130_fd_sc_hd__mux2_1
X_17973_ _02203_ _02208_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__or2_1
X_13096_ net8265 _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16924_ _09262_ _08403_ vssd1 vssd1 vccd1 vccd1 _09946_ sky130_fd_sc_hd__nor2_1
X_12047_ _05234_ _05235_ _05206_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__mux2_1
X_19712_ net41 net40 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__or2_2
X_16855_ _09868_ _09875_ _09876_ _09877_ vssd1 vssd1 vccd1 vccd1 _09878_ sky130_fd_sc_hd__a211oi_2
X_19643_ net6520 net3592 _03441_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
X_15806_ _08417_ _08691_ _08899_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__o21bai_1
X_19574_ net7303 net2205 _03403_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
X_16786_ _09814_ _09815_ vssd1 vssd1 vccd1 vccd1 _09816_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13998_ _06673_ _06698_ _07167_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__o21ai_1
X_18525_ net4603 net4554 _02691_ _02627_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a211oi_1
X_15737_ _08778_ _08780_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ net3965 net4044 vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__xor2_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18456_ _02607_ _02633_ _02634_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15668_ _08725_ _08751_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _10333_ _10394_ _10424_ vssd1 vssd1 vccd1 vccd1 _10425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14619_ _07434_ _07453_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__and2_2
XFILLER_0_172_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18387_ net3661 net3565 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__nand2_1
X_15599_ _08692_ _08693_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__or2b_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17338_ _10355_ _10356_ vssd1 vssd1 vccd1 vccd1 _10357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17269_ net8035 _06124_ _09413_ vssd1 vssd1 vccd1 vccd1 _10288_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19008_ net1613 net5784 _02992_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20280_ _09733_ _03793_ _03810_ net3996 _09725_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o221a_1
Xhold4005 net8130 vssd1 vssd1 vccd1 vccd1 net4532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4016 net8190 vssd1 vssd1 vccd1 vccd1 net4543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4027 rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 net4554 sky130_fd_sc_hd__buf_2
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4038 net2877 vssd1 vssd1 vccd1 vccd1 net4565 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_179_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3304 net7964 vssd1 vssd1 vccd1 vccd1 net3831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4049 net4256 vssd1 vssd1 vccd1 vccd1 net4576 sky130_fd_sc_hd__clkbuf_2
Xhold3315 net7742 vssd1 vssd1 vccd1 vccd1 net3842 sky130_fd_sc_hd__buf_1
Xhold3326 _00748_ vssd1 vssd1 vccd1 vccd1 net3853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3337 _03085_ vssd1 vssd1 vccd1 vccd1 net3864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2603 _01581_ vssd1 vssd1 vccd1 vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3348 net626 vssd1 vssd1 vccd1 vccd1 net3875 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2614 net5960 vssd1 vssd1 vccd1 vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3359 _00623_ vssd1 vssd1 vccd1 vccd1 net3886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2625 net7491 vssd1 vssd1 vccd1 vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2636 net2866 vssd1 vssd1 vccd1 vccd1 net3163 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1902 net6718 vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 _03545_ vssd1 vssd1 vccd1 vccd1 net3174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 _01582_ vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 rbzero.pov.spi_buffer\[20\] vssd1 vssd1 vccd1 vccd1 net3185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 _04156_ vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2669 _03023_ vssd1 vssd1 vccd1 vccd1 net3196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 net7350 vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1946 _01440_ vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1957 _01364_ vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 net5693 vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1979 net3044 vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21803_ net245 net2980 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10__f_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ clknet_leaf_96_i_clk net4736 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19791__69 clknet_1_1__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21665_ clknet_leaf_122_i_clk net2192 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20616_ clknet_1_0__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__buf_1
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21596_ net230 net2362 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ net4083 net4862 vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5240 rbzero.debug_overlay.playerX\[-4\] vssd1 vssd1 vccd1 vccd1 net5767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5251 _00633_ vssd1 vssd1 vccd1 vccd1 net5778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5262 _04058_ vssd1 vssd1 vccd1 vccd1 net5789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5273 _02986_ vssd1 vssd1 vccd1 vccd1 net5800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5284 rbzero.pov.spi_buffer\[66\] vssd1 vssd1 vccd1 vccd1 net5811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5295 _02548_ vssd1 vssd1 vccd1 vccd1 net5822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4550 net701 vssd1 vssd1 vccd1 vccd1 net5077 sky130_fd_sc_hd__dlygate4sd3_1
X_22148_ clknet_leaf_51_i_clk _01635_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4561 rbzero.spi_registers.texadd1\[23\] vssd1 vssd1 vccd1 vccd1 net5088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4572 net734 vssd1 vssd1 vccd1 vccd1 net5099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4583 _00824_ vssd1 vssd1 vccd1 vccd1 net5110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4594 net731 vssd1 vssd1 vccd1 vccd1 net5121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3860 net8320 vssd1 vssd1 vccd1 vccd1 net4387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22079_ net521 net2252 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
Xhold3871 net7915 vssd1 vssd1 vccd1 vccd1 net4398 sky130_fd_sc_hd__dlygate4sd3_1
X_14970_ net4401 _07998_ _08079_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3893 net8173 vssd1 vssd1 vccd1 vccd1 net4420 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13921_ _06992_ _07029_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__and2_4
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ net3957 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__clkbuf_1
X_13852_ _07020_ _07021_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12803_ net7746 net4838 vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__nor2_1
X_16571_ _09657_ _09660_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__xnor2_1
X_20520__260 clknet_1_0__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__inv_2
X_13783_ _06720_ net577 vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10995_ net6345 net2845 _04238_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
X_18310_ net6428 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__clkbuf_1
X_15522_ _08611_ _08530_ _08616_ _08531_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__o31a_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19290_ net5161 _03236_ _03241_ _03230_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__o211a_1
X_12734_ _05904_ _05905_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _02456_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__clkbuf_1
X_15453_ _08544_ _08547_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__nand2_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12665_ _05837_ _05839_ _05840_ _05799_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a221o_2
XFILLER_0_155_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14404_ _07572_ _07574_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11616_ _04758_ _04759_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__nand2_1
X_18172_ net4526 net4496 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15384_ _08467_ _08471_ _08478_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__nand3_1
XFILLER_0_154_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ net4133 net4089 _05749_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17123_ _10034_ _10035_ _10142_ vssd1 vssd1 vccd1 vccd1 _10143_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03861_ _03861_ vssd1 vssd1 vccd1 vccd1 clknet_0__03861_ sky130_fd_sc_hd__clkbuf_16
X_14335_ _07455_ _07505_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11547_ net3982 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17054_ _10072_ _10074_ vssd1 vssd1 vccd1 vccd1 _10075_ sky130_fd_sc_hd__nor2_1
Xhold509 net5423 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ _07109_ _07342_ _07346_ _07363_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__a211o_1
X_11478_ net4132 _04667_ net4145 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_204_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16005_ _09088_ _09098_ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13217_ _06307_ _06387_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__or2_2
X_14197_ _07355_ _07367_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__nand2_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _06317_ _06318_ _06306_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__mux2_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17956_ _10316_ _09345_ _02099_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__or3_1
X_13079_ _06249_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__xor2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1209 net5539 vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16907_ _09927_ _09928_ vssd1 vssd1 vccd1 vccd1 _09929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17887_ _01983_ _01990_ _01988_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a21oi_1
X_20603__335 clknet_1_1__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__inv_2
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ net6542 net3816 _03430_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
X_16838_ _09858_ _09861_ _09845_ vssd1 vssd1 vccd1 vccd1 _09863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ _08980_ _08982_ _09800_ vssd1 vssd1 vccd1 vccd1 _09801_ sky130_fd_sc_hd__a21o_1
X_19557_ net6816 net1622 net1882 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
X_18508_ _02666_ _02672_ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a21oi_1
X_19488_ net1626 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18439_ net3604 rbzero.wall_tracer.rayAddendX\[1\] net4724 vssd1 vssd1 vccd1 vccd1
+ _02620_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21450_ clknet_leaf_38_i_clk net1584 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21381_ clknet_leaf_3_i_clk net5003 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20332_ net6178 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20263_ _05673_ _09733_ net4096 _03794_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a22o_1
X_22002_ net444 net2621 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold3101 _04655_ vssd1 vssd1 vccd1 vccd1 net3628 sky130_fd_sc_hd__clkbuf_2
Xhold3112 _02595_ vssd1 vssd1 vccd1 vccd1 net3639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20194_ _03728_ net3662 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__or2_1
Xhold3123 _00522_ vssd1 vssd1 vccd1 vccd1 net3650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3134 _05151_ vssd1 vssd1 vccd1 vccd1 net3661 sky130_fd_sc_hd__clkbuf_4
Xhold2400 net2863 vssd1 vssd1 vccd1 vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3145 _03318_ vssd1 vssd1 vccd1 vccd1 net3672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 _04341_ vssd1 vssd1 vccd1 vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3156 _06059_ vssd1 vssd1 vccd1 vccd1 net3683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2422 _01533_ vssd1 vssd1 vccd1 vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3167 rbzero.spi_registers.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 net3694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2433 _04119_ vssd1 vssd1 vccd1 vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3178 _03494_ vssd1 vssd1 vccd1 vccd1 net3705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03850_ clknet_0__03850_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03850_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2444 _04214_ vssd1 vssd1 vccd1 vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3189 net5831 vssd1 vssd1 vccd1 vccd1 net3716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1710 _01385_ vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2455 _04072_ vssd1 vssd1 vccd1 vccd1 net2982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1721 net7010 vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2466 net7440 vssd1 vssd1 vccd1 vccd1 net2993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1732 net7062 vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2477 _00948_ vssd1 vssd1 vccd1 vccd1 net3004 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1743 _00983_ vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2488 net5897 vssd1 vssd1 vccd1 vccd1 net3015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 _01080_ vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2499 net2262 vssd1 vssd1 vccd1 vccd1 net3026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1765 _04251_ vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1776 net2946 vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20578__312 clknet_1_1__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__inv_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1787 _01157_ vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1798 _04096_ vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10780_ net6116 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__clkbuf_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ clknet_leaf_103_i_clk net4597 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _05632_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21648_ clknet_leaf_126_i_clk net2803 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ _04558_ _04559_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__nor2_1
X_12381_ rbzero.tex_b1\[3\] rbzero.tex_b1\[2\] _04924_ vssd1 vssd1 vccd1 vccd1 _05566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21579_ net213 net1984 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_80 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_91 net4912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _07288_ _07289_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11332_ rbzero.spi_registers.texadd3\[6\] rbzero.spi_registers.texadd1\[6\] rbzero.spi_registers.texadd0\[6\]
+ rbzero.spi_registers.texadd2\[6\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__mux4_2
XFILLER_0_160_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ _07164_ _07174_ _07172_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__a21oi_1
X_11263_ _04459_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_8
Xhold5070 _00498_ vssd1 vssd1 vccd1 vccd1 net5597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5081 rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 net5608 sky130_fd_sc_hd__dlygate4sd3_1
X_13002_ net4565 _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nor2_1
X_11194_ _04264_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__clkbuf_4
Xhold5092 _00389_ vssd1 vssd1 vccd1 vccd1 net5619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4380 net4705 vssd1 vssd1 vccd1 vccd1 net4907 sky130_fd_sc_hd__clkbuf_1
X_17810_ _02047_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__or2_2
Xhold4391 _08130_ vssd1 vssd1 vccd1 vccd1 net4918 sky130_fd_sc_hd__dlymetal6s2s_1
X_18790_ _02935_ _02936_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17741_ _08167_ _10289_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__nor2_1
Xhold3690 net8303 vssd1 vssd1 vccd1 vccd1 net4217 sky130_fd_sc_hd__dlygate4sd3_1
X_14953_ net4583 _07938_ _08068_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__mux2_1
X_13904_ _06706_ _06771_ _06796_ _06703_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__o22a_1
X_17672_ _01910_ _01911_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__nor2_1
X_14884_ _08033_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
X_20444__191 clknet_1_1__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__inv_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16623_ _09105_ net4189 vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__xnor2_1
X_19411_ net1733 net3902 _03141_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _07004_ _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap82 _06464_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_6
XFILLER_0_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16554_ _09640_ _09643_ vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__xnor2_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ net6275 _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__or2_1
X_13766_ _06935_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ net2716 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15505_ _08537_ _08538_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__or2_1
X_19273_ net5057 _03200_ _03229_ _03230_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__o211a_1
X_12717_ net32 net33 _05876_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__and4_1
X_16485_ _09461_ _09575_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__xor2_4
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13697_ net79 _06769_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _02441_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15436_ _08529_ _08142_ _08132_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__or3b_1
XFILLER_0_26_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ net25 _05823_ _05826_ _05801_ net26 vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18155_ net4567 net4461 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15367_ rbzero.wall_tracer.visualWallDist\[-10\] _08117_ vssd1 vssd1 vccd1 vccd1
+ _08462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ net4128 _05043_ net16 vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__mux2_1
X_17106_ _09891_ _10126_ vssd1 vssd1 vccd1 vccd1 _10127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03844_ _03844_ vssd1 vssd1 vccd1 vccd1 clknet_0__03844_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14318_ _06754_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__clkbuf_4
X_18086_ _02318_ net3749 _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
X_15298_ _08389_ _08391_ _08392_ _08221_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__o22ai_1
Xhold306 net5329 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold317 net5200 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 net5381 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17037_ _10024_ _10057_ vssd1 vssd1 vccd1 vccd1 _10058_ sky130_fd_sc_hd__xnor2_2
Xhold339 net5251 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14249_ _06758_ _07342_ _07419_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ net3159 net7587 _03058_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _03347_ vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 net6447 vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _02174_ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nor2_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 net6551 vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 _00913_ vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20950_ clknet_leaf_63_i_clk _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19609_ net3770 _02472_ net92 net1777 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__and4_1
X_20881_ net4879 _02508_ _02559_ net8249 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21502_ clknet_leaf_15_i_clk net1268 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21433_ clknet_leaf_40_i_clk net2258 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21364_ clknet_leaf_4_i_clk net5015 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_20674__19 clknet_1_1__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_0_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20315_ net6570 net3592 _03825_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21295_ clknet_leaf_35_i_clk net5394 vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold840 net4231 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold851 _03432_ vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 net6330 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold873 net6137 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_20246_ net3337 net5984 _03788_ _03783_ _03689_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_102_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold884 net6266 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 net6334 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ net7565 _03743_ net4417 _03732_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__o211a_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2230 _01505_ vssd1 vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 _04087_ vssd1 vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2252 _01318_ vssd1 vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2263 net2040 vssd1 vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2274 net1145 vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2285 _01468_ vssd1 vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1540 _03158_ vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2296 net5648 vssd1 vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1551 rbzero.pov.ready_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ rbzero.debug_overlay.facingX\[-5\] _05108_ _05114_ rbzero.debug_overlay.facingX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a22o_1
Xhold1562 _03041_ vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1573 _00939_ vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1584 net6712 vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10901_ net7057 net7033 _04265_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1595 net6962 vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_108 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_108/HI o_rgb[19]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_119 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_119/HI zeros[8] sky130_fd_sc_hd__conb_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ net4117 _05066_ net3517 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__and3b_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _06788_ _06789_ _06790_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ net3250 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _06589_ _06590_ _06607_ _06617_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__a211oi_4
X_10763_ net6245 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net9 net8 _05658_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__and4_1
X_16270_ _09360_ _09361_ vssd1 vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__nor2_1
X_13482_ _06652_ _06566_ _06492_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__mux2_1
X_10694_ net6152 net3356 _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15221_ net4399 _08124_ _06119_ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__a21oi_1
X_12433_ _05465_ _04949_ _05031_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__a21oi_1
X_20632__361 clknet_1_1__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__inv_2
XFILLER_0_63_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ _08243_ _08244_ _08245_ _08246_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _05250_ vssd1 vssd1 vccd1 vccd1 _05549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14103_ _07272_ _07273_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__and2_1
X_11315_ _04504_ _04505_ rbzero.spi_registers.texadd3\[14\] vssd1 vssd1 vccd1 vccd1
+ _04507_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19960_ net3010 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
X_15083_ _06033_ _08177_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12295_ _05233_ _05476_ _05480_ _05263_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14034_ _06576_ _06914_ net3579 vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__o21ai_1
X_18911_ net1916 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
X_11246_ net7260 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19891_ net1359 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18842_ net3485 _02947_ _02979_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__and3_1
X_11177_ net2674 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15985_ _08759_ _08656_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__and2b_1
X_18773_ _02919_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17724_ _01741_ _01943_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nand2_1
X_14936_ net3933 _06235_ net1791 vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__o21ai_1
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17655_ _10062_ _09181_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__or2_1
X_14867_ net7794 _07967_ _08019_ _08020_ _07869_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__a221o_2
XFILLER_0_188_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _09653_ _09695_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__xnor2_2
X_13818_ net537 _06986_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__or2b_1
XFILLER_0_203_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17586_ _01680_ _01705_ _01703_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14798_ net7824 _07960_ net7806 vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16537_ _09624_ _09625_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__and2_1
X_19325_ net1602 _03251_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13749_ _06915_ _06916_ _06917_ _06919_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16468_ _09533_ _09558_ vssd1 vssd1 vccd1 vccd1 _09559_ sky130_fd_sc_hd__xnor2_1
X_19256_ net5145 _03216_ _03221_ _03219_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__o211a_1
Xhold7208 rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 net7735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7219 net4002 vssd1 vssd1 vccd1 vccd1 net7746 sky130_fd_sc_hd__clkbuf_2
X_15419_ _08502_ _08503_ _08513_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__a21bo_1
X_18207_ _02426_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__clkbuf_1
X_19187_ net5240 _03168_ _03180_ _03176_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__o211a_1
X_16399_ _09488_ _09489_ vssd1 vssd1 vccd1 vccd1 _09490_ sky130_fd_sc_hd__nor2_1
Xhold6507 rbzero.tex_r0\[6\] vssd1 vssd1 vccd1 vccd1 net7034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6518 net2125 vssd1 vssd1 vccd1 vccd1 net7045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6529 rbzero.tex_g0\[44\] vssd1 vssd1 vccd1 vccd1 net7056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18138_ net3768 net4392 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5806 net1390 vssd1 vssd1 vccd1 vccd1 net6333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5817 rbzero.tex_b1\[62\] vssd1 vssd1 vccd1 vccd1 net6344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 net6033 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5828 net1286 vssd1 vssd1 vccd1 vccd1 net6355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 net4969 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5839 rbzero.spi_registers.new_texadd\[0\]\[5\] vssd1 vssd1 vccd1 vccd1 net6366
+ sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ _02266_ _02304_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__xnor2_1
Xhold125 net8096 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold136 net7464 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold147 net4802 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ _03690_ _03691_ _03484_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a21oi_1
Xhold158 net5016 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ clknet_leaf_70_i_clk _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold169 net5086 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20031_ net5907 _03615_ _03606_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__o211a_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20460__206 clknet_1_0__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__inv_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21982_ net424 net2909 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20933_ clknet_leaf_78_i_clk net4685 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20864_ _03312_ net1093 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20795_ _03878_ _03962_ _03963_ _03883_ net5692 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7720 _02939_ vssd1 vssd1 vccd1 vccd1 net8247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7731 _02672_ vssd1 vssd1 vccd1 vccd1 net8258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7742 net8029 vssd1 vssd1 vccd1 vccd1 net8269 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7775 net4216 vssd1 vssd1 vccd1 vccd1 net8302 sky130_fd_sc_hd__dlygate4sd3_1
X_21416_ clknet_leaf_2_i_clk net3908 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7786 net4340 vssd1 vssd1 vccd1 vccd1 net8313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7797 net4402 vssd1 vssd1 vccd1 vccd1 net8324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21347_ clknet_leaf_13_i_clk net5270 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11100_ net6271 net2978 _04364_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__mux2_1
X_12080_ rbzero.tex_r1\[55\] rbzero.tex_r1\[54\] _05237_ vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__mux2_1
Xhold670 net6459 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21278_ clknet_leaf_27_i_clk net5538 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold681 _01498_ vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold692 net6179 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net2000 net6118 _04331_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20229_ _04459_ net3679 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__or2_1
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 net8150 vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 net3815 vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2082 _01047_ vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _08253_ _08464_ _08573_ _08864_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__a22o_1
X_19812__87 clknet_1_1__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__inv_2
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2093 _04154_ vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ net4779 _06148_ _06150_ _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 net6829 vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1381 _00694_ vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ _07843_ _07883_ _07885_ _07890_ net7839 vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__a311o_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ net3372 _05102_ _05108_ rbzero.debug_overlay.playerY\[-5\] _05121_ vssd1
+ vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__a221o_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 net5610 vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _09537_ _10346_ _10350_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__or3_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _06699_ _07807_ _07305_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11864_ net45 vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__buf_6
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13603_ _06772_ _06773_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__xor2_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _10287_ _10290_ _10285_ vssd1 vssd1 vccd1 vccd1 _10389_ sky130_fd_sc_hd__a21oi_1
X_10815_ net2522 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _07489_ _07391_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__nor2_1
X_11795_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _04979_ vssd1 vssd1 vccd1 vccd1 _04985_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19110_ net1817 _03125_ net5527 _03128_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__o211a_1
X_16322_ _07989_ _07979_ _08027_ _08020_ _07869_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__a221oi_2
X_13534_ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__clkbuf_4
X_10746_ net7262 net7427 _04182_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20556__292 clknet_1_0__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__inv_2
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19041_ net3399 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__clkbuf_1
X_16253_ _09344_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__buf_4
X_13465_ _06538_ _06599_ _06602_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ net7220 net7129 _04149_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15204_ net4284 net3445 _08256_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__or3_4
X_12416_ _04922_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ _09275_ _09276_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13396_ _06565_ _06566_ _06551_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15135_ net3317 net4344 _08188_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__or3_1
X_12347_ _05527_ _05529_ _05532_ _05233_ _04942_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03512_ clknet_0__03512_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03512_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15066_ _08160_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__buf_2
X_19943_ net3061 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
X_12278_ net5049 net7719 _04845_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _07186_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__xnor2_1
X_11229_ net2346 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19874_ net1689 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
X_18825_ net5845 _02947_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18756_ _02865_ net3761 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__or2_1
X_15968_ _08127_ _09062_ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__or2_1
X_17707_ _01944_ _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14919_ net4589 _08050_ _08052_ net3751 net4695 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__o221a_1
XFILLER_0_210_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15899_ _08399_ _08359_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__or2b_1
X_18687_ _02839_ _02840_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17638_ _01876_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20639__367 clknet_1_0__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__inv_2
XFILLER_0_37_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _01808_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19308_ net1435 _03251_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__05946_ clknet_0__05946_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05946_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7005 net3246 vssd1 vssd1 vccd1 vccd1 net7532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7016 rbzero.pov.ready_buffer\[28\] vssd1 vssd1 vccd1 vccd1 net7543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7027 net2764 vssd1 vssd1 vccd1 vccd1 net7554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19239_ net5141 _03201_ _03211_ _03206_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__o211a_1
Xhold7038 net876 vssd1 vssd1 vccd1 vccd1 net7565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6304 _04427_ vssd1 vssd1 vccd1 vccd1 net6831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7049 _02730_ vssd1 vssd1 vccd1 vccd1 net7576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6315 net1846 vssd1 vssd1 vccd1 vccd1 net6842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6326 rbzero.tex_g0\[36\] vssd1 vssd1 vccd1 vccd1 net6853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6337 net2269 vssd1 vssd1 vccd1 vccd1 net6864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5603 net1018 vssd1 vssd1 vccd1 vccd1 net6130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6348 _04314_ vssd1 vssd1 vccd1 vccd1 net6875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6359 net2015 vssd1 vssd1 vccd1 vccd1 net6886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5614 _04047_ vssd1 vssd1 vccd1 vccd1 net6141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5625 net1089 vssd1 vssd1 vccd1 vccd1 net6152 sky130_fd_sc_hd__dlygate4sd3_1
X_21201_ clknet_leaf_116_i_clk net3133 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5636 rbzero.tex_g0\[42\] vssd1 vssd1 vccd1 vccd1 net6163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4902 _00388_ vssd1 vssd1 vccd1 vccd1 net5429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5647 net1073 vssd1 vssd1 vccd1 vccd1 net6174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5658 _04371_ vssd1 vssd1 vccd1 vccd1 net6185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4913 net1050 vssd1 vssd1 vccd1 vccd1 net5440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5669 rbzero.tex_g0\[12\] vssd1 vssd1 vccd1 vccd1 net6196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4924 rbzero.spi_registers.vshift\[5\] vssd1 vssd1 vccd1 vccd1 net5451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4935 net1137 vssd1 vssd1 vccd1 vccd1 net5462 sky130_fd_sc_hd__dlygate4sd3_1
X_21132_ clknet_leaf_29_i_clk net4036 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_1
Xhold4946 _00525_ vssd1 vssd1 vccd1 vccd1 net5473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4957 net1209 vssd1 vssd1 vccd1 vccd1 net5484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4968 rbzero.pov.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 net5495 sky130_fd_sc_hd__dlygate4sd3_1
X_21063_ clknet_leaf_60_i_clk _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4979 _00771_ vssd1 vssd1 vccd1 vccd1 net5506 sky130_fd_sc_hd__dlygate4sd3_1
X_20384__137 clknet_1_1__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__inv_2
X_20014_ net5849 _08263_ _03614_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21965_ net407 net2290 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ clknet_leaf_66_i_clk _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21896_ net338 net1082 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20847_ _04000_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__buf_1
XFILLER_0_194_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ net2531 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__clkbuf_1
X_11580_ _04766_ _04767_ net1284 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20778_ net1009 net5622 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10531_ net1939 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7550 _00602_ vssd1 vssd1 vccd1 vccd1 net8077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ net8275 _06266_ _06264_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__o21a_1
X_10462_ net2349 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7561 net4912 vssd1 vssd1 vccd1 vccd1 net8088 sky130_fd_sc_hd__buf_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7572 rbzero.wall_tracer.rayAddendY\[-8\] vssd1 vssd1 vccd1 vccd1 net8099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7583 _00604_ vssd1 vssd1 vccd1 vccd1 net8110 sky130_fd_sc_hd__dlygate4sd3_1
X_12201_ _04930_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or2_1
Xhold7594 _00511_ vssd1 vssd1 vccd1 vccd1 net8121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6860 net2917 vssd1 vssd1 vccd1 vccd1 net7387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13181_ _06335_ _06337_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a21oi_2
Xhold6871 rbzero.tex_g1\[35\] vssd1 vssd1 vccd1 vccd1 net7398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6882 net2943 vssd1 vssd1 vccd1 vccd1 net7409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6893 _02996_ vssd1 vssd1 vccd1 vccd1 net7420 sky130_fd_sc_hd__dlygate4sd3_1
X_12132_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _04933_ vssd1 vssd1 vccd1 vccd1 _05320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _09956_ _09961_ vssd1 vssd1 vccd1 vccd1 _09962_ sky130_fd_sc_hd__xor2_1
X_12063_ rbzero.tex_r1\[35\] rbzero.tex_r1\[34\] _05237_ vssd1 vssd1 vccd1 vccd1 _05252_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ net2545 net7157 _04320_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__mux2_1
X_16871_ _09891_ _09892_ vssd1 vssd1 vccd1 vccd1 _09893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18610_ _05164_ net4423 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__or2_1
X_15822_ _08916_ _08329_ _08897_ _08900_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__o31a_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ net6742 net3562 net1779 vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19797__75 clknet_1_0__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _08830_ _08847_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__xor2_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18541_ net4053 _09788_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__o21ai_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _06068_ net4642 _06138_ _06139_ _06140_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a2111o_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _05067_ _05098_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__or2_1
X_14704_ _07828_ _07816_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15684_ _08767_ _08769_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__nand2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _02634_ _02649_ _02647_ _04481_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a31o_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ net4436 _06043_ net4044 _04674_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _08326_ _09664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__nor2_1
X_14635_ _06839_ _07251_ _07305_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__a21oi_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ _05018_ _05036_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__nand2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _10371_ _10372_ vssd1 vssd1 vccd1 vccd1 _10373_ sky130_fd_sc_hd__xor2_2
X_14566_ _07734_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__nand2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _04836_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16305_ _09286_ _09290_ _09287_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__o21ai_1
X_13517_ _06343_ _06564_ net562 vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__and3_1
X_17285_ _10302_ _10303_ vssd1 vssd1 vccd1 vccd1 _10304_ sky130_fd_sc_hd__nor2_1
X_10729_ net2049 net6818 _04097_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14497_ _07665_ _07667_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__nor2_1
X_19024_ net4017 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
X_16236_ _09326_ net5769 vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__or2_1
X_13448_ _06441_ _06549_ _06614_ _06491_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16167_ _08389_ _08309_ _08392_ _08308_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ net82 _06489_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or2_2
Xhold4209 net639 vssd1 vssd1 vccd1 vccd1 net4736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15118_ _08187_ _08208_ _08212_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__a21bo_2
X_16098_ _09189_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3508 _02736_ vssd1 vssd1 vccd1 vccd1 net4035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3519 _00615_ vssd1 vssd1 vccd1 vccd1 net4046 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_8__f_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15049_ _08132_ _08143_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__nand2_1
X_19926_ net5710 net7367 _03572_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2807 _03381_ vssd1 vssd1 vccd1 vccd1 net3334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2818 net7604 vssd1 vssd1 vccd1 vccd1 net3345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 net7517 vssd1 vssd1 vccd1 vccd1 net3356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19857_ net1707 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
X_18808_ net3695 net5799 _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__or3_1
XFILLER_0_183_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19788_ clknet_1_1__leaf__03506_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_89_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18739_ _02873_ _02888_ _02886_ _04481_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21750_ clknet_leaf_99_i_clk net3681 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20701_ _03880_ _03881_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21681_ clknet_leaf_113_i_clk net5820 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6101 rbzero.spi_registers.new_texadd\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net6628
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6112 net1828 vssd1 vssd1 vccd1 vccd1 net6639 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_27_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold6123 rbzero.tex_r0\[33\] vssd1 vssd1 vccd1 vccd1 net6650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20494_ clknet_1_1__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__buf_1
Xhold6134 net1579 vssd1 vssd1 vccd1 vccd1 net6661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5400 net3309 vssd1 vssd1 vccd1 vccd1 net5927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6145 rbzero.tex_b0\[25\] vssd1 vssd1 vccd1 vccd1 net6672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6156 net2220 vssd1 vssd1 vccd1 vccd1 net6683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5411 _02714_ vssd1 vssd1 vccd1 vccd1 net5938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6167 _03000_ vssd1 vssd1 vccd1 vccd1 net6694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5422 _09729_ vssd1 vssd1 vccd1 vccd1 net5949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6178 net1872 vssd1 vssd1 vccd1 vccd1 net6705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5433 rbzero.wall_tracer.rayAddendX\[-4\] vssd1 vssd1 vccd1 vccd1 net5960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6189 _04081_ vssd1 vssd1 vccd1 vccd1 net6716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5444 _02605_ vssd1 vssd1 vccd1 vccd1 net5971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5455 _05678_ vssd1 vssd1 vccd1 vccd1 net5982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4710 _00785_ vssd1 vssd1 vccd1 vccd1 net5237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4721 net818 vssd1 vssd1 vccd1 vccd1 net5248 sky130_fd_sc_hd__dlygate4sd3_1
X_22164_ clknet_leaf_96_i_clk net4426 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5466 rbzero.spi_registers.new_sky\[0\] vssd1 vssd1 vccd1 vccd1 net5993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5477 rbzero.spi_registers.new_sky\[4\] vssd1 vssd1 vccd1 vccd1 net6004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4732 rbzero.spi_registers.texadd2\[10\] vssd1 vssd1 vccd1 vccd1 net5259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5488 net3734 vssd1 vssd1 vccd1 vccd1 net6015 sky130_fd_sc_hd__clkbuf_2
Xhold4743 net802 vssd1 vssd1 vccd1 vccd1 net5270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5499 net623 vssd1 vssd1 vccd1 vccd1 net6026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4754 _01015_ vssd1 vssd1 vccd1 vccd1 net5281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21115_ clknet_leaf_93_i_clk net4728 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold4765 net911 vssd1 vssd1 vccd1 vccd1 net5292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4776 rbzero.spi_registers.texadd2\[22\] vssd1 vssd1 vccd1 vccd1 net5303 sky130_fd_sc_hd__dlygate4sd3_1
X_22095_ net157 net2440 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
Xhold4787 net932 vssd1 vssd1 vccd1 vccd1 net5314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4798 _00792_ vssd1 vssd1 vccd1 vccd1 net5325 sky130_fd_sc_hd__dlygate4sd3_1
X_21046_ clknet_leaf_58_i_clk _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12750_ net4111 _05673_ net4071 net4092 _05901_ net36 vssd1 vssd1 vccd1 vccd1 _05927_
+ sky130_fd_sc_hd__mux4_1
X_21948_ net390 net2972 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ net3405 net3955 _04584_ net3406 _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__o221a_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ net4149 net4141 net4164 net7727 _05851_ net31 vssd1 vssd1 vccd1 vccd1 _05859_
+ sky130_fd_sc_hd__mux4_1
X_21879_ net321 net2219 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _07072_ net569 _07281_ _06754_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__o22ai_2
X_11632_ _04776_ _04801_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__and2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _07240_ _07390_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11563_ net1079 net1228 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _06398_ _06403_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nor2_1
X_17070_ _10084_ _10085_ _10090_ vssd1 vssd1 vccd1 vccd1 _10091_ sky130_fd_sc_hd__o21a_1
X_10514_ net5645 net7295 _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__mux2_1
X_14282_ _07451_ _07452_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ net4106 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__buf_4
X_16021_ _06122_ _09114_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__or2_1
X_13233_ _06382_ _06383_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__nand2_4
Xhold7380 net3406 vssd1 vssd1 vccd1 vccd1 net7907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7391 rbzero.wall_tracer.stepDistY\[3\] vssd1 vssd1 vccd1 vccd1 net7918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ net4133 net4089 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6690 rbzero.tex_b1\[41\] vssd1 vssd1 vccd1 vccd1 net7217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13164_ _06305_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _05258_ vssd1 vssd1 vccd1 vccd1 _05303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17972_ _02203_ _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__nand2_1
X_13095_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19711_ net6209 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__clkbuf_1
X_16923_ _09943_ _09944_ vssd1 vssd1 vccd1 vccd1 _09945_ sky130_fd_sc_hd__xor2_1
X_12046_ rbzero.tex_r1\[29\] rbzero.tex_r1\[28\] _05220_ vssd1 vssd1 vccd1 vccd1 _05235_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19642_ net1771 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__clkbuf_1
X_16854_ net4581 net4397 vssd1 vssd1 vccd1 vccd1 _09877_ sky130_fd_sc_hd__nor2_1
X_15805_ _08417_ _08691_ _08899_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__or3b_1
XFILLER_0_172_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19573_ net2105 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
X_16785_ net4569 net4485 vssd1 vssd1 vccd1 vccd1 _09815_ sky130_fd_sc_hd__nand2_1
X_13997_ _06673_ _06698_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18524_ _02697_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__xor2_1
X_15736_ _08821_ _08822_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__xor2_1
X_12948_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__buf_4
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18455_ _02633_ _02634_ _02607_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a21oi_1
X_15667_ _08754_ _08761_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__nand2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ net3975 _04476_ net3871 vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or3b_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _10406_ _10423_ vssd1 vssd1 vccd1 vccd1 _10424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _07511_ _07787_ _07788_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__o21bai_4
X_15598_ _08342_ _08345_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__xor2_2
X_18386_ net3509 _05155_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__xor2_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17337_ _10218_ _10230_ _10229_ vssd1 vssd1 vccd1 vccd1 _10356_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14549_ _07710_ _07718_ _07719_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17268_ _10285_ _10286_ vssd1 vssd1 vccd1 vccd1 _10287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20415__166 clknet_1_0__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__inv_2
XFILLER_0_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ net7512 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16219_ _09153_ _09193_ _09192_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_183_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17199_ _09666_ _09667_ vssd1 vssd1 vccd1 vccd1 _10219_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__05645_ clknet_0__05645_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05645_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4006 net1003 vssd1 vssd1 vccd1 vccd1 net4533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4017 _00413_ vssd1 vssd1 vccd1 vccd1 net4544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4028 _03762_ vssd1 vssd1 vccd1 vccd1 net4555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4039 net7955 vssd1 vssd1 vccd1 vccd1 net4566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3305 net8339 vssd1 vssd1 vccd1 vccd1 net3832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3316 _03421_ vssd1 vssd1 vccd1 vccd1 net3843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3327 net7988 vssd1 vssd1 vccd1 vccd1 net3854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3338 _00727_ vssd1 vssd1 vccd1 vccd1 net3865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3349 rbzero.spi_registers.spi_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net3876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2604 net7460 vssd1 vssd1 vccd1 vccd1 net3131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 net5962 vssd1 vssd1 vccd1 vccd1 net3142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2626 net7493 vssd1 vssd1 vccd1 vccd1 net3153 sky130_fd_sc_hd__dlygate4sd3_1
X_19909_ net3260 net2974 _03561_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__mux2_1
Xhold2637 _04325_ vssd1 vssd1 vccd1 vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1903 net6720 vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 _01111_ vssd1 vssd1 vccd1 vccd1 net3175 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03509_ _03509_ vssd1 vssd1 vccd1 vccd1 clknet_0__03509_ sky130_fd_sc_hd__clkbuf_16
Xhold2659 net1946 vssd1 vssd1 vccd1 vccd1 net3186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1914 net6004 vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1925 _01487_ vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1936 net5663 vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1947 net5621 vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__buf_1
Xhold1958 net6953 vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 net6951 vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19776__56 clknet_1_0__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21802_ net244 net1227 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20496__238 clknet_1_1__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__inv_2
XFILLER_0_151_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21733_ clknet_leaf_96_i_clk net4805 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21664_ clknet_leaf_23_i_clk net2929 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21595_ net229 net2650 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5230 net2630 vssd1 vssd1 vccd1 vccd1 net5757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5241 net3339 vssd1 vssd1 vccd1 vccd1 net5768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5252 net3967 vssd1 vssd1 vccd1 vccd1 net5779 sky130_fd_sc_hd__clkbuf_1
Xhold5263 net585 vssd1 vssd1 vccd1 vccd1 net5790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5274 _00645_ vssd1 vssd1 vccd1 vccd1 net5801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4540 net720 vssd1 vssd1 vccd1 vccd1 net5067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5285 net1709 vssd1 vssd1 vccd1 vccd1 net5812 sky130_fd_sc_hd__dlygate4sd3_1
X_22147_ clknet_leaf_53_i_clk _01634_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5296 net3635 vssd1 vssd1 vccd1 vccd1 net5823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4551 _00815_ vssd1 vssd1 vccd1 vccd1 net5078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4562 net842 vssd1 vssd1 vccd1 vccd1 net5089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4573 rbzero.spi_registers.texadd3\[14\] vssd1 vssd1 vccd1 vccd1 net5100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4584 net798 vssd1 vssd1 vccd1 vccd1 net5111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3850 net3474 vssd1 vssd1 vccd1 vccd1 net4377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4595 _00797_ vssd1 vssd1 vccd1 vccd1 net5122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3861 net8322 vssd1 vssd1 vccd1 vccd1 net4388 sky130_fd_sc_hd__buf_1
X_22078_ net520 net2375 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold3872 net7917 vssd1 vssd1 vccd1 vccd1 net4399 sky130_fd_sc_hd__buf_1
XFILLER_0_195_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3883 net7945 vssd1 vssd1 vccd1 vccd1 net4410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3894 _00769_ vssd1 vssd1 vccd1 vccd1 net4421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21029_ clknet_leaf_53_i_clk net4235 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13920_ _07071_ _07089_ _07090_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13851_ _07020_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12802_ net7744 net6046 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16570_ _09658_ _09659_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__nor2_1
X_13782_ _06917_ _06919_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__xnor2_1
X_10994_ net2846 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ _08535_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__clkbuf_4
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _05906_ _05907_ _05908_ _05909_ net38 vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a32o_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15452_ _08546_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__inv_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ _02455_ net3835 _02393_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05797_ _05802_ _05841_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a31o_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ _07571_ _07573_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11615_ _04769_ _04803_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a21o_1
X_15383_ _08414_ _08433_ _08476_ _08477_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__a31o_1
X_18171_ net4526 net4496 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12595_ _04648_ _04461_ _04468_ _04023_ _05749_ _05747_ vssd1 vssd1 vccd1 vccd1 _05775_
+ sky130_fd_sc_hd__mux4_1
X_17122_ _10036_ _10037_ vssd1 vssd1 vccd1 vccd1 _10142_ sky130_fd_sc_hd__or2b_1
XFILLER_0_170_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03860_ _03860_ vssd1 vssd1 vccd1 vccd1 clknet_0__03860_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _07456_ _07501_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__o21a_1
X_11546_ _04727_ _04730_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__and3b_1
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17053_ _09945_ _09946_ _10073_ vssd1 vssd1 vccd1 vccd1 _10074_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ _07341_ _07353_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ net4105 _04666_ net4115 net3516 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__o211a_1
X_16004_ _09088_ _09098_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__or2_1
X_13216_ net8015 _06266_ _06264_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__o21a_1
XFILLER_0_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14196_ _07359_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ net4293 _05997_ _06265_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__mux2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17955_ _10316_ _09225_ _09345_ _08472_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__o22a_1
X_13078_ _06051_ _06250_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or3_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16906_ _09650_ _09895_ _09926_ vssd1 vssd1 vccd1 vccd1 _09928_ sky130_fd_sc_hd__nand3_1
X_12029_ rbzero.tex_r1\[15\] rbzero.tex_r1\[14\] _04979_ vssd1 vssd1 vccd1 vccd1 _05218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17886_ _02113_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__xnor2_1
X_19625_ net1296 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
X_16837_ _09858_ _09861_ vssd1 vssd1 vccd1 vccd1 _09862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19556_ _04458_ net1881 vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__nor2_1
X_16768_ _08980_ _08982_ _06057_ vssd1 vssd1 vccd1 vccd1 _09800_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18507_ _02681_ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__nand2_1
X_15719_ _08200_ _08318_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__nor2_1
X_19487_ net1426 net6056 _03354_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__mux2_1
X_16699_ net1009 _09745_ _09746_ net8012 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18438_ net4724 rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02619_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18369_ _02553_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21380_ clknet_leaf_9_i_clk net5027 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20331_ net6176 net3631 _03813_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20262_ net4113 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22001_ net443 net1522 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3102 _01623_ vssd1 vssd1 vccd1 vccd1 net3629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3113 net4727 vssd1 vssd1 vccd1 vccd1 net3640 sky130_fd_sc_hd__dlygate4sd3_1
X_20193_ net3661 net2161 _03723_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3124 net7724 vssd1 vssd1 vccd1 vccd1 net3651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3135 _03755_ vssd1 vssd1 vccd1 vccd1 net3662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2401 _03589_ vssd1 vssd1 vccd1 vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3146 _00888_ vssd1 vssd1 vccd1 vccd1 net3673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2412 _01320_ vssd1 vssd1 vccd1 vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3157 net7606 vssd1 vssd1 vccd1 vccd1 net3684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2423 net7325 vssd1 vssd1 vccd1 vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3168 net3394 vssd1 vssd1 vccd1 vccd1 net3695 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2434 _01521_ vssd1 vssd1 vccd1 vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3179 _01016_ vssd1 vssd1 vccd1 vccd1 net3706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2445 _01435_ vssd1 vssd1 vccd1 vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 net6819 vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 rbzero.tex_b1\[27\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2456 _01560_ vssd1 vssd1 vccd1 vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1722 _01522_ vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2467 _04129_ vssd1 vssd1 vccd1 vccd1 net2994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 net7412 vssd1 vssd1 vccd1 vccd1 net3005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _04057_ vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1744 net6921 vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2489 _03071_ vssd1 vssd1 vccd1 vccd1 net3016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1755 net7166 vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1766 _01401_ vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1777 _04107_ vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 net7022 vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1799 _01538_ vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21716_ clknet_leaf_127_i_clk net3610 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21647_ clknet_leaf_126_i_clk net1887 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11400_ _04591_ _04557_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12380_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _05369_ vssd1 vssd1 vccd1 vccd1 _05565_
+ sky130_fd_sc_hd__mux2_1
X_21578_ net212 net2806 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_70 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11331_ rbzero.texu_hot\[1\] _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_92 net8002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050_ _07203_ _07220_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5060 _04373_ vssd1 vssd1 vccd1 vccd1 net5587 sky130_fd_sc_hd__dlygate4sd3_1
X_13001_ net4541 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__inv_2
Xhold5071 net5676 vssd1 vssd1 vccd1 vccd1 net5598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5082 net1918 vssd1 vssd1 vccd1 vccd1 net5609 sky130_fd_sc_hd__dlygate4sd3_1
X_11193_ net6944 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__clkbuf_1
Xhold5093 net2059 vssd1 vssd1 vccd1 vccd1 net5620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4370 net3668 vssd1 vssd1 vccd1 vccd1 net4897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4381 _09223_ vssd1 vssd1 vccd1 vccd1 net4908 sky130_fd_sc_hd__clkbuf_2
Xhold4392 rbzero.wall_tracer.trackDistX\[-3\] vssd1 vssd1 vccd1 vccd1 net4919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3680 net8134 vssd1 vssd1 vccd1 vccd1 net4207 sky130_fd_sc_hd__dlygate4sd3_1
X_17740_ _01977_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__nor2_1
Xhold3691 net7899 vssd1 vssd1 vccd1 vccd1 net4218 sky130_fd_sc_hd__dlygate4sd3_1
X_14952_ _08073_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
X_13903_ _07054_ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__or2_1
Xhold2990 net5913 vssd1 vssd1 vccd1 vccd1 net3517 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17671_ _01907_ _01909_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__and2_1
X_14883_ net4413 _08032_ net3775 vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__mux2_1
X_19410_ net3902 _03140_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nand2_2
X_16622_ net4188 net2898 _08111_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__mux2_1
X_13834_ _07003_ _06998_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19341_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__clkbuf_4
X_16553_ _09641_ _09642_ vssd1 vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__xor2_1
X_13765_ _06928_ _06929_ _06934_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__a21oi_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ net7314 net7013 _04309_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
X_15504_ _08588_ _08590_ _08598_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__a21bo_1
X_19272_ _03205_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__clkbuf_4
X_12716_ _05890_ _05893_ _05850_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__mux2_1
X_16484_ _09462_ _09574_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_169_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13696_ _06662_ _06673_ _06771_ _06796_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__or4_4
XFILLER_0_73_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18223_ _02440_ net4575 _02393_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
X_15435_ _08127_ _08142_ _08529_ _08338_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__o22a_1
X_12647_ _05797_ _05802_ net4147 _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15366_ _08460_ _08443_ _06121_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__a21o_1
X_18154_ net4567 net4461 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__or2_1
X_12578_ net4103 net4024 _05730_ net3996 net16 net19 vssd1 vssd1 vccd1 vccd1 _05758_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _10123_ _10125_ vssd1 vssd1 vccd1 vccd1 _10126_ sky130_fd_sc_hd__xor2_2
Xclkbuf_0__03843_ _03843_ vssd1 vssd1 vccd1 vccd1 clknet_0__03843_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14317_ _07467_ _07487_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__and2_4
X_11529_ _04679_ net1803 net4309 _04465_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__o22a_1
X_15297_ _08384_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__buf_2
XFILLER_0_145_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18085_ net4782 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__buf_4
Xhold307 net8203 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 net5202 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ _10055_ _10056_ vssd1 vssd1 vccd1 vccd1 _10057_ sky130_fd_sc_hd__nand2_1
X_14248_ _07413_ _07305_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__nor2_1
Xhold329 net5299 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14179_ _07345_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ net3270 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _00905_ vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17938_ _10327_ _08799_ _01693_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__nor3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _03435_ vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 _03816_ vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
X_17869_ _02104_ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor2_1
X_19608_ net1021 net4816 _03312_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20880_ _02757_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19539_ _08092_ _03386_ net1777 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__and3_2
XFILLER_0_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21501_ clknet_leaf_22_i_clk net1434 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21432_ clknet_leaf_40_i_clk net1645 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21363_ clknet_leaf_3_i_clk net4197 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20314_ net1356 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold830 _01268_ vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_21294_ clknet_leaf_34_i_clk net5422 vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold841 net6373 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold852 _00967_ vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20245_ _05673_ net4111 net4025 _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__and4_1
Xhold863 net6332 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _01274_ vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 net6268 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 net6336 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ net4416 _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or2_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2220 net7116 vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2231 net3439 vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2242 _01547_ vssd1 vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2253 net7364 vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2264 _04061_ vssd1 vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1530 _00753_ vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2275 _03571_ vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2286 net7392 vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1541 net4385 vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2297 net5650 vssd1 vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1552 net628 vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1563 _00690_ vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1574 net6821 vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ net2590 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__clkbuf_1
Xhold1585 _01362_ vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1596 net5545 vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11880_ net4058 net5912 net4107 net5205 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__o22ai_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_109 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_109/HI o_rgb[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_95_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10831_ net7492 net7514 _04227_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ _06719_ _06720_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ net2750 net6243 _04194_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _05676_ _05682_ net5 vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__mux2_1
X_13481_ _06392_ _06558_ _06561_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__o21a_1
X_10693_ _04104_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ _08312_ net8045 _08124_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__a21o_1
X_12432_ net4080 _05015_ _05021_ net3781 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _08240_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ net7725 net4956 _04845_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14102_ _07246_ _07247_ _07271_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__nand3_1
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11314_ _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__and2_2
X_15082_ _08175_ _08176_ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__nand2_2
XFILLER_0_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ _05276_ _05477_ _05479_ _04919_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _06576_ net3579 _06914_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__or3_1
X_18910_ net6357 net7143 _03014_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__mux2_1
X_11245_ net7258 net3005 _04445_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19890_ net6436 net3273 _03550_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18841_ net3937 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__clkbuf_1
X_11176_ net7391 net6156 _04412_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18772_ _02865_ net6046 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__or2_1
X_15984_ _09076_ _09078_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__xor2_1
X_17723_ _01940_ _01942_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14935_ net3943 _06239_ _08035_ net3926 net4661 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__o221a_1
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17654_ _01813_ _01806_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__or2b_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _07934_ net8362 vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__nor2_2
XFILLER_0_188_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16605_ _09692_ _09694_ vssd1 vssd1 vccd1 vccd1 _09695_ sky130_fd_sc_hd__xor2_2
XFILLER_0_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ _06986_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__xnor2_2
X_17585_ _01805_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14797_ _07864_ _07926_ _07944_ _07959_ net532 net7785 vssd1 vssd1 vccd1 vccd1 _07960_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19324_ net5276 _03250_ _03260_ _03259_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__o211a_1
X_16536_ _09624_ _09625_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__nor2_1
X_13748_ _06918_ _06916_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19255_ net6370 _03217_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__or2_1
X_16467_ _09555_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ _06838_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__xor2_1
Xhold7209 rbzero.color_sky\[1\] vssd1 vssd1 vccd1 vccd1 net7736 sky130_fd_sc_hd__dlygate4sd3_1
X_18206_ _02425_ net3669 _02393_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15418_ _08500_ _08501_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19186_ net6281 _03170_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__or2_1
X_16398_ _09487_ _09485_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6508 net2761 vssd1 vssd1 vccd1 vccd1 net7035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6519 _03011_ vssd1 vssd1 vccd1 vccd1 net7046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ net8039 _02358_ _02359_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__o21a_1
X_15349_ net8065 _06120_ _08133_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__or4_4
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5807 rbzero.spi_registers.new_texadd\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net6334
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5818 net1298 vssd1 vssd1 vccd1 vccd1 net6345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 net6035 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5829 rbzero.pov.spi_buffer\[26\] vssd1 vssd1 vccd1 vccd1 net6356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold115 net6071 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18068_ _02270_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__xnor2_1
Xhold126 net4425 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _03693_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net4804 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17019_ _08167_ _09351_ vssd1 vssd1 vccd1 vccd1 _10040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold159 net5018 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20030_ net3990 _03634_ _03615_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__o21ai_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21981_ net423 net2812 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ clknet_leaf_80_i_clk net4510 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ net4932 net6122 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20794_ _03960_ _03961_ _03959_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_187_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7721 rbzero.debug_overlay.vplaneY\[-8\] vssd1 vssd1 vccd1 vccd1 net8248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7732 rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 net8259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7743 net7799 vssd1 vssd1 vccd1 vccd1 net8270 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21415_ clknet_leaf_38_i_clk net5454 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7776 net1079 vssd1 vssd1 vccd1 vccd1 net8303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7787 net3388 vssd1 vssd1 vccd1 vccd1 net8314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7798 net3491 vssd1 vssd1 vccd1 vccd1 net8325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21346_ clknet_leaf_13_i_clk net5163 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold660 _01313_ vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
X_21277_ clknet_leaf_25_i_clk net4308 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold671 net6461 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11030_ net2736 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
Xhold682 net5483 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
X_20228_ net3678 net2468 _03709_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__mux2_1
Xhold693 net6181 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ _03728_ net7627 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or2_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2050 _01392_ vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2061 net5615 vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 _03411_ vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2083 net7468 vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _06151_ _06152_ _06154_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and4_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2094 _01489_ vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _01134_ vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 net6831 vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14720_ net7811 _07887_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__a21oi_1
Xhold1382 net6867 vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ gpout0.vpos\[5\] net4126 net4160 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__or3b_1
Xhold1393 net6775 vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _07805_ _07810_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__nand2_2
X_11863_ _04485_ _04653_ _04656_ _05048_ net4148 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__o221a_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ net6808 net7336 _04216_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
X_13602_ _06729_ _06726_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__nand2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17370_ _10310_ _10276_ vssd1 vssd1 vccd1 vccd1 _10388_ sky130_fd_sc_hd__or2b_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _04938_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14582_ _07413_ _07457_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__nor2_1
X_16321_ _08491_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10745_ net7031 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13533_ _06589_ _06590_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19040_ net3745 net3596 net3398 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
X_16252_ _06123_ net4913 vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__or2_1
X_13464_ _06492_ _06612_ _06613_ _06615_ _06564_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__a311o_1
X_10676_ net7151 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12415_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _04924_ vssd1 vssd1 vccd1 vccd1 _05600_
+ sky130_fd_sc_hd__mux2_1
X_15203_ _08297_ net2898 _08194_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__mux2_2
XFILLER_0_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16183_ _08221_ _08411_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13395_ _06398_ _06403_ _06528_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _05530_ _05531_ _04984_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__mux2_1
X_15134_ _08228_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03511_ clknet_0__03511_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03511_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19942_ net3060 net7455 _03572_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux2_1
X_15065_ _08147_ net7835 _08157_ _08159_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__a2bb2o_2
X_12277_ _05463_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _07138_ _07136_ _07135_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11228_ net7332 net6780 _04434_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19873_ net6649 net6357 _03539_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ net4062 _04102_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nor2_2
X_11159_ net7244 net2488 _04401_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18755_ _02865_ net3761 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nand2_1
X_15967_ _09061_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__clkbuf_4
X_17706_ _10390_ _01837_ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14918_ net4917 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__o21a_1
X_18686_ _02828_ _02832_ _02838_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__o21ai_2
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _08550_ _08560_ _08558_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17637_ _10163_ _09114_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14849_ _08005_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17568_ _08918_ _10211_ _01693_ _10346_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19307_ _03237_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__clkbuf_4
X_16519_ _09607_ _09608_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _10404_ _10405_ _10402_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7006 rbzero.pov.spi_buffer\[41\] vssd1 vssd1 vccd1 vccd1 net7533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7017 net1055 vssd1 vssd1 vccd1 vccd1 net7544 sky130_fd_sc_hd__dlygate4sd3_1
X_19238_ net6419 _03203_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__or2_1
Xhold7028 rbzero.pov.spi_buffer\[28\] vssd1 vssd1 vccd1 vccd1 net7555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7039 rbzero.pov.ready_buffer\[52\] vssd1 vssd1 vccd1 vccd1 net7566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6305 net1898 vssd1 vssd1 vccd1 vccd1 net6832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6316 rbzero.spi_registers.new_leak\[2\] vssd1 vssd1 vccd1 vccd1 net6843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6327 net2563 vssd1 vssd1 vccd1 vccd1 net6854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19169_ net6305 _03170_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__or2_1
Xhold6338 rbzero.tex_b1\[30\] vssd1 vssd1 vccd1 vccd1 net6865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5604 rbzero.spi_registers.new_texadd\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net6131
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6349 net2117 vssd1 vssd1 vccd1 vccd1 net6876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21200_ clknet_leaf_127_i_clk net2586 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5615 net1041 vssd1 vssd1 vccd1 vccd1 net6142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5626 _04161_ vssd1 vssd1 vccd1 vccd1 net6153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5637 net1080 vssd1 vssd1 vccd1 vccd1 net6164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4903 net1007 vssd1 vssd1 vccd1 vccd1 net5430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5648 rbzero.spi_registers.new_texadd\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net6175
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5659 rbzero.tex_r0\[54\] vssd1 vssd1 vccd1 vccd1 net6186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4914 _00879_ vssd1 vssd1 vccd1 vccd1 net5441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21131_ clknet_leaf_30_i_clk net3963 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_1
Xhold4925 net1122 vssd1 vssd1 vccd1 vccd1 net5452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4936 rbzero.spi_registers.vshift\[4\] vssd1 vssd1 vccd1 vccd1 net5463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4947 net1162 vssd1 vssd1 vccd1 vccd1 net5474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4958 _00881_ vssd1 vssd1 vccd1 vccd1 net5485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4969 net1253 vssd1 vssd1 vccd1 vccd1 net5496 sky130_fd_sc_hd__buf_1
X_21062_ clknet_leaf_68_i_clk _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20013_ net3339 _03607_ net4443 _03339_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21964_ net406 net1193 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ clknet_leaf_77_i_clk _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21895_ net337 net2284 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _09721_ clknet_1_0__leaf__05946_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__and2_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20777_ net1009 net5622 vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10530_ net2719 net7087 _04064_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7540 net1028 vssd1 vssd1 vccd1 vccd1 net8067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ net6888 net6902 _04031_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7551 rbzero.traced_texa\[10\] vssd1 vssd1 vccd1 vccd1 net8078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7562 _00518_ vssd1 vssd1 vccd1 vccd1 net8089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7573 net681 vssd1 vssd1 vccd1 vccd1 net8100 sky130_fd_sc_hd__dlygate4sd3_1
X_12200_ rbzero.tex_g1\[11\] rbzero.tex_g1\[10\] _04923_ vssd1 vssd1 vccd1 vccd1 _05387_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6850 net2488 vssd1 vssd1 vccd1 vccd1 net7377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7595 rbzero.traced_texa\[-3\] vssd1 vssd1 vccd1 vccd1 net8122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _06305_ _06338_ _06341_ _06346_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__a2111o_1
Xhold6861 rbzero.tex_b1\[59\] vssd1 vssd1 vccd1 vccd1 net7388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6872 net2471 vssd1 vssd1 vccd1 vccd1 net7399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6883 _03006_ vssd1 vssd1 vccd1 vccd1 net7410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ _04847_ _05318_ _04829_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__o21a_1
Xhold6894 net2765 vssd1 vssd1 vccd1 vccd1 net7421 sky130_fd_sc_hd__dlygate4sd3_1
X_21329_ clknet_leaf_12_i_clk net5063 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12062_ rbzero.tex_r1\[33\] rbzero.tex_r1\[32\] _05250_ vssd1 vssd1 vccd1 vccd1 _05251_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold490 net6127 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ net2254 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16870_ _09630_ _09889_ _09890_ vssd1 vssd1 vccd1 vccd1 _09892_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15821_ _08402_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__clkbuf_4
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18540_ _08103_ _06042_ _02711_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__or3_1
X_15752_ _08831_ _08845_ _08846_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__a21oi_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _06104_ net3893 _06039_ net4034 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__a22o_1
Xhold1190 _01352_ vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _07873_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__clkbuf_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _02634_ _02647_ _02649_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11915_ net3370 _05102_ _05103_ net2898 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a22o_1
X_15683_ _08773_ _08777_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__xnor2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ net4033 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__clkbuf_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _08799_ _09403_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14634_ _07796_ _07798_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__nor2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _05024_ _05034_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17353_ _10146_ _10244_ _10243_ vssd1 vssd1 vccd1 vccd1 _10372_ sky130_fd_sc_hd__a21oi_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11777_ _04942_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14565_ _07735_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16304_ _09394_ _09395_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10728_ net2748 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__clkbuf_1
X_13516_ _06505_ _06545_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__nand2_1
X_17284_ _10162_ _10172_ _10170_ vssd1 vssd1 vccd1 vccd1 _10303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14496_ _07658_ _07662_ _07664_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19023_ net1426 net4016 _03078_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16235_ _09326_ net5769 vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__nand2_1
X_10659_ net2156 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ _06589_ _06590_ _06607_ _06617_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__a211o_4
Xclkbuf_leaf_8_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16166_ _08389_ _08308_ _08309_ _08392_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__or4_1
X_13378_ _06531_ _06533_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nand2_4
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15117_ _08160_ _08168_ net8414 _08211_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__or4_1
X_12329_ _05233_ _05510_ _05514_ _05263_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a211o_1
XFILLER_0_181_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16097_ _09024_ _09046_ _09190_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3509 _00619_ vssd1 vssd1 vccd1 vccd1 net4036 sky130_fd_sc_hd__dlygate4sd3_1
X_15048_ _08139_ _08142_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19925_ net3228 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2808 _00931_ vssd1 vssd1 vccd1 vccd1 net3335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2819 net7511 vssd1 vssd1 vccd1 vccd1 net3346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19856_ net1752 net7498 _03528_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18807_ net3485 _02951_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__nor2_1
X_16999_ _09905_ _09906_ _09903_ vssd1 vssd1 vccd1 vccd1 _10020_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18738_ _02873_ _02886_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18669_ net4764 net8092 _02822_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__and3_1
X_20700_ _03878_ _03881_ _03882_ _03883_ net4984 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a32o_1
XFILLER_0_176_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21680_ clknet_leaf_114_i_clk net5748 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6102 net1745 vssd1 vssd1 vccd1 vccd1 net6629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6113 rbzero.tex_g0\[11\] vssd1 vssd1 vccd1 vccd1 net6640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6124 net1833 vssd1 vssd1 vccd1 vccd1 net6651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6135 _03524_ vssd1 vssd1 vccd1 vccd1 net6662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6146 net1730 vssd1 vssd1 vccd1 vccd1 net6673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5401 rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 net5928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6157 _03835_ vssd1 vssd1 vccd1 vccd1 net6684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5412 rbzero.spi_registers.got_new_sky vssd1 vssd1 vccd1 vccd1 net5939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5423 _00481_ vssd1 vssd1 vccd1 vccd1 net5950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6168 net1683 vssd1 vssd1 vccd1 vccd1 net6695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6179 rbzero.pov.ready_buffer\[18\] vssd1 vssd1 vccd1 vccd1 net6706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5434 net3141 vssd1 vssd1 vccd1 vccd1 net5961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5445 net3605 vssd1 vssd1 vccd1 vccd1 net5972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4700 rbzero.spi_registers.texadd1\[6\] vssd1 vssd1 vccd1 vccd1 net5227 sky130_fd_sc_hd__dlygate4sd3_1
X_22163_ clknet_leaf_94_i_clk net4854 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5456 _03784_ vssd1 vssd1 vccd1 vccd1 net5983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4711 net937 vssd1 vssd1 vccd1 vccd1 net5238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4722 _00876_ vssd1 vssd1 vccd1 vccd1 net5249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5467 net1733 vssd1 vssd1 vccd1 vccd1 net5994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4733 net758 vssd1 vssd1 vccd1 vccd1 net5260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5478 net2441 vssd1 vssd1 vccd1 vccd1 net6005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4744 rbzero.spi_registers.texadd3\[22\] vssd1 vssd1 vccd1 vccd1 net5271 sky130_fd_sc_hd__dlygate4sd3_1
X_21114_ clknet_leaf_105_i_clk net3829 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold5489 _02694_ vssd1 vssd1 vccd1 vccd1 net6016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4755 net974 vssd1 vssd1 vccd1 vccd1 net5282 sky130_fd_sc_hd__dlygate4sd3_1
X_22094_ net156 net3130 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
Xhold4766 _00794_ vssd1 vssd1 vccd1 vccd1 net5293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4777 net814 vssd1 vssd1 vccd1 vccd1 net5304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4788 rbzero.spi_registers.texadd2\[13\] vssd1 vssd1 vccd1 vccd1 net5315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21045_ clknet_leaf_59_i_clk _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4799 net963 vssd1 vssd1 vccd1 vccd1 net5326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21947_ net389 net3171 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ net3406 _04584_ _04502_ net1361 vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a211o_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05851_ net4068 net32 _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0__f__03514_ clknet_0__03514_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03514_
+ sky130_fd_sc_hd__clkbuf_16
X_21878_ net320 net2302 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11631_ _04814_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__or2_4
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ net4086 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__clkbuf_1
X_20473__217 clknet_1_0__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__inv_2
XFILLER_0_38_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14350_ _07519_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11562_ net4154 _04748_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10513_ _04030_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__clkbuf_4
X_13301_ _06438_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ _07449_ _07450_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ net4105 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7370 net4212 vssd1 vssd1 vccd1 vccd1 net7897 sky130_fd_sc_hd__dlygate4sd3_1
X_16020_ net8002 _08129_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__nand2_2
X_13232_ _06310_ _06402_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__xnor2_4
Xhold7381 rbzero.traced_texVinit\[7\] vssd1 vssd1 vccd1 vccd1 net7908 sky130_fd_sc_hd__dlygate4sd3_1
X_10444_ net4145 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__clkbuf_1
Xhold7392 net4429 vssd1 vssd1 vccd1 vccd1 net7919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6680 rbzero.tex_r0\[18\] vssd1 vssd1 vccd1 vccd1 net7207 sky130_fd_sc_hd__dlygate4sd3_1
X_13163_ _06273_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__xnor2_1
Xhold6691 net2777 vssd1 vssd1 vccd1 vccd1 net7218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _04943_ _05301_ _04947_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17971_ _02206_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__xnor2_1
Xhold5990 _03451_ vssd1 vssd1 vccd1 vccd1 net6517 sky130_fd_sc_hd__dlygate4sd3_1
X_13094_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__clkbuf_4
X_20367__122 clknet_1_1__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__inv_2
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19710_ net6207 net3631 _03456_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux2_1
X_16922_ _08309_ _08411_ vssd1 vssd1 vccd1 vccd1 _09944_ sky130_fd_sc_hd__nor2_1
X_12045_ rbzero.tex_r1\[31\] rbzero.tex_r1\[30\] _05220_ vssd1 vssd1 vccd1 vccd1 _05234_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19641_ net6697 net3738 _03441_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
X_16853_ net4581 net4397 vssd1 vssd1 vccd1 vccd1 _09876_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15804_ _08897_ _08898_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19572_ net5613 net4016 _03403_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__mux2_1
X_16784_ net4569 net4485 vssd1 vssd1 vccd1 vccd1 _09814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _06719_ _06695_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__or2_1
X_18523_ net8258 _02683_ _02681_ net8257 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__o211a_1
X_15735_ _08793_ _08795_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12947_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__clkbuf_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _02610_ _02614_ _02632_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a21o_1
X_15666_ _08759_ _08760_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__nor2b_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _06029_ _06052_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17405_ _10421_ _10422_ vssd1 vssd1 vccd1 vccd1 _10423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07454_ _07509_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__and2_1
X_11829_ net4271 net4335 net4259 vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__nand3_1
X_18385_ _02559_ net8049 net4785 net3514 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a31o_1
X_15597_ _08308_ _08309_ _08329_ _08691_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__or4_4
XFILLER_0_173_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _10345_ _10354_ vssd1 vssd1 vccd1 vccd1 _10355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14548_ _07711_ _07717_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17267_ _10283_ _10284_ vssd1 vssd1 vccd1 vccd1 _10286_ sky130_fd_sc_hd__and2_1
X_14479_ _07625_ _07648_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19006_ net7510 net3345 _02992_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
X_16218_ _09271_ _09310_ vssd1 vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ _10208_ _10217_ vssd1 vssd1 vccd1 vccd1 _10218_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4007 net7857 vssd1 vssd1 vccd1 vccd1 net4534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16149_ _09226_ _09241_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__xor2_2
Xhold4018 net3383 vssd1 vssd1 vccd1 vccd1 net4545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4029 _01227_ vssd1 vssd1 vccd1 vccd1 net4556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3306 net7982 vssd1 vssd1 vccd1 vccd1 net3833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3317 _03422_ vssd1 vssd1 vccd1 vccd1 net3844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3328 net7974 vssd1 vssd1 vccd1 vccd1 net3855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3339 net7628 vssd1 vssd1 vccd1 vccd1 net3866 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2605 net7462 vssd1 vssd1 vccd1 vccd1 net3132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2616 _00597_ vssd1 vssd1 vccd1 vccd1 net3143 sky130_fd_sc_hd__dlygate4sd3_1
X_19908_ net3167 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
Xhold2627 _01417_ vssd1 vssd1 vccd1 vccd1 net3154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2638 _01335_ vssd1 vssd1 vccd1 vccd1 net3165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 net7436 vssd1 vssd1 vccd1 vccd1 net3176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 _01442_ vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03508_ _03508_ vssd1 vssd1 vccd1 vccd1 clknet_0__03508_ sky130_fd_sc_hd__clkbuf_16
Xhold1915 _03350_ vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1926 net7032 vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_19839_ net2312 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__clkbuf_4
Xhold1937 _01408_ vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1948 net5623 vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1959 _03021_ vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21801_ net243 net2666 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21732_ clknet_leaf_96_i_clk net3568 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21663_ clknet_leaf_23_i_clk net3161 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21594_ net228 net625 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5220 _01167_ vssd1 vssd1 vccd1 vccd1 net5747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5231 rbzero.pov.ready_buffer\[58\] vssd1 vssd1 vccd1 vccd1 net5758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5242 _09327_ vssd1 vssd1 vccd1 vccd1 net5769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5253 net8218 vssd1 vssd1 vccd1 vccd1 net5780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5264 net5906 vssd1 vssd1 vccd1 vccd1 net5791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5275 net1252 vssd1 vssd1 vccd1 vccd1 net5802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4530 net689 vssd1 vssd1 vccd1 vccd1 net5057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5286 _03066_ vssd1 vssd1 vccd1 vccd1 net5813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4541 rbzero.spi_registers.texadd2\[21\] vssd1 vssd1 vccd1 vccd1 net5068 sky130_fd_sc_hd__dlygate4sd3_1
X_22146_ clknet_leaf_81_i_clk _01633_ vssd1 vssd1 vccd1 vccd1 reg_vsync sky130_fd_sc_hd__dfxtp_1
Xhold5297 _00598_ vssd1 vssd1 vccd1 vccd1 net5824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4552 net702 vssd1 vssd1 vccd1 vccd1 net5079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4563 _00830_ vssd1 vssd1 vccd1 vccd1 net5090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4574 net742 vssd1 vssd1 vccd1 vccd1 net5101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4585 rbzero.spi_registers.texadd3\[4\] vssd1 vssd1 vccd1 vccd1 net5112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3840 _00774_ vssd1 vssd1 vccd1 vccd1 net4367 sky130_fd_sc_hd__dlygate4sd3_1
X_22077_ net519 net2799 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold4596 net732 vssd1 vssd1 vccd1 vccd1 net5123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3851 net7851 vssd1 vssd1 vccd1 vccd1 net4378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3862 net8056 vssd1 vssd1 vccd1 vccd1 net4389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3873 net7830 vssd1 vssd1 vccd1 vccd1 net4400 sky130_fd_sc_hd__dlygate4sd3_1
X_21028_ clknet_leaf_53_i_clk net4249 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3884 net1058 vssd1 vssd1 vccd1 vccd1 net4411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3895 net1205 vssd1 vssd1 vccd1 vccd1 net4422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13850_ _06976_ net548 vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ net7744 net6046 vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__nand2_2
X_10993_ net2845 net51 _04238_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
X_13781_ _06926_ _06951_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__xnor2_2
X_15520_ _08611_ _08614_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__or2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ net4149 net4141 net4164 net4173 _05901_ net37 vssd1 vssd1 vccd1 vccd1 _05909_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _08338_ _08529_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__nor3_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_73_i_clk clknet_4_12__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _06914_ _07390_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nor2_1
X_11614_ _04766_ _04768_ _04765_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a21oi_1
X_18170_ _02394_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__clkbuf_1
X_15382_ _08427_ _08428_ net8042 _08475_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ _05756_ _05762_ _05767_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _10057_ _10024_ vssd1 vssd1 vccd1 vccd1 _10141_ sky130_fd_sc_hd__or2b_1
XFILLER_0_167_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ _07502_ _07503_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__or2b_1
XFILLER_0_53_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11545_ net4095 _04731_ _04733_ net4357 _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__o221a_1
X_17052_ _09943_ _09944_ vssd1 vssd1 vccd1 vccd1 _10073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14264_ _07237_ _07354_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__or2b_1
X_11476_ net7562 _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__or2_2
XFILLER_0_151_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16003_ _09089_ net7766 _09097_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__a21oi_1
X_13215_ _06308_ _06310_ _06367_ _06381_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a41o_1
XFILLER_0_123_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _07284_ _07360_ _07365_ net5902 vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13146_ _06281_ _06312_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__xor2_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _02075_ _02089_ _02190_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a21bo_1
X_13077_ net5531 net5605 _06244_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__o21a_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16905_ _09650_ _09895_ _09926_ vssd1 vssd1 vccd1 vccd1 _09927_ sky130_fd_sc_hd__a21o_1
X_12028_ _05215_ _05216_ _05206_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17885_ _02121_ _02122_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19624_ net6297 net3863 _03430_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__mux2_1
X_16836_ _09859_ net3798 vssd1 vssd1 vccd1 vccd1 _09861_ sky130_fd_sc_hd__or2b_1
XFILLER_0_189_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19555_ net1880 net1777 vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nand2_1
X_16767_ net3805 _09798_ vssd1 vssd1 vccd1 vccd1 _09799_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13979_ _07100_ _07131_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nand2_1
X_18506_ _02626_ net6015 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15718_ _08805_ _08807_ _08806_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__a21o_1
X_19486_ net6012 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20421__171 clknet_1_1__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__inv_2
X_16698_ net864 _09745_ _09746_ net7999 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18437_ _02617_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02618_
+ sky130_fd_sc_hd__nand2_1
X_15649_ _08674_ _08728_ _08740_ _08741_ _08743_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__a32o_1
X_19781__60 clknet_1_0__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18368_ net3493 rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1 vccd1 _02554_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_161_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17319_ _10223_ _10224_ vssd1 vssd1 vccd1 vccd1 _10338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ net6339 net3738 _02493_ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330_ net6182 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20261_ _09721_ _03798_ net4112 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22000_ net442 net2452 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3103 net8395 vssd1 vssd1 vccd1 vccd1 net3630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20192_ net2079 _03743_ net4502 _03732_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3114 net6037 vssd1 vssd1 vccd1 vccd1 net3641 sky130_fd_sc_hd__buf_2
Xhold3125 _03321_ vssd1 vssd1 vccd1 vccd1 net3652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3136 _03756_ vssd1 vssd1 vccd1 vccd1 net3663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3147 net7614 vssd1 vssd1 vccd1 vccd1 net3674 sky130_fd_sc_hd__clkbuf_2
Xhold2402 _01151_ vssd1 vssd1 vccd1 vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2413 net3059 vssd1 vssd1 vccd1 vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3158 _01180_ vssd1 vssd1 vccd1 vccd1 net3685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 _04135_ vssd1 vssd1 vccd1 vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3169 _02988_ vssd1 vssd1 vccd1 vccd1 net3696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2435 net7458 vssd1 vssd1 vccd1 vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1701 _01466_ vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2446 rbzero.pov.spi_buffer\[43\] vssd1 vssd1 vccd1 vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1712 net1988 vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2457 net7267 vssd1 vssd1 vccd1 vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 _01512_ vssd1 vssd1 vccd1 vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1723 net5644 vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _01574_ vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2479 _04451_ vssd1 vssd1 vccd1 vccd1 net3006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1745 _04089_ vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1756 net7168 vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1767 net7148 vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1778 _01532_ vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
X_20504__246 clknet_1_1__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__inv_2
Xhold1789 _04452_ vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21715_ clknet_leaf_127_i_clk net3693 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21646_ clknet_leaf_117_i_clk net3136 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21577_ net211 net2656 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_60 _05794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_71 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_82 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ rbzero.spi_registers.texadd3\[7\] rbzero.spi_registers.texadd1\[7\] rbzero.spi_registers.texadd0\[7\]
+ rbzero.spi_registers.texadd2\[7\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux4_2
XANTENNA_93 net8012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ _04102_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__clkbuf_8
X_20585__318 clknet_1_0__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__inv_2
XFILLER_0_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5050 rbzero.tex_r0\[48\] vssd1 vssd1 vccd1 vccd1 net5577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5061 net2884 vssd1 vssd1 vccd1 vccd1 net5588 sky130_fd_sc_hd__dlygate4sd3_1
X_13000_ net3749 _06174_ net4506 _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_162_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ net6942 net2744 _04412_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__mux2_1
Xhold5072 _04060_ vssd1 vssd1 vccd1 vccd1 net5599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5083 _01621_ vssd1 vssd1 vccd1 vccd1 net5610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5094 rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 net5621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4360 net789 vssd1 vssd1 vccd1 vccd1 net4887 sky130_fd_sc_hd__dlygate4sd3_1
X_22129_ clknet_leaf_53_i_clk net5694 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold4371 rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 net4898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4382 _09602_ vssd1 vssd1 vccd1 vccd1 net4909 sky130_fd_sc_hd__buf_1
XFILLER_0_203_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4393 net3887 vssd1 vssd1 vccd1 vccd1 net4920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3670 net841 vssd1 vssd1 vccd1 vccd1 net4197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3681 net8136 vssd1 vssd1 vccd1 vccd1 net4208 sky130_fd_sc_hd__dlygate4sd3_1
X_14951_ net4630 _07929_ _08068_ vssd1 vssd1 vccd1 vccd1 _08073_ sky130_fd_sc_hd__mux2_1
Xhold3692 net7901 vssd1 vssd1 vccd1 vccd1 net4219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13902_ _07051_ _07053_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__nor2_1
X_17670_ _01907_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__nor2_1
Xhold2980 net7797 vssd1 vssd1 vccd1 vccd1 net3507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2991 _00478_ vssd1 vssd1 vccd1 vccd1 net3518 sky130_fd_sc_hd__dlygate4sd3_1
X_14882_ _07869_ net8370 _07996_ vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__nor3_1
X_16621_ _09589_ _09710_ vssd1 vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_134_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13833_ _06998_ _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__nand2b_1
X_20479__223 clknet_1_1__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__inv_2
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19340_ net1020 _03140_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__nand2_2
X_16552_ _08326_ _08411_ vssd1 vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13764_ _06928_ _06929_ _06934_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__and3_1
X_10976_ _04264_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__buf_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _08591_ _08587_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19271_ net2075 _03202_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__or2_1
X_12715_ _05891_ _05892_ _05862_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__mux2_1
X_16483_ _09464_ _09573_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__xnor2_4
X_13695_ _06744_ _06745_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18222_ _02438_ _02439_ _01953_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ _08528_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12646_ net43 _05798_ _05818_ net44 _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ _02379_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__clkbuf_1
X_15365_ net3531 _08133_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ net4111 _05673_ net4071 net4092 _05749_ net18 vssd1 vssd1 vccd1 vccd1 _05757_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17104_ _09893_ _09999_ _10124_ vssd1 vssd1 vccd1 vccd1 _10125_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_29_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03842_ _03842_ vssd1 vssd1 vccd1 vccd1 clknet_0__03842_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _07464_ _07465_ _07466_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__a21o_1
X_11528_ net4309 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__inv_2
X_18084_ net4646 _09413_ _06239_ net4781 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__o211ai_1
X_15296_ _08241_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold308 net8020 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17035_ _10025_ _10026_ _10054_ vssd1 vssd1 vccd1 vccd1 _10056_ sky130_fd_sc_hd__nand3_1
Xhold319 net5355 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14247_ net569 _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20451__197 clknet_1_1__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__inv_2
X_11459_ _04465_ _04612_ _04622_ _04650_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14178_ _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__xor2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ net4513 net6015 _06296_ _06299_ _06297_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a221o_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ net7449 net7536 _03058_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 net5815 vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ _10327_ _08799_ _01693_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a21o_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1019 _00970_ vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17868_ _09915_ _09612_ _01973_ _02105_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o31a_1
XFILLER_0_205_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19607_ net4815 _03363_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__nand2_1
X_16819_ net4633 _09843_ _09845_ vssd1 vssd1 vccd1 vccd1 _09846_ sky130_fd_sc_hd__a21o_1
X_17799_ _02035_ _02036_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19538_ net3906 _02948_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19469_ net1493 net5996 _03345_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21500_ clknet_leaf_3_i_clk net1651 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21431_ clknet_leaf_40_i_clk net2449 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7914 _06571_ vssd1 vssd1 vccd1 vccd1 net8441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21362_ clknet_leaf_3_i_clk net5135 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20313_ net6372 net3738 _03825_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21293_ clknet_leaf_34_i_clk net5418 vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold820 _03462_ vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 net3272 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 net6375 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 net6338 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
X_20244_ net4103 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold864 _00595_ vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 net5561 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 _01278_ vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _00574_ vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
X_20175_ _03710_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2210 _01324_ vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2221 _04178_ vssd1 vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2232 _03042_ vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2243 net7528 vssd1 vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2254 _04044_ vssd1 vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20428__177 clknet_1_1__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__inv_2
Xhold2265 _01570_ vssd1 vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1520 _03111_ vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1531 net5617 vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__buf_1
Xhold2276 _01135_ vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2287 _04413_ vssd1 vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1542 net7177 vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1553 _03009_ vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2298 _01306_ vssd1 vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1564 net6702 vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 net6823 vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1586 net7100 vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1597 _01479_ vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10830_ net6213 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10761_ net2289 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _05679_ _05681_ _05649_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__mux2_1
X_10692_ net2188 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__clkbuf_1
X_13480_ _06557_ _06647_ _06650_ _06605_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a211o_1
X_19760__41 clknet_1_0__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_0_168_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12431_ _04818_ _05590_ _05598_ _04821_ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a311o_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21629_ clknet_leaf_129_i_clk net3304 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15150_ _08226_ _08227_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ _05547_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14101_ _07246_ _07247_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11313_ net7748 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__buf_4
X_12293_ _04976_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__or2_1
X_15081_ net3489 net3417 net5859 vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__o21ai_1
X_11244_ net6934 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__clkbuf_1
X_14032_ _07114_ _07162_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net2814 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
X_18840_ _02969_ net3936 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4190 net694 vssd1 vssd1 vccd1 vccd1 net4717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18771_ _02866_ net6046 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ _08354_ _08655_ _09077_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__a21boi_2
X_17722_ _01958_ _01959_ _09845_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a21o_1
X_14934_ net7821 _06237_ _04482_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__o21a_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _01807_ _01812_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__nand2_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _07877_ _07978_ net7846 vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__mux2_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16604_ _09533_ _09558_ _09693_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_203_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13816_ _06945_ _06947_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17584_ _01823_ _01824_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__nor2_1
X_14796_ _07804_ _07853_ _07818_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ net1718 _03251_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16535_ _09478_ _09490_ _09488_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ _06683_ _06737_ _06705_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10959_ net6778 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19254_ net5424 _03216_ _03220_ _03219_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__o211a_1
X_16466_ _09408_ _09425_ _09556_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13678_ _06841_ _06848_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18205_ _09809_ _02424_ _01729_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__o21ai_1
X_15417_ _08508_ _08510_ _08511_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12629_ _05797_ net24 _05801_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__nand4_1
X_19185_ net5256 _03168_ _03179_ _03176_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__o211a_1
X_16397_ _09485_ _09487_ vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6509 _04169_ vssd1 vssd1 vccd1 vccd1 net7036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18136_ _02364_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__clkbuf_1
X_15348_ net3453 _08438_ _08439_ _08442_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__a31o_4
X_20533__272 clknet_1_1__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__inv_2
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5808 net1422 vssd1 vssd1 vccd1 vccd1 net6335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5819 rbzero.spi_registers.new_texadd\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net6346
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 _01413_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
X_18067_ _02297_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__xnor2_1
Xhold116 net6073 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
X_20664__10 clknet_1_1__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
X_15279_ _08372_ _08373_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__or2_4
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold127 net8297 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net4437 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _09912_ _09913_ _09911_ vssd1 vssd1 vccd1 vccd1 _10039_ sky130_fd_sc_hd__a21bo_1
Xhold149 net7507 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ net3121 net6687 net2874 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ net422 net2749 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
X_20931_ clknet_leaf_60_i_clk net4549 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20862_ net4932 net63 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20793_ _03959_ _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7700 net3536 vssd1 vssd1 vccd1 vccd1 net8227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7711 _08045_ vssd1 vssd1 vccd1 vccd1 net8238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7722 _04013_ vssd1 vssd1 vccd1 vccd1 net8249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7733 _02700_ vssd1 vssd1 vccd1 vccd1 net8260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21414_ clknet_leaf_52_i_clk net5466 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7788 rbzero.texu_hot\[5\] vssd1 vssd1 vccd1 vccd1 net8315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21345_ clknet_leaf_13_i_clk net4200 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7799 rbzero.wall_tracer.stepDistX\[-8\] vssd1 vssd1 vccd1 vccd1 net8326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21276_ clknet_leaf_25_i_clk net4326 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 _03150_ vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 net6226 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold672 _01067_ vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold683 net5485 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
X_20227_ net6693 _03706_ net4687 _03765_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 _01276_ vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
X_20158_ rbzero.debug_overlay.facingY\[-7\] net3289 _03723_ vssd1 vssd1 vccd1 vccd1
+ _03733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2040 _04213_ vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2051 rbzero.tex_b1\[8\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2062 net7278 vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20089_ net3326 _08299_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__nand2_1
X_12980_ net4309 _06068_ net3965 _04722_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__o221a_1
Xhold2073 _00952_ vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2084 net7370 vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2095 net2734 vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1350 _00665_ vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 net6865 vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1372 _01050_ vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _04664_ _04660_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__nor2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 net6869 vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 net6777 vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14650_ net7795 vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__buf_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11862_ net4147 net4066 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nor2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _06693_ _06771_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__or2_1
X_10813_ net7173 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__clkbuf_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14581_ _07072_ _07327_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__or2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04977_ _04980_ _04982_ _04919_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__o211a_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16320_ _08905_ _09411_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__clkbuf_4
X_10744_ net2999 net7029 _04182_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16251_ net8275 _08129_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__nand2_1
X_13463_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__clkbuf_8
X_10675_ net7149 net2635 _04149_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15202_ _08295_ _08296_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__and2_1
X_12414_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _05369_ vssd1 vssd1 vccd1 vccd1 _05599_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ _08241_ _08403_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13394_ _06389_ _06401_ _06549_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _08226_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__or2_1
X_12345_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _04913_ vssd1 vssd1 vccd1 vccd1 _05531_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03510_ clknet_0__03510_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03510_
+ sky130_fd_sc_hd__clkbuf_16
X_19941_ net2861 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
X_15064_ _08156_ _08158_ _08148_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__o21a_1
X_12276_ reg_rgb\[15\] _05462_ _05054_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__mux2_4
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14015_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__inv_2
X_11227_ net6770 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__clkbuf_1
X_19872_ net3174 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
X_18823_ _02947_ net3486 vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__and2_1
X_11158_ net6105 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11089_ net7308 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
X_15966_ _08128_ _09060_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__or2_1
X_20563__298 clknet_1_0__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__inv_2
X_18754_ net5842 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__clkbuf_1
X_17705_ _01835_ _01836_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__nor2_1
X_14917_ net4669 _08050_ _08052_ net4526 net4585 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__o221a_1
X_15897_ _08656_ _08762_ _08989_ _08991_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__a2bb2o_4
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18685_ _02828_ _02832_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__or3_1
XFILLER_0_188_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17636_ _01874_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__xnor2_1
X_14848_ net4430 _08004_ _07976_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17567_ _08918_ _01693_ _10346_ _10211_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_59_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14779_ _07851_ _07855_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _08611_ _09470_ _09472_ _09468_ vssd1 vssd1 vccd1 vccd1 _09608_ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19306_ _03235_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__buf_4
X_17498_ _10427_ _10393_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16449_ _09419_ _09296_ _06123_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__a21o_2
Xhold7007 net3166 vssd1 vssd1 vccd1 vccd1 net7534 sky130_fd_sc_hd__dlygate4sd3_1
X_19237_ net5097 _03201_ _03210_ _03206_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7018 _03024_ vssd1 vssd1 vccd1 vccd1 net7545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7029 net3179 vssd1 vssd1 vccd1 vccd1 net7556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6306 rbzero.tex_r0\[12\] vssd1 vssd1 vccd1 vccd1 net6833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19168_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6317 net2256 vssd1 vssd1 vccd1 vccd1 net6844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6328 _04279_ vssd1 vssd1 vccd1 vccd1 net6855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6339 net1888 vssd1 vssd1 vccd1 vccd1 net6866 sky130_fd_sc_hd__dlygate4sd3_1
X_18119_ _02349_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__clkbuf_1
Xhold5605 net2137 vssd1 vssd1 vccd1 vccd1 net6132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5616 rbzero.tex_r1\[10\] vssd1 vssd1 vccd1 vccd1 net6143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5627 net1090 vssd1 vssd1 vccd1 vccd1 net6154 sky130_fd_sc_hd__dlygate4sd3_1
X_19099_ _09721_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__clkbuf_4
Xhold5638 _04272_ vssd1 vssd1 vccd1 vccd1 net6165 sky130_fd_sc_hd__dlygate4sd3_1
X_21130_ clknet_leaf_32_i_clk net3449 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4904 rbzero.map_overlay.i_mapdx\[5\] vssd1 vssd1 vccd1 vccd1 net5431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5649 net1386 vssd1 vssd1 vccd1 vccd1 net6176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4915 net1051 vssd1 vssd1 vccd1 vccd1 net5442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4926 _00902_ vssd1 vssd1 vccd1 vccd1 net5453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4937 net1156 vssd1 vssd1 vccd1 vccd1 net5464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4948 rbzero.pov.ready_buffer\[21\] vssd1 vssd1 vccd1 vccd1 net5475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4959 net1210 vssd1 vssd1 vccd1 vccd1 net5486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21061_ clknet_leaf_68_i_clk _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20012_ _03609_ net4442 vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21963_ net405 net2752 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ clknet_leaf_65_i_clk _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21894_ net336 net3072 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _03999_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20776_ _03878_ _03945_ _03947_ _03883_ net5488 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7530 net4389 vssd1 vssd1 vccd1 vccd1 net8057 sky130_fd_sc_hd__dlygate4sd3_1
X_10460_ net6583 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__clkbuf_1
Xhold7541 net8467 vssd1 vssd1 vccd1 vccd1 net8068 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7552 net850 vssd1 vssd1 vccd1 vccd1 net8079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7563 net4291 vssd1 vssd1 vccd1 vccd1 net8090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7574 _01652_ vssd1 vssd1 vccd1 vccd1 net8101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7585 _02845_ vssd1 vssd1 vccd1 vccd1 net8112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6840 net2411 vssd1 vssd1 vccd1 vccd1 net7367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6851 _04406_ vssd1 vssd1 vccd1 vccd1 net7378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7596 net896 vssd1 vssd1 vccd1 vccd1 net8123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6862 net2285 vssd1 vssd1 vccd1 vccd1 net7389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6873 rbzero.tex_b1\[39\] vssd1 vssd1 vccd1 vccd1 net7400 sky130_fd_sc_hd__dlygate4sd3_1
X_12130_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _04950_ vssd1 vssd1 vccd1 vccd1 _05318_
+ sky130_fd_sc_hd__mux2_1
Xhold6884 net2944 vssd1 vssd1 vccd1 vccd1 net7411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6895 rbzero.tex_g0\[37\] vssd1 vssd1 vccd1 vccd1 net7422 sky130_fd_sc_hd__dlygate4sd3_1
X_21328_ clknet_leaf_47_i_clk net5079 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__clkbuf_8
X_21259_ clknet_leaf_22_i_clk net3772 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold480 net5429 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold491 net6129 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11012_ net7157 net7240 _04320_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__mux2_1
X_15820_ _08896_ _08913_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__xor2_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _08832_ _08844_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__nor2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ net3960 _06061_ net3848 net3965 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a22o_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 _03537_ vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ net4381 _07870_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__mux2_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 net6602 vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _02630_ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__xnor2_1
X_11914_ _04684_ _05079_ _05098_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__nor3_4
X_15682_ _08775_ _08776_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__nand2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ net4053 net4641 _06048_ net3552 _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__a221o_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _10437_ _10438_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__and2_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14633_ _07789_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__xnor2_4
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ net3781 _05015_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__nor2_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _10275_ _10370_ vssd1 vssd1 vccd1 vccd1 _10371_ sky130_fd_sc_hd__xnor2_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _07308_ _07457_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__or2_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _04941_ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__nor2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _08509_ _08403_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ _06669_ _06685_ _06493_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__mux2_1
X_17283_ _10292_ _10301_ vssd1 vssd1 vccd1 vccd1 _10302_ sky130_fd_sc_hd__xnor2_1
X_10727_ net6818 net7117 _04097_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14495_ _07630_ _07643_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__xnor2_1
X_19022_ net4077 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ net7781 net5768 _08111_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__mux2_1
X_13446_ _06611_ _06616_ _06540_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__a21oi_2
X_10658_ net7299 net7224 _04138_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ _09256_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13377_ _06451_ _06452_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__xor2_1
X_10589_ net49 net2947 _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15116_ _08210_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__clkbuf_4
X_12328_ _04911_ _05511_ _05513_ _04919_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16096_ _09043_ _09045_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__and2b_1
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ _08141_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__clkbuf_4
X_19924_ net3227 net5710 _03572_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__mux2_1
X_12259_ rbzero.tex_g1\[59\] rbzero.tex_g1\[58\] _04968_ vssd1 vssd1 vccd1 vccd1 _05446_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2809 net4185 vssd1 vssd1 vccd1 vccd1 net3336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20645__373 clknet_1_1__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__inv_2
X_19855_ net3064 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
X_18806_ net4832 _02948_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a21oi_2
X_20344__101 clknet_1_0__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__inv_2
XFILLER_0_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _09929_ _09894_ vssd1 vssd1 vccd1 vccd1 _10019_ sky130_fd_sc_hd__or2b_1
X_18737_ _02869_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__xnor2_1
X_15949_ _08453_ _08468_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18668_ net4764 net8092 _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17619_ _01804_ _01781_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18599_ net4528 net4848 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20561_ clknet_1_0__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__buf_1
XFILLER_0_55_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20390__143 clknet_1_0__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__inv_2
Xhold6103 _03477_ vssd1 vssd1 vccd1 vccd1 net6630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6114 net1715 vssd1 vssd1 vccd1 vccd1 net6641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6125 _04140_ vssd1 vssd1 vccd1 vccd1 net6652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6136 net1580 vssd1 vssd1 vccd1 vccd1 net6663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6147 _04431_ vssd1 vssd1 vccd1 vccd1 net6674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5402 net3417 vssd1 vssd1 vccd1 vccd1 net5929 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6158 net2221 vssd1 vssd1 vccd1 vccd1 net6685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5413 net3902 vssd1 vssd1 vccd1 vccd1 net5940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6169 rbzero.spi_registers.new_texadd\[0\]\[14\] vssd1 vssd1 vccd1 vccd1 net6696
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5424 net4090 vssd1 vssd1 vccd1 vccd1 net5951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5435 _02538_ vssd1 vssd1 vccd1 vccd1 net5962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22162_ clknet_leaf_94_i_clk net4889 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5446 rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 net5973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4701 net852 vssd1 vssd1 vccd1 vccd1 net5228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4712 rbzero.spi_registers.texadd0\[8\] vssd1 vssd1 vccd1 vccd1 net5239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5457 _03785_ vssd1 vssd1 vccd1 vccd1 net5984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5468 rbzero.spi_registers.new_sky\[2\] vssd1 vssd1 vccd1 vccd1 net5995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4723 net819 vssd1 vssd1 vccd1 vccd1 net5250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5479 rbzero.spi_registers.new_sky\[5\] vssd1 vssd1 vccd1 vccd1 net6006 sky130_fd_sc_hd__dlygate4sd3_1
X_21113_ clknet_leaf_105_i_clk net4787 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold4734 _00841_ vssd1 vssd1 vccd1 vccd1 net5261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4745 net982 vssd1 vssd1 vccd1 vccd1 net5272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22093_ net155 net2986 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
Xhold4756 rbzero.spi_registers.texadd1\[16\] vssd1 vssd1 vccd1 vccd1 net5283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4767 net912 vssd1 vssd1 vccd1 vccd1 net5294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4778 _00853_ vssd1 vssd1 vccd1 vccd1 net5305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21044_ clknet_leaf_61_i_clk _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4789 net874 vssd1 vssd1 vccd1 vccd1 net5316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21946_ net388 net1085 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03513_ clknet_0__03513_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03513_
+ sky130_fd_sc_hd__clkbuf_16
X_21877_ net319 net2484 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11630_ _04805_ _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__xnor2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20828_ _08038_ net4085 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__and2_1
X_11561_ _04691_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__or2_1
X_20759_ _03930_ _03931_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13300_ _06399_ _06470_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nor2_1
X_10512_ net6261 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _07449_ _07450_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__nor2_1
X_11492_ net4138 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7360 rbzero.traced_texVinit\[3\] vssd1 vssd1 vccd1 vccd1 net7887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13231_ _06367_ _06381_ _06385_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a21oi_2
Xhold7371 net1075 vssd1 vssd1 vccd1 vccd1 net7898 sky130_fd_sc_hd__dlygate4sd3_1
X_10443_ net4132 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__clkbuf_1
Xhold7382 net4223 vssd1 vssd1 vccd1 vccd1 net7909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6670 _04343_ vssd1 vssd1 vccd1 vccd1 net7197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13162_ _06274_ _06275_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__and2b_1
Xhold6681 net2450 vssd1 vssd1 vccd1 vccd1 net7208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6692 rbzero.tex_r0\[22\] vssd1 vssd1 vccd1 vccd1 net7219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _04951_ vssd1 vssd1 vccd1 vccd1 _05301_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5980 _04299_ vssd1 vssd1 vccd1 vccd1 net6507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17970_ _01760_ _09114_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__nor2_1
Xhold5991 net1571 vssd1 vssd1 vccd1 vccd1 net6518 sky130_fd_sc_hd__dlygate4sd3_1
X_13093_ net8217 _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _04988_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__buf_4
X_16921_ _08326_ _09025_ vssd1 vssd1 vccd1 vccd1 _09943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ net1406 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__clkbuf_1
X_16852_ net3799 _09867_ vssd1 vssd1 vccd1 vccd1 _09875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15803_ _08402_ _08328_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16783_ _09804_ _09805_ _09806_ vssd1 vssd1 vccd1 vccd1 _09813_ sky130_fd_sc_hd__o21a_1
X_19571_ net3003 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13995_ _07111_ _07112_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15734_ _08826_ _08828_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__nor2_1
X_18522_ _02695_ _02696_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12946_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15665_ _08756_ _08758_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__nand2_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _02610_ _02614_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nand3_1
X_12877_ _06029_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _10419_ _10420_ vssd1 vssd1 vccd1 vccd1 _10422_ sky130_fd_sc_hd__and2_1
X_14616_ _07508_ _07559_ _07784_ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__a22oi_4
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ net3781 _05015_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__nand2_1
X_18384_ _04490_ _02567_ _02568_ _09736_ rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15596_ _08341_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__clkbuf_4
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _10352_ _10353_ vssd1 vssd1 vccd1 vccd1 _10354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _07711_ _07717_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _04921_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ _10283_ _10284_ vssd1 vssd1 vccd1 vccd1 _10285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14478_ _07625_ _07648_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__xor2_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16217_ _09307_ _09309_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__xor2_2
X_19005_ net3016 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13429_ _06530_ _06532_ _06522_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17197_ _10210_ _10216_ vssd1 vssd1 vccd1 vccd1 _10217_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ _09239_ _09240_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__xor2_2
Xhold4008 net3725 vssd1 vssd1 vccd1 vccd1 net4535 sky130_fd_sc_hd__clkbuf_2
Xhold4019 net7987 vssd1 vssd1 vccd1 vccd1 net4546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16079_ _08010_ _08017_ net565 _08021_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__o31a_1
Xhold3307 net7993 vssd1 vssd1 vccd1 vccd1 net3834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3318 _00962_ vssd1 vssd1 vccd1 vccd1 net3845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3329 net7976 vssd1 vssd1 vccd1 vccd1 net3856 sky130_fd_sc_hd__dlygate4sd3_1
X_19907_ net7534 net3260 _03561_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__mux2_1
Xhold2606 _00688_ vssd1 vssd1 vccd1 vccd1 net3133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2617 rbzero.pov.spi_buffer\[9\] vssd1 vssd1 vccd1 vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2628 net7497 vssd1 vssd1 vccd1 vccd1 net3155 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03507_ _03507_ vssd1 vssd1 vccd1 vccd1 clknet_0__03507_ sky130_fd_sc_hd__clkbuf_16
Xhold2639 net7533 vssd1 vssd1 vccd1 vccd1 net3166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 net7090 vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1916 _00908_ vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_19838_ net1857 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
Xhold1927 _04271_ vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 net7191 vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1949 net2502 vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 i_debug_map_overlay vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21800_ net242 net2603 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21731_ clknet_leaf_108_i_clk net4005 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21662_ clknet_leaf_23_i_clk net2714 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21593_ net227 net2281 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5210 net4374 vssd1 vssd1 vccd1 vccd1 net5737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5221 net3387 vssd1 vssd1 vccd1 vccd1 net5748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5232 net5733 vssd1 vssd1 vccd1 vccd1 net5759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5243 rbzero.pov.ready_buffer\[51\] vssd1 vssd1 vccd1 vccd1 net5770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5254 net3968 vssd1 vssd1 vccd1 vccd1 net5781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4520 net611 vssd1 vssd1 vccd1 vccd1 net5047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5265 _03069_ vssd1 vssd1 vccd1 vccd1 net5792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4531 _00827_ vssd1 vssd1 vccd1 vccd1 net5058 sky130_fd_sc_hd__dlygate4sd3_1
X_22145_ clknet_leaf_56_i_clk net901 vssd1 vssd1 vccd1 vccd1 reg_hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5287 net1710 vssd1 vssd1 vccd1 vccd1 net5814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4542 net707 vssd1 vssd1 vccd1 vccd1 net5069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5298 rbzero.pov.ready_buffer\[67\] vssd1 vssd1 vccd1 vccd1 net5825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4553 rbzero.spi_registers.texadd0\[4\] vssd1 vssd1 vccd1 vccd1 net5080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4564 net843 vssd1 vssd1 vccd1 vccd1 net5091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4575 _00869_ vssd1 vssd1 vccd1 vccd1 net5102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3830 net8165 vssd1 vssd1 vccd1 vccd1 net4357 sky130_fd_sc_hd__clkbuf_2
Xhold4586 net769 vssd1 vssd1 vccd1 vccd1 net5113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3841 net959 vssd1 vssd1 vccd1 vccd1 net4368 sky130_fd_sc_hd__dlygate4sd3_1
X_22076_ net518 net977 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4597 rbzero.spi_registers.texadd1\[2\] vssd1 vssd1 vccd1 vccd1 net5124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3852 net7853 vssd1 vssd1 vccd1 vccd1 net4379 sky130_fd_sc_hd__buf_1
Xhold3863 net8058 vssd1 vssd1 vccd1 vccd1 net4390 sky130_fd_sc_hd__buf_1
Xhold3874 net3484 vssd1 vssd1 vccd1 vccd1 net4401 sky130_fd_sc_hd__buf_1
X_21027_ clknet_leaf_53_i_clk net4264 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3885 net7796 vssd1 vssd1 vccd1 vccd1 net4412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3896 net8252 vssd1 vssd1 vccd1 vccd1 net4423 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19767__47 clknet_1_1__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
X_12800_ _05969_ _05973_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a21o_4
XFILLER_0_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13780_ _06949_ _06950_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__xor2_2
X_10992_ net5716 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _05901_ net4068 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nand2_1
X_21929_ net371 net2850 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20397__149 clknet_1_1__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__inv_2
XFILLER_0_132_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _08142_ _08277_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ net6627 _05799_ _05837_ net54 vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _07240_ _07145_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__nor2_1
X_11613_ _04771_ _04775_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__o21bai_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _08427_ _08428_ net8042 _08475_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12593_ net20 _05769_ _05772_ net21 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__and4b_1
XFILLER_0_93_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17120_ _10013_ _10138_ _10136_ _10137_ vssd1 vssd1 vccd1 vccd1 _10140_ sky130_fd_sc_hd__o211ai_2
X_14332_ _07459_ _07460_ _07481_ _07479_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ _04731_ net4095 _04682_ net4384 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_108_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17051_ _10070_ _10071_ vssd1 vssd1 vccd1 vccd1 _10072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14263_ _07383_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nor2_2
X_11475_ net5946 _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _09089_ net7766 _09093_ _09096_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13214_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__clkbuf_4
Xhold7190 _01251_ vssd1 vssd1 vccd1 vccd1 net7717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14194_ _07361_ _07362_ _07364_ _07290_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ _06265_ _06025_ _06315_ _04491_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _06029_ _06031_ _06050_ _06243_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__and4_1
X_17953_ _02090_ _02072_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__or2b_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16904_ _09907_ _09925_ vssd1 vssd1 vccd1 vccd1 _09926_ sky130_fd_sc_hd__xnor2_1
X_12027_ rbzero.tex_r1\[9\] rbzero.tex_r1\[8\] _04968_ vssd1 vssd1 vccd1 vccd1 _05216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17884_ _02114_ _02019_ _02120_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__and3_1
X_19623_ net1375 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
X_16835_ net3888 net4776 vssd1 vssd1 vccd1 vccd1 _09860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19554_ net3980 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
X_16766_ _09796_ _09797_ vssd1 vssd1 vccd1 vccd1 _09798_ sky130_fd_sc_hd__nand2_1
X_13978_ _07102_ _07130_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__or2b_1
X_18505_ _02627_ net6015 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15717_ _08810_ _08811_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__and2_1
X_12929_ net4354 _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__or2_1
X_16697_ _09738_ vssd1 vssd1 vccd1 vccd1 _09746_ sky130_fd_sc_hd__clkbuf_4
X_19485_ net1493 net6010 _03354_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20456__202 clknet_1_0__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__inv_2
X_18436_ net4724 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ _08742_ _08740_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__xnor2_2
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15579_ _08665_ _08672_ _08673_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__nand3_1
X_18367_ net3494 rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1 vccd1 _02553_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17318_ _10213_ _10215_ _10212_ vssd1 vssd1 vccd1 vccd1 _10337_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ net1678 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17249_ _10267_ _10256_ vssd1 vssd1 vccd1 vccd1 _10268_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20260_ net4024 net4103 net4111 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20191_ net4501 _03744_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or2_1
Xhold3104 rbzero.spi_registers.spi_buffer\[23\] vssd1 vssd1 vccd1 vccd1 net3631 sky130_fd_sc_hd__clkbuf_2
Xhold3115 _04497_ vssd1 vssd1 vccd1 vccd1 net3642 sky130_fd_sc_hd__buf_1
XFILLER_0_122_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3126 _03322_ vssd1 vssd1 vccd1 vccd1 net3653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3137 _01223_ vssd1 vssd1 vccd1 vccd1 net3664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2403 net7341 vssd1 vssd1 vccd1 vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3148 net7616 vssd1 vssd1 vccd1 vccd1 net3675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2414 net5734 vssd1 vssd1 vccd1 vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2425 _01506_ vssd1 vssd1 vccd1 vccd1 net2952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2436 _04429_ vssd1 vssd1 vccd1 vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1702 net6974 vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2447 net2088 vssd1 vssd1 vccd1 vccd1 net2974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 _04359_ vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 _04050_ vssd1 vssd1 vccd1 vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2469 net7428 vssd1 vssd1 vccd1 vccd1 net2996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1724 net5646 vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1735 net3025 vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1746 _01545_ vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1757 _01382_ vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1768 net7150 vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1779 net5672 vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ clknet_leaf_127_i_clk net3438 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ clknet_leaf_117_i_clk net3140 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_50 _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21576_ net210 net2815 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_61 _08038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20527_ clknet_1_1__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__buf_1
XFILLER_0_127_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_83 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_94 net8264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ net5568 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5040 _04457_ vssd1 vssd1 vccd1 vccd1 net5567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5051 _04123_ vssd1 vssd1 vccd1 vccd1 net5578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5062 rbzero.tex_b1\[32\] vssd1 vssd1 vccd1 vccd1 net5589 sky130_fd_sc_hd__dlygate4sd3_1
X_11191_ net6540 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
Xhold5073 net2041 vssd1 vssd1 vccd1 vccd1 net5600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5084 net1919 vssd1 vssd1 vccd1 vccd1 net5611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4350 _08462_ vssd1 vssd1 vccd1 vccd1 net4877 sky130_fd_sc_hd__buf_2
Xhold5095 net2474 vssd1 vssd1 vccd1 vccd1 net5622 sky130_fd_sc_hd__buf_1
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22128_ clknet_leaf_53_i_clk net5583 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold4361 _01649_ vssd1 vssd1 vccd1 vccd1 net4888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4372 net3784 vssd1 vssd1 vccd1 vccd1 net4899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4383 rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1 vccd1 net4910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4394 gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3660 _04477_ vssd1 vssd1 vccd1 vccd1 net4187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3671 net8117 vssd1 vssd1 vccd1 vccd1 net4198 sky130_fd_sc_hd__dlygate4sd3_1
X_14950_ _08072_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
X_22059_ net501 net2882 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold3682 net988 vssd1 vssd1 vccd1 vccd1 net4209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3693 rbzero.wall_tracer.visualWallDist\[2\] vssd1 vssd1 vccd1 vccd1 net4220 sky130_fd_sc_hd__buf_1
Xhold2970 _01226_ vssd1 vssd1 vccd1 vccd1 net3497 sky130_fd_sc_hd__dlygate4sd3_1
X_13901_ _06703_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__clkbuf_4
X_14881_ _08031_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
Xhold2981 net8037 vssd1 vssd1 vccd1 vccd1 net3508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2992 net5931 vssd1 vssd1 vccd1 vccd1 net3519 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16620_ _09590_ _09709_ vssd1 vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__xnor2_2
X_13832_ _06999_ _07001_ _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ _08509_ _09025_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13763_ _06930_ _06932_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__a21bo_1
X_10975_ net7256 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap85 _04851_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _08287_ _08335_ _08596_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ net4128 _05043_ net28 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16482_ _09570_ _09572_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__xor2_4
X_19270_ net5412 _03216_ _03228_ _03219_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13694_ _06752_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15433_ _08315_ _08316_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__and2_1
X_18221_ _02436_ _02437_ _09845_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a21o_1
X_12645_ net46 _05817_ _05799_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15364_ _08410_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18152_ _02378_ net3785 _02320_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ net21 net20 _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__and3_1
X_17103_ _09997_ _09998_ vssd1 vssd1 vccd1 vccd1 _10124_ sky130_fd_sc_hd__or2b_1
Xclkbuf_0__03841_ _03841_ vssd1 vssd1 vccd1 vccd1 clknet_0__03841_ sky130_fd_sc_hd__clkbuf_16
X_14315_ _07417_ _07421_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__xnor2_4
X_18083_ _09788_ net3700 _02317_ _09793_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a31o_1
X_11527_ net4152 _04464_ _04501_ net8170 _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a221o_1
X_15295_ _08389_ _08221_ _08241_ _08384_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__or4_1
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17034_ _10025_ _10026_ _10054_ vssd1 vssd1 vccd1 vccd1 _10055_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _07310_ _07416_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__xnor2_4
Xhold309 net7084 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _04500_ _04647_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14177_ _07240_ _07281_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_108_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11389_ _04545_ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13128_ _06297_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nor2_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ net3412 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17936_ _01794_ _10220_ _02083_ _02081_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__o31a_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _06190_ _06197_ _06200_ _06220_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a41o_1
Xhold1009 _03060_ vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17867_ _01971_ _01972_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19606_ net1020 _03139_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16818_ net4865 vssd1 vssd1 vccd1 vccd1 _09845_ sky130_fd_sc_hd__buf_4
X_17798_ _02035_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19746__28 clknet_1_1__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
XFILLER_0_191_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19537_ net3770 net4833 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nor2_1
X_16749_ net2968 _09103_ _09782_ vssd1 vssd1 vccd1 vccd1 _09783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19468_ net1533 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18419_ _02589_ _02593_ _02599_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__o21ai_2
X_19399_ net5440 _03302_ _03304_ _03299_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7915 net7807 vssd1 vssd1 vccd1 vccd1 net8442 sky130_fd_sc_hd__dlygate4sd3_1
X_21430_ clknet_leaf_26_i_clk net3522 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21361_ clknet_leaf_6_i_clk net5278 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20312_ net1503 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold810 net6340 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
X_21292_ clknet_leaf_34_i_clk net5159 vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold821 _00994_ vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold832 _03555_ vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20510__251 clknet_1_1__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__inv_2
Xhold843 _01256_ vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
X_20243_ net4024 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__inv_2
Xhold854 _02498_ vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 net3744 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _03391_ vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 net5508 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_20174_ _03706_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__clkbuf_4
Xhold898 net4073 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2200 _01056_ vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2211 net7004 vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2222 _01467_ vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2233 _00691_ vssd1 vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 net1194 vssd1 vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1510 _01387_ vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2255 _01586_ vssd1 vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1521 _00750_ vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2266 rbzero.tex_r0\[1\] vssd1 vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 net7446 vssd1 vssd1 vccd1 vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1532 net5619 vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2288 _01063_ vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1543 _03567_ vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2299 net7430 vssd1 vssd1 vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1554 _00661_ vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1565 _04148_ vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1576 _01508_ vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1587 _04326_ vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 net7044 vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_87_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10760_ net6243 net7015 _04194_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10691_ net7095 net6152 _04149_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_10_i_clk clknet_4_2__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12430_ _05263_ _05602_ _05606_ _05614_ _04991_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o311a_1
XFILLER_0_191_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21628_ clknet_leaf_129_i_clk net3344 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ reg_rgb\[22\] _05546_ _05054_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21559_ net193 net1732 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ _07268_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__xnor2_1
X_11312_ net7747 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__buf_4
X_15080_ net5859 net3489 net3417 vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_25_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12292_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _04916_ vssd1 vssd1 vccd1 vccd1 _05478_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14031_ _07163_ _07175_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or2_1
X_11243_ net6932 net2832 _04445_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__mux2_1
X_11174_ net7393 net7391 _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4180 _00431_ vssd1 vssd1 vccd1 vccd1 net4707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4191 net4233 vssd1 vssd1 vccd1 vccd1 net4718 sky130_fd_sc_hd__clkbuf_2
X_18770_ _09739_ net4858 net8243 net3762 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__a31o_1
X_15982_ _08624_ _08654_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3490 _03083_ vssd1 vssd1 vccd1 vccd1 net4017 sky130_fd_sc_hd__dlygate4sd3_1
X_17721_ _01958_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__nor2_1
X_14933_ net4655 _06239_ _08052_ net3835 net4675 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__o221a_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _01790_ _01800_ _01798_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a21o_1
X_14864_ _08018_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ _09555_ _09557_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__and2b_1
X_13815_ _06982_ _06984_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_187_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17583_ _01821_ _01822_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14795_ _07958_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19322_ net5181 _03250_ _03258_ _03259_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__o211a_1
X_16534_ _09615_ _09623_ vssd1 vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__xnor2_1
X_13746_ _06703_ _06808_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nor2_1
X_10958_ net6776 net2017 _04298_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19253_ net6325 _03217_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16465_ _09422_ _09424_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__or2b_1
X_13677_ _06846_ _06847_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__nor2_1
X_10889_ net7051 net2900 _04253_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18204_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15416_ _08211_ _08207_ _08221_ _08241_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__or4_1
X_12628_ _05803_ _05805_ _05806_ net26 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a2bb2o_1
X_16396_ _09486_ _09378_ _09376_ vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19184_ net6542 _03170_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15347_ _08441_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__inv_2
X_18135_ _02363_ net3757 _02320_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
X_12559_ net14 _05721_ _05739_ net15 vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5809 _02482_ vssd1 vssd1 vccd1 vccd1 net6336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20568__303 clknet_1_1__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__inv_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold106 net6029 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
X_15278_ net3777 _08118_ _08137_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__o21ai_2
X_18066_ _02298_ _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__xnor2_1
Xhold117 _01373_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold128 net7211 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17017_ _10036_ _10037_ vssd1 vssd1 vccd1 vccd1 _10038_ sky130_fd_sc_hd__xnor2_1
Xhold139 net5032 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _07311_ _07396_ _07398_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ net2427 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _02156_ net4655 _10260_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ net1947 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
X_20930_ clknet_leaf_60_i_clk net4573 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20861_ net4204 _04001_ _04002_ _10257_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20792_ net969 net5692 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20337__95 clknet_1_0__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__inv_2
XFILLER_0_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7701 rbzero.traced_texa\[6\] vssd1 vssd1 vccd1 vccd1 net8228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7723 rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 net8250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7734 net8071 vssd1 vssd1 vccd1 vccd1 net8261 sky130_fd_sc_hd__clkbuf_2
X_21413_ clknet_leaf_38_i_clk net4232 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7745 rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 net8272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7789 net7751 vssd1 vssd1 vccd1 vccd1 net8316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21344_ clknet_leaf_46_i_clk net5131 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 _01147_ vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_21275_ clknet_leaf_25_i_clk net5543 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold651 net4370 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 net6228 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20226_ net4686 _03710_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__or2_1
Xhold673 net6256 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 net6252 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 net6511 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
X_20157_ net1057 _03707_ _03731_ _03732_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__o211a_1
Xhold2030 net7382 vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2041 _01436_ vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2052 net6891 vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2063 _04269_ vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2074 net7096 vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
X_20088_ net3326 _08299_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__or2_2
Xhold2085 _01516_ vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1340 _03598_ vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2096 net5670 vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1351 net3769 vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ net3431 _05100_ _05104_ net4169 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a2111o_1
Xhold1362 _04356_ vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1373 net6761 vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1384 _01034_ vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 _01358_ vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ net5965 _05050_ net6044 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a21o_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06722_ _06723_ _06724_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__o21a_2
XFILLER_0_95_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ net2521 net7171 _04216_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _07741_ _07744_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _04938_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__buf_2
X_10743_ net6617 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16250_ _09248_ _09269_ _09341_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13462_ _06624_ _06628_ _06631_ _06632_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__o22a_1
XFILLER_0_165_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20517__257 clknet_1_1__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__inv_2
X_10674_ net6086 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ net3461 _08261_ net2898 vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__o21ai_1
X_12413_ _05465_ _05593_ _05597_ _05263_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a211o_1
XFILLER_0_211_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16181_ _09163_ _09166_ _09164_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13393_ _06516_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15132_ net4583 _08137_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__nor2_1
X_12344_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _05249_ vssd1 vssd1 vccd1 vccd1 _05530_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19940_ net3283 net3060 _03572_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__mux2_1
X_15063_ net3536 net4168 vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__xnor2_2
X_12275_ net3871 _04653_ net4148 _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ _07183_ _07184_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__or2_1
X_11226_ net6768 net2345 _04434_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux2_1
X_19871_ net3173 net6649 _03539_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
X_18822_ net3485 _02951_ _02953_ net7695 vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__a211o_1
X_11157_ net6103 net2572 _04401_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18753_ rbzero.wall_tracer.rayAddendY\[6\] _02902_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02903_ sky130_fd_sc_hd__mux2_1
X_11088_ net2557 net7306 _04364_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
X_15965_ net8015 _08129_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__nand2_4
X_17704_ _01741_ _01943_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__xnor2_1
X_14916_ net8029 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__o21a_1
X_18684_ net3678 net4528 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__xor2_2
XFILLER_0_37_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15896_ _08656_ _08990_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__xnor2_4
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _10186_ _09060_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ net7794 _07946_ _08003_ net4704 vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__a211o_2
XFILLER_0_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ _09537_ _10350_ _10348_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_129_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14778_ net7843 _07821_ _07863_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ net5137 _03236_ _03249_ _03246_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__o211a_1
X_16517_ _09605_ _09606_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13729_ _06897_ net539 _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__a21oi_2
X_17497_ _10273_ _01717_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ net6440 _03203_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or2_1
X_16448_ _09536_ _09538_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7008 rbzero.pov.ready_buffer\[62\] vssd1 vssd1 vccd1 vccd1 net7535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7019 net3180 vssd1 vssd1 vccd1 vccd1 net7546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6307 net1926 vssd1 vssd1 vccd1 vccd1 net6834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19167_ net3842 _03123_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__nand2_2
X_16379_ _09468_ _09469_ vssd1 vssd1 vccd1 vccd1 _09470_ sky130_fd_sc_hd__nand2_1
Xhold6318 rbzero.tex_b1\[21\] vssd1 vssd1 vccd1 vccd1 net6845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6329 net2564 vssd1 vssd1 vccd1 vccd1 net6856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18118_ _02348_ net4565 _02320_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5606 _03481_ vssd1 vssd1 vccd1 vccd1 net6133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5617 net1064 vssd1 vssd1 vccd1 vccd1 net6144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19098_ net3367 _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__or2_1
Xhold5628 rbzero.tex_b0\[40\] vssd1 vssd1 vccd1 vccd1 net6155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5639 net1081 vssd1 vssd1 vccd1 vccd1 net6166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4905 net1024 vssd1 vssd1 vccd1 vccd1 net5432 sky130_fd_sc_hd__dlygate4sd3_1
X_18049_ _10316_ _09345_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4916 rbzero.spi_registers.texadd0\[23\] vssd1 vssd1 vccd1 vccd1 net5443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4927 net1123 vssd1 vssd1 vccd1 vccd1 net5454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4938 _00901_ vssd1 vssd1 vccd1 vccd1 net5465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4949 net1108 vssd1 vssd1 vccd1 vccd1 net5476 sky130_fd_sc_hd__dlygate4sd3_1
X_21060_ clknet_leaf_68_i_clk _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20011_ net4441 _08238_ _03614_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20622__352 clknet_1_1__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__inv_2
X_21962_ net404 net2378 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20913_ clknet_4_12__leaf_i_clk _00400_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21893_ net335 net1902 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _09721_ clknet_1_0__leaf__05898_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__and2_2
XFILLER_0_77_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20775_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7520 _02562_ vssd1 vssd1 vccd1 vccd1 net8047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7531 net3468 vssd1 vssd1 vccd1 vccd1 net8058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7542 _00517_ vssd1 vssd1 vccd1 vccd1 net8069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7553 _00520_ vssd1 vssd1 vccd1 vccd1 net8080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6830 net2887 vssd1 vssd1 vccd1 vccd1 net7357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7575 rbzero.pov.ready_buffer\[13\] vssd1 vssd1 vccd1 vccd1 net8102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6841 rbzero.tex_r0\[47\] vssd1 vssd1 vccd1 vccd1 net7368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7586 net1675 vssd1 vssd1 vccd1 vccd1 net8113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6852 net2489 vssd1 vssd1 vccd1 vccd1 net7379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7597 _00507_ vssd1 vssd1 vccd1 vccd1 net8124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6863 rbzero.tex_b0\[41\] vssd1 vssd1 vccd1 vccd1 net7390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6874 net2333 vssd1 vssd1 vccd1 vccd1 net7401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21327_ clknet_leaf_45_i_clk net5031 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6885 rbzero.tex_b0\[7\] vssd1 vssd1 vccd1 vccd1 net7412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6896 net2604 vssd1 vssd1 vccd1 vccd1 net7423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12060_ _04923_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__clkbuf_8
Xhold470 net6117 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
X_21258_ clknet_leaf_22_i_clk net3795 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold481 net7891 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11011_ net6550 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
Xhold492 _01303_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20209_ _09725_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__buf_4
X_21189_ clknet_leaf_129_i_clk net3294 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _08832_ _08844_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__xor2_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _06062_ _06043_ net4044 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 net6622 vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 _01104_ vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _05101_ _05089_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__nor2_4
X_14701_ net3775 vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__buf_4
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 net6604 vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
X_15681_ _08180_ _08252_ _08254_ _08245_ net7836 vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__a32o_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ net3469 _06030_ _06068_ net3990 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _10435_ _10436_ vssd1 vssd1 vccd1 vccd1 _10438_ sky130_fd_sc_hd__or2_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ net4080 _05025_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a21bo_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _07790_ _07802_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__xnor2_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _10367_ _10369_ vssd1 vssd1 vccd1 vccd1 _10370_ sky130_fd_sc_hd__xor2_2
XFILLER_0_173_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14563_ _07306_ _07391_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__nor2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ _04942_ _04948_ _04956_ _04964_ _04817_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__o311a_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _09392_ _09393_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__xnor2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ net2811 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13514_ _06430_ _06432_ _06553_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__mux2_1
X_17282_ _10299_ _10300_ vssd1 vssd1 vccd1 vccd1 _10301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14494_ _07658_ _07662_ _07664_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19021_ net1493 net4076 _03078_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
X_16233_ _09323_ _09325_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__xor2_4
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13445_ _06492_ _06612_ _06613_ _06615_ _06538_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__a311o_1
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10657_ net6920 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16164_ _09253_ _09255_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _06527_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__clkbuf_4
X_10588_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ _04915_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__or2_1
X_15115_ net3637 _08162_ _08185_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16095_ _09162_ _09188_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__xnor2_1
X_15046_ _06120_ net8072 vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__or2_1
X_19923_ net2312 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12258_ _04847_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11209_ net6673 net1758 _04423_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__mux2_1
X_19854_ net7540 net1752 _03528_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__mux2_1
X_12189_ _04706_ _05375_ _05376_ net4139 vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18805_ net3940 net4814 net3084 vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__and3b_1
X_16997_ _09888_ _10002_ vssd1 vssd1 vccd1 vccd1 _10018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18736_ _02856_ net4686 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__xor2_1
X_15948_ _09030_ _09042_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18667_ _02813_ _02814_ _02815_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a21bo_1
X_15879_ _08938_ _08955_ _08973_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17618_ _01758_ _01775_ _01773_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18598_ _02752_ _02757_ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17549_ _01788_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19219_ net6321 _03169_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6104 net1746 vssd1 vssd1 vccd1 vccd1 net6631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6115 rbzero.tex_g1\[25\] vssd1 vssd1 vccd1 vccd1 net6642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6126 net1834 vssd1 vssd1 vccd1 vccd1 net6653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6137 rbzero.pov.spi_buffer\[73\] vssd1 vssd1 vccd1 vccd1 net6664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6148 net1731 vssd1 vssd1 vccd1 vccd1 net6675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5403 _01182_ vssd1 vssd1 vccd1 vccd1 net5930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5414 _03353_ vssd1 vssd1 vccd1 vccd1 net5941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6159 rbzero.pov.ready_buffer\[54\] vssd1 vssd1 vccd1 vccd1 net6686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5425 net3778 vssd1 vssd1 vccd1 vccd1 net5952 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5436 net3142 vssd1 vssd1 vccd1 vccd1 net5963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22161_ clknet_leaf_96_i_clk net4717 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5447 net3893 vssd1 vssd1 vccd1 vccd1 net5974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4702 _00813_ vssd1 vssd1 vccd1 vccd1 net5229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5458 _01242_ vssd1 vssd1 vccd1 vccd1 net5985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4713 net799 vssd1 vssd1 vccd1 vccd1 net5240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4724 rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 net5251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5469 net2321 vssd1 vssd1 vccd1 vccd1 net5996 sky130_fd_sc_hd__dlygate4sd3_1
X_21112_ clknet_leaf_95_i_clk net3717 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold4735 net759 vssd1 vssd1 vccd1 vccd1 net5262 sky130_fd_sc_hd__dlygate4sd3_1
X_22092_ net154 net2130 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4746 _00877_ vssd1 vssd1 vccd1 vccd1 net5273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4757 net878 vssd1 vssd1 vccd1 vccd1 net5284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4768 rbzero.spi_registers.texadd2\[7\] vssd1 vssd1 vccd1 vccd1 net5295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4779 net815 vssd1 vssd1 vccd1 vccd1 net5306 sky130_fd_sc_hd__dlygate4sd3_1
X_21043_ clknet_leaf_61_i_clk _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21945_ net387 net1987 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03512_ clknet_0__03512_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03512_
+ sky130_fd_sc_hd__clkbuf_16
X_21876_ net318 net926 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20827_ net4084 _04485_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _04749_ _04660_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__or2_1
X_20758_ _03925_ _03928_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10511_ net2774 net6259 _04053_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11491_ net3431 _04501_ _04600_ net3991 _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20689_ _09727_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7350 net4350 vssd1 vssd1 vccd1 vccd1 net7877 sky130_fd_sc_hd__dlygate4sd3_1
X_13230_ _06308_ _06400_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__xor2_2
Xhold7361 net4210 vssd1 vssd1 vccd1 vccd1 net7888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10442_ _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__buf_4
Xhold7372 rbzero.traced_texVinit\[6\] vssd1 vssd1 vccd1 vccd1 net7899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7383 net1105 vssd1 vssd1 vccd1 vccd1 net7910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7394 _00501_ vssd1 vssd1 vccd1 vccd1 net7921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6660 rbzero.pov.ready_buffer\[20\] vssd1 vssd1 vccd1 vccd1 net7187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _04491_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nand2_1
Xhold6671 net2555 vssd1 vssd1 vccd1 vccd1 net7198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6682 rbzero.tex_g1\[34\] vssd1 vssd1 vccd1 vccd1 net7209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6693 net2635 vssd1 vssd1 vccd1 vccd1 net7220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _04949_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5970 _03832_ vssd1 vssd1 vccd1 vccd1 net6497 sky130_fd_sc_hd__dlygate4sd3_1
X_13092_ _05980_ _05983_ net8051 _05984_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__a211oi_4
Xhold5981 net1270 vssd1 vssd1 vccd1 vccd1 net6508 sky130_fd_sc_hd__dlygate4sd3_1
X_20629__358 clknet_1_1__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__inv_2
Xhold5992 rbzero.spi_registers.new_texadd\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 net6519
+ sky130_fd_sc_hd__dlygate4sd3_1
X_16920_ _09640_ _09643_ vssd1 vssd1 vccd1 vccd1 _09942_ sky130_fd_sc_hd__nand2_1
X_12043_ _05204_ _05229_ _05231_ _05213_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f__05946_ clknet_0__05946_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05946_
+ sky130_fd_sc_hd__clkbuf_16
X_16851_ _09874_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__clkbuf_1
X_15802_ _08161_ _08318_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ net7395 net1426 _03403_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
X_16782_ _09812_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__clkbuf_1
X_13994_ _07108_ _07110_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__and2_1
X_18521_ _02627_ net4828 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__nand2_1
X_15733_ _08825_ _08824_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__and2b_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__buf_4
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18452_ _02630_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__or2_1
X_15664_ _08756_ _08758_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__nor2_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _06031_ _06050_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__a21o_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _10419_ _10420_ vssd1 vssd1 vccd1 vccd1 _10421_ sky130_fd_sc_hd__nor2_1
X_14615_ _07508_ _07785_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__xnor2_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _05014_ _05016_ _04909_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__a21oi_1
X_18383_ net3661 _02566_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__nand2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _08658_ _08689_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__xor2_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _10105_ _10226_ vssd1 vssd1 vccd1 vccd1 _10353_ sky130_fd_sc_hd__and2_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20374__128 clknet_1_0__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__inv_2
X_11758_ _04943_ _04944_ _04946_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o211a_1
X_14546_ _07712_ _07715_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10709_ net2319 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17265_ _10153_ _10154_ _10152_ vssd1 vssd1 vccd1 vccd1 _10284_ sky130_fd_sc_hd__a21boi_1
X_14477_ _07627_ _07646_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__a21oi_2
X_11689_ net4057 _04868_ _04867_ net4105 _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__o221a_1
XFILLER_0_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19004_ net6327 net5898 _02992_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16216_ _09162_ _09188_ _09308_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__05742_ _05742_ vssd1 vssd1 vccd1 vccd1 clknet_0__05742_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13428_ _06491_ _06597_ _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__and3_1
X_17196_ _10214_ _10215_ vssd1 vssd1 vccd1 vccd1 _10216_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ _09122_ _09120_ _09119_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13359_ _06455_ _06459_ _06461_ _06463_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__o31a_1
Xhold4009 net8332 vssd1 vssd1 vccd1 vccd1 net4536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _08010_ _08017_ _08021_ _08439_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__nor4_4
Xhold3308 net3380 vssd1 vssd1 vccd1 vccd1 net3835 sky130_fd_sc_hd__clkbuf_2
Xhold3319 net7971 vssd1 vssd1 vccd1 vccd1 net3846 sky130_fd_sc_hd__dlygate4sd3_1
X_19906_ net3215 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
X_15029_ _08123_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__buf_4
Xhold2607 net7452 vssd1 vssd1 vccd1 vccd1 net3134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 net2956 vssd1 vssd1 vccd1 vccd1 net3145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _03538_ vssd1 vssd1 vccd1 vccd1 net3156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03506_ _03506_ vssd1 vssd1 vccd1 vccd1 clknet_0__03506_ sky130_fd_sc_hd__clkbuf_16
Xhold1906 _04201_ vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_19837_ net3019 net3145 _03517_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
Xhold1917 net7199 vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1928 _01384_ vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 _04076_ vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 i_debug_trace_overlay vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
XFILLER_0_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18719_ _02869_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19699_ net6625 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21730_ clknet_leaf_109_i_clk net3930 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21661_ clknet_leaf_24_i_clk net3288 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21592_ net226 net1763 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5200 _01618_ vssd1 vssd1 vccd1 vccd1 net5727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5211 rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 net5738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5222 rbzero.pov.ready_buffer\[47\] vssd1 vssd1 vccd1 vccd1 net5749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5233 _03704_ vssd1 vssd1 vccd1 vccd1 net5760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5244 net3323 vssd1 vssd1 vccd1 vccd1 net5771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5255 rbzero.pov.ready_buffer\[64\] vssd1 vssd1 vccd1 vccd1 net5782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4510 net703 vssd1 vssd1 vccd1 vccd1 net5037 sky130_fd_sc_hd__dlygate4sd3_1
X_22144_ clknet_leaf_40_i_clk _01631_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold4521 rbzero.color_sky\[4\] vssd1 vssd1 vccd1 vccd1 net5048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5266 net3192 vssd1 vssd1 vccd1 vccd1 net5793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5277 _02798_ vssd1 vssd1 vccd1 vccd1 net5804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4532 net690 vssd1 vssd1 vccd1 vccd1 net5059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5288 rbzero.pov.ready_buffer\[60\] vssd1 vssd1 vccd1 vccd1 net5815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4543 _00852_ vssd1 vssd1 vccd1 vccd1 net5070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4554 net711 vssd1 vssd1 vccd1 vccd1 net5081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5299 net1703 vssd1 vssd1 vccd1 vccd1 net5826 sky130_fd_sc_hd__buf_1
Xhold3820 net8170 vssd1 vssd1 vccd1 vccd1 net4347 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold4565 rbzero.spi_registers.texadd0\[0\] vssd1 vssd1 vccd1 vccd1 net5092 sky130_fd_sc_hd__dlygate4sd3_1
X_22075_ net517 net3116 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold4576 net743 vssd1 vssd1 vccd1 vccd1 net5103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3831 _00777_ vssd1 vssd1 vccd1 vccd1 net4358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4587 _00859_ vssd1 vssd1 vccd1 vccd1 net5114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3842 net8164 vssd1 vssd1 vccd1 vccd1 net4369 sky130_fd_sc_hd__clkbuf_2
Xhold3853 net7869 vssd1 vssd1 vccd1 vccd1 net4380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4598 net752 vssd1 vssd1 vccd1 vccd1 net5125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3864 net7940 vssd1 vssd1 vccd1 vccd1 net4391 sky130_fd_sc_hd__dlygate4sd3_1
X_21026_ clknet_leaf_53_i_clk net4255 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3875 net8323 vssd1 vssd1 vccd1 vccd1 net4402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3886 net7798 vssd1 vssd1 vccd1 vccd1 net4413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3897 _02754_ vssd1 vssd1 vccd1 vccd1 net4424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_92_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10991_ net5640 net5714 _04309_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _05901_ net4156 vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__or2_1
X_21928_ net370 net2740 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ net48 _05817_ _05818_ clknet_1_1__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _05840_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21859_ net301 net1893 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _04776_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__nor2_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _07033_ _07326_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__or2_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15380_ _08472_ _08474_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__nor2_1
X_12592_ _05747_ _05749_ net4147 _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14331_ _07456_ _07501_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__xnor2_1
X_11543_ net1163 _04732_ _04679_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17050_ _09262_ _08411_ vssd1 vssd1 vccd1 vccd1 _10071_ sky130_fd_sc_hd__nor2_1
X_14262_ _07385_ _07428_ _07432_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ net3955 net3858 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__nor2_2
X_16001_ _09091_ net8542 _09094_ net3418 vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13213_ _06382_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__and2_1
Xhold7180 gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 net7707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7191 rbzero.color_floor\[4\] vssd1 vssd1 vccd1 vccd1 net7718 sky130_fd_sc_hd__dlygate4sd3_1
X_14193_ _07347_ _07363_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6490 net2094 vssd1 vssd1 vccd1 vccd1 net7017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ net8263 _06265_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17952_ _02111_ _02128_ _02126_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a21o_1
X_13075_ _06247_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__nor2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16903_ _09923_ _09924_ vssd1 vssd1 vccd1 vccd1 _09925_ sky130_fd_sc_hd__nor2_1
X_12026_ rbzero.tex_r1\[11\] rbzero.tex_r1\[10\] _04968_ vssd1 vssd1 vccd1 vccd1 _05215_
+ sky130_fd_sc_hd__mux2_1
X_17883_ _02114_ _02019_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19622_ net6367 net2205 _03430_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
X_16834_ net3888 net4776 vssd1 vssd1 vccd1 vccd1 _09859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _03320_ net3979 vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__and2_1
X_16765_ net4506 net4535 vssd1 vssd1 vccd1 vccd1 _09797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13977_ _07142_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__nand2_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18504_ _02559_ net4869 net8258 net3615 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a31o_1
X_15716_ _08708_ _08753_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__xor2_4
XFILLER_0_158_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12928_ net7687 vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__clkbuf_4
X_19484_ net1594 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
X_16696_ _09736_ vssd1 vssd1 vccd1 vccd1 _09745_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ _02601_ _02612_ _02613_ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15647_ _08674_ _08728_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__nand2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ net4043 vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__buf_1
XFILLER_0_68_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18366_ net3493 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__clkbuf_1
X_15578_ _08634_ _08660_ _08664_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__a21o_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _10313_ _10335_ vssd1 vssd1 vccd1 vccd1 _10336_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14529_ _07308_ _07391_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18297_ net6585 net3562 _02493_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17248_ _10253_ vssd1 vssd1 vccd1 vccd1 _10267_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17179_ _10197_ _10198_ vssd1 vssd1 vccd1 vccd1 _10199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20190_ net8103 _03743_ net4734 _03732_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3105 net7602 vssd1 vssd1 vccd1 vccd1 net3632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3116 net5209 vssd1 vssd1 vccd1 vccd1 net3643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3127 _00890_ vssd1 vssd1 vccd1 vccd1 net3654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3138 net8367 vssd1 vssd1 vccd1 vccd1 net3665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2404 _04384_ vssd1 vssd1 vccd1 vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3149 _00739_ vssd1 vssd1 vccd1 vccd1 net3676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 _00705_ vssd1 vssd1 vccd1 vccd1 net2942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2426 net7697 vssd1 vssd1 vccd1 vccd1 net2953 sky130_fd_sc_hd__buf_2
Xhold2437 _01048_ vssd1 vssd1 vccd1 vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 net6976 vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _03566_ vssd1 vssd1 vccd1 vccd1 net2975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _01304_ vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 _01580_ vssd1 vssd1 vccd1 vccd1 net2986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 _01566_ vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1736 _03525_ vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1747 net6947 vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1758 net7388 vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 _01492_ vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21713_ clknet_leaf_103_i_clk net4465 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_1__f_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21644_ clknet_leaf_117_i_clk net2071 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21575_ net209 net2675 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_40 net4490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 rbzero.tex_b0\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_73 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_95 net8270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5030 rbzero.tex_r1\[0\] vssd1 vssd1 vccd1 vccd1 net5557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5041 net1837 vssd1 vssd1 vccd1 vccd1 net5568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5052 net2582 vssd1 vssd1 vccd1 vccd1 net5579 sky130_fd_sc_hd__dlygate4sd3_1
X_11190_ net6538 net1773 _04412_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__mux2_1
Xhold5063 _04354_ vssd1 vssd1 vccd1 vccd1 net5590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5074 rbzero.tex_r0\[2\] vssd1 vssd1 vccd1 vccd1 net5601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4340 _02669_ vssd1 vssd1 vccd1 vccd1 net4867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5085 rbzero.spi_registers.new_mapd\[4\] vssd1 vssd1 vccd1 vccd1 net5612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5096 _01614_ vssd1 vssd1 vccd1 vccd1 net5623 sky130_fd_sc_hd__dlygate4sd3_1
X_22127_ clknet_leaf_53_i_clk net5624 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold4351 rbzero.wall_tracer.rayAddendY\[-7\] vssd1 vssd1 vccd1 vccd1 net4878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4362 net790 vssd1 vssd1 vccd1 vccd1 net4889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4373 rbzero.pov.ready_buffer\[53\] vssd1 vssd1 vccd1 vccd1 net4900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4384 net3765 vssd1 vssd1 vccd1 vccd1 net4911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3650 _04670_ vssd1 vssd1 vccd1 vccd1 net4177 sky130_fd_sc_hd__buf_2
Xhold4395 net602 vssd1 vssd1 vccd1 vccd1 net4922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22058_ net500 net2273 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold3661 net4283 vssd1 vssd1 vccd1 vccd1 net4188 sky130_fd_sc_hd__clkbuf_2
Xhold3672 _00832_ vssd1 vssd1 vccd1 vccd1 net4199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3683 net7887 vssd1 vssd1 vccd1 vccd1 net4210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3694 net8000 vssd1 vssd1 vccd1 vccd1 net4221 sky130_fd_sc_hd__dlygate4sd3_1
X_21009_ clknet_leaf_37_i_clk net4337 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13900_ _07030_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xnor2_2
Xhold2960 net5865 vssd1 vssd1 vccd1 vccd1 net3487 sky130_fd_sc_hd__dlygate4sd3_1
X_14880_ net4608 _08030_ net3775 vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__mux2_1
Xhold2982 net7735 vssd1 vssd1 vccd1 vccd1 net3509 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_2_2_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
Xhold2993 _03361_ vssd1 vssd1 vccd1 vccd1 net3520 sky130_fd_sc_hd__dlygate4sd3_1
X_13831_ _06715_ _06708_ _06813_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f__05645_ clknet_0__05645_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05645_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16550_ _08799_ _08403_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ net7254 net2715 _04298_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__mux2_1
X_13762_ _06729_ _06931_ _06727_ _06758_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__nand4_2
XFILLER_0_35_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap75 _09172_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_6
X_15501_ _08325_ _08334_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__nor2_1
Xmax_cap86 net87 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ net4102 net4024 net5965 net6044 net28 net31 vssd1 vssd1 vccd1 vccd1 _05891_
+ sky130_fd_sc_hd__mux4_1
X_16481_ _09370_ _09439_ _09571_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__a21oi_4
X_13693_ _06827_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18220_ _02436_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nor2_1
X_15432_ _08311_ _08318_ _08323_ _08307_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__o31a_1
X_12644_ _05814_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _02376_ _02377_ _09864_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__o21ai_1
X_15363_ _08457_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12575_ _05747_ net18 net19 vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17102_ _10023_ _10122_ vssd1 vssd1 vccd1 vccd1 _10123_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_0__03840_ _03840_ vssd1 vssd1 vccd1 vccd1 clknet_0__03840_ sky130_fd_sc_hd__clkbuf_16
X_14314_ _07471_ _07477_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__xor2_4
XFILLER_0_145_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18082_ net3749 net4381 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__or2_1
X_11526_ net2185 _04022_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__xor2_1
X_15294_ _08168_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__buf_2
XFILLER_0_124_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _10038_ _10053_ vssd1 vssd1 vccd1 vccd1 _10054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14245_ _07284_ _07281_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nor2_2
X_11457_ _04500_ _04461_ _04648_ _04468_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14176_ _07314_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__xor2_2
X_20486__229 clknet_1_1__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__inv_2
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11388_ rbzero.spi_registers.texadd2\[23\] _04506_ _04548_ rbzero.spi_registers.texadd1\[23\]
+ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a221o_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13127_ net3719 net3614 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nor2_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ net7520 net5835 _03058_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _02170_ _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__and2_1
X_13058_ _06182_ _06233_ _06168_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__o21a_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _05190_ _05192_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__o21ai_1
X_17866_ _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19605_ _02475_ net4844 _03312_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16817_ net4633 _09843_ vssd1 vssd1 vccd1 vccd1 _09844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17797_ _01917_ _01929_ _01927_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19536_ _03352_ net3624 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__nor2_1
X_16748_ net2968 _09103_ _09780_ vssd1 vssd1 vccd1 vccd1 _09782_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19467_ net1396 net6014 _03345_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ net4271 _09741_ _09742_ net3502 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18418_ _02589_ _02593_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19398_ net2447 _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18349_ _02536_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__buf_4
XFILLER_0_174_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7916 _06553_ vssd1 vssd1 vccd1 vccd1 net8443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21360_ clknet_leaf_6_i_clk net5183 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20311_ net6470 net3562 _03825_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold800 _01006_ vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_21291_ clknet_leaf_26_i_clk net5470 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03869_ clknet_0__03869_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03869_
+ sky130_fd_sc_hd__clkbuf_16
Xhold811 net6342 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 net6324 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _01120_ vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
X_20242_ net4111 net4103 net5983 _05673_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__or4b_1
Xhold844 net6383 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 _00586_ vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold866 _03415_ vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 _00938_ vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold888 net5510 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
X_20173_ net3713 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
Xhold899 net4075 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__buf_4
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2201 net7347 vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2212 _04236_ vssd1 vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2223 net7078 vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2234 net7034 vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1500 _04035_ vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 _03532_ vssd1 vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2256 net7339 vssd1 vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 net8161 vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__clkbuf_2
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2267 net5602 vssd1 vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 rbzero.tex_g1\[60\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 _04410_ vssd1 vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 net6006 vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1544 _01131_ vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2289 rbzero.tex_r0\[45\] vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1555 net6945 vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 _01494_ vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1577 net5612 vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1588 _01334_ vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1599 net7046 vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20591__324 clknet_1_1__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__inv_2
XFILLER_0_48_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ net2729 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21627_ clknet_leaf_127_i_clk net3150 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ net4163 _05544_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__and3_1
X_21558_ net192 net1760 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _04913_ vssd1 vssd1 vccd1 vccd1 _05477_
+ sky130_fd_sc_hd__mux2_1
X_21489_ clknet_leaf_11_i_clk net1470 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14030_ _07179_ _07181_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or2_1
X_11242_ net6217 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11173_ _04264_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4170 net2197 vssd1 vssd1 vccd1 vccd1 net4697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4181 net3422 vssd1 vssd1 vccd1 vccd1 net4708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4192 _08060_ vssd1 vssd1 vccd1 vccd1 net4719 sky130_fd_sc_hd__dlygate4sd3_1
X_15981_ _08621_ _09075_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17720_ _01847_ _01850_ _01848_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__o21a_1
Xhold3480 _06064_ vssd1 vssd1 vccd1 vccd1 net4007 sky130_fd_sc_hd__clkbuf_2
Xhold3491 _00725_ vssd1 vssd1 vccd1 vccd1 net4018 sky130_fd_sc_hd__dlygate4sd3_1
X_14932_ net8088 _06237_ _04482_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__o21a_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _01858_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__xnor2_1
Xhold2790 net7780 vssd1 vssd1 vccd1 vccd1 net3317 sky130_fd_sc_hd__clkbuf_2
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ net4440 _08017_ _07976_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__mux2_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16602_ _09690_ _09691_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__or2_2
X_13814_ _06981_ _06980_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__or2b_1
X_17582_ _01821_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14794_ net4392 net7825 _07872_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19321_ _03205_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__buf_4
X_16533_ _09621_ _09622_ vssd1 vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__nor2_1
X_13745_ _06708_ net3607 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__nor2_1
X_10957_ net6508 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19252_ net5388 _03216_ _03218_ _03219_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__o211a_1
X_16464_ _09539_ _09554_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__xnor2_2
X_13676_ _06842_ _06843_ _06845_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__nor3_1
X_10888_ net6886 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18203_ _02414_ _02416_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15415_ _08229_ _08509_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ net4149 net4141 net4164 net7727 _05802_ net25 vssd1 vssd1 vccd1 vccd1 _05806_
+ sky130_fd_sc_hd__mux4_1
X_19183_ net5364 _03168_ _03178_ _03176_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__o211a_1
X_16395_ _09374_ _09375_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18134_ _02361_ _02362_ _09847_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__o21ai_1
X_15346_ _08113_ _08440_ _08123_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12558_ net12 _05690_ _05723_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18065_ _02299_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__xnor2_1
X_11509_ net2898 net3955 _04584_ net3461 _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a221o_1
X_15277_ _08113_ _08369_ _08371_ _08118_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__o211a_2
Xhold107 net6031 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net8 _05670_ net9 vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__and3b_1
Xhold118 net7489 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _08543_ net7818 vssd1 vssd1 vccd1 vccd1 _10037_ sky130_fd_sc_hd__and2_1
Xhold129 net5641 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14228_ _07311_ _07396_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159_ _07195_ _07329_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ net6201 net4901 net2874 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _09788_ _02059_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a21o_1
X_18898_ net3186 net7188 _03014_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
X_17849_ _01794_ _10096_ _02024_ _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20540__278 clknet_1_1__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__inv_2
X_20860_ net4217 _04001_ _04002_ _10132_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19519_ net1493 net6494 net3086 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__mux2_1
X_20791_ net969 net5692 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7702 _03968_ vssd1 vssd1 vccd1 vccd1 net8229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7713 _08046_ vssd1 vssd1 vccd1 vccd1 net8240 sky130_fd_sc_hd__dlygate4sd3_1
X_21412_ clknet_leaf_38_i_clk net5565 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7724 net4167 vssd1 vssd1 vccd1 vccd1 net8251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7735 rbzero.debug_overlay.vplaneY\[-7\] vssd1 vssd1 vccd1 vccd1 net8262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7746 rbzero.wall_tracer.trackDistX\[9\] vssd1 vssd1 vccd1 vccd1 net8273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21343_ clknet_leaf_19_i_clk net5091 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7779 rbzero.row_render.size\[0\] vssd1 vssd1 vccd1 vccd1 net8306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20434__183 clknet_1_0__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__inv_2
XFILLER_0_170_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold630 net5465 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21274_ clknet_leaf_25_i_clk net5529 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 net6230 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 net6222 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold663 _01463_ vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20225_ net3577 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold674 _03828_ vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 net6254 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 net6513 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
X_20156_ _09725_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__clkbuf_4
Xhold2020 _01330_ vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 net7384 vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2042 net7179 vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2053 _01285_ vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
X_20087_ net4284 _03662_ net2397 _03316_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a211o_1
Xhold2064 _01386_ vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 _04378_ vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1330 _03527_ vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1341 _01160_ vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2086 net6626 vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 _01325_ vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 _02471_ vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1363 _01307_ vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _04275_ vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1385 net6751 vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1396 net6646 vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11860_ net7716 net4138 net4177 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and3_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ net2652 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11791_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _04978_ vssd1 vssd1 vccd1 vccd1 _04981_
+ sky130_fd_sc_hd__mux2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20989_ clknet_leaf_112_i_clk net4060 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13530_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__buf_2
X_10742_ net2417 net6615 _04182_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ net6084 net2294 _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__mux2_1
X_13461_ _06505_ _06543_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__nand2_2
XFILLER_0_153_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15200_ net2898 net3461 _08261_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__or3_4
X_12412_ _05517_ _05594_ _05596_ _05306_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16180_ _09272_ _08392_ _09158_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13392_ _06557_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__or3_1
XFILLER_0_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15131_ _08225_ vssd1 vssd1 vccd1 vccd1 _08226_ sky130_fd_sc_hd__buf_4
X_12343_ _04943_ _05528_ _04947_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12274_ net4172 _05460_ _04656_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__a21o_1
X_15062_ net3536 _08156_ vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11225_ net2918 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__clkbuf_1
X_14013_ _07149_ _07150_ _07182_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__and3_1
X_19870_ net2180 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11156_ net2540 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__clkbuf_1
X_18821_ _02963_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18752_ _02893_ _02894_ _02901_ _02526_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a2bb2o_1
X_15964_ _08544_ _08549_ _08546_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__a21o_1
X_11087_ net3244 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
X_17703_ _01940_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__xor2_1
X_14915_ net3796 _08050_ _08052_ net3790 net4577 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__o221a_1
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18683_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__xnor2_1
X_15895_ _08754_ _08760_ _08759_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__a21o_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _10432_ _08612_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__or2_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ _07934_ _08000_ _08002_ net7824 vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17565_ _01684_ _01686_ _01683_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ net7813 _07895_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__a21oi_1
X_11989_ net4127 _04600_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19304_ net1514 _03238_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ _09601_ _09604_ _09599_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ _06885_ _06896_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__and2b_1
X_17496_ _01714_ _01716_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19235_ net5352 _03201_ _03209_ _03206_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__o211a_1
X_16447_ _09537_ _09170_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13659_ net83 _06771_ _06829_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__o21ai_1
Xhold7009 net3269 vssd1 vssd1 vccd1 vccd1 net7536 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_71_i_clk clknet_4_13__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19166_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__buf_4
X_16378_ _08543_ _09225_ _09347_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6308 rbzero.tex_r1\[57\] vssd1 vssd1 vccd1 vccd1 net6835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6319 net2107 vssd1 vssd1 vccd1 vccd1 net6846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ _02346_ net3733 _09829_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__o21ai_1
X_15329_ _08422_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5607 net2138 vssd1 vssd1 vccd1 vccd1 net6134 sky130_fd_sc_hd__dlygate4sd3_1
X_19097_ net3623 _03123_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nand2_4
Xhold5618 _04091_ vssd1 vssd1 vccd1 vccd1 net6145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5629 net1052 vssd1 vssd1 vccd1 vccd1 net6156 sky130_fd_sc_hd__dlygate4sd3_1
X_18048_ _02164_ _02182_ _02181_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_197_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4906 _00772_ vssd1 vssd1 vccd1 vccd1 net5433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4917 net1067 vssd1 vssd1 vccd1 vccd1 net5444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4928 rbzero.spi_registers.texadd2\[14\] vssd1 vssd1 vccd1 vccd1 net5455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4939 net1157 vssd1 vssd1 vccd1 vccd1 net5466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20010_ net5904 _03607_ net3545 _03339_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__o211a_1
X_19999_ net5816 _08158_ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21961_ net403 net2553 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ clknet_leaf_78_i_clk _00399_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_21892_ net334 net1141 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20843_ _03998_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__buf_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20774_ _03942_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_i_clk clknet_4_9__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7510 net4414 vssd1 vssd1 vccd1 vccd1 net8037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7521 _02563_ vssd1 vssd1 vccd1 vccd1 net8048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7543 net4226 vssd1 vssd1 vccd1 vccd1 net8070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7554 rbzero.wall_tracer.stepDistY\[-8\] vssd1 vssd1 vccd1 vccd1 net8081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6820 rbzero.tex_r0\[16\] vssd1 vssd1 vccd1 vccd1 net7347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7565 _02821_ vssd1 vssd1 vccd1 vccd1 net8092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6831 rbzero.tex_r1\[48\] vssd1 vssd1 vccd1 vccd1 net7358 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7576 net638 vssd1 vssd1 vccd1 vccd1 net8103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6842 net2581 vssd1 vssd1 vccd1 vccd1 net7369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7587 _00632_ vssd1 vssd1 vccd1 vccd1 net8114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6853 rbzero.tex_g1\[40\] vssd1 vssd1 vccd1 vccd1 net7380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7598 rbzero.traced_texa\[-7\] vssd1 vssd1 vccd1 vccd1 net8125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6864 net2673 vssd1 vssd1 vccd1 vccd1 net7391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21326_ clknet_leaf_45_i_clk net5230 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6875 rbzero.tex_r0\[52\] vssd1 vssd1 vccd1 vccd1 net7402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6886 net3005 vssd1 vssd1 vccd1 vccd1 net7413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6897 rbzero.pov.sclk_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net7424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21257_ clknet_leaf_22_i_clk net3633 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold460 _03223_ vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold471 net6119 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net2253 net6548 _04320_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__mux2_1
Xhold482 net8223 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20208_ _02627_ _03744_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__or2_1
Xhold493 net8174 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_1
XFILLER_0_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21188_ clknet_leaf_127_i_clk net3181 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_20139_ _03689_ net7653 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or2_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _06104_ net4034 net3965 _06060_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__or4_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 _01269_ vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 net6624 vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net3774 _04485_ _04479_ _06117_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__and4_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 net5811 vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _04684_ _05073_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nand2_1
X_15680_ net8414 _08774_ _08271_ _08252_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__or4b_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _00589_ vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ net7712 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__inv_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _07800_ _07801_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__nor2_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net4079 _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__or2_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _10182_ _10240_ _10368_ vssd1 vssd1 vccd1 vccd1 _10369_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _07704_ _07728_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__nand2_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _04958_ _04960_ _04963_ _04928_ _04824_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a221o_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _08244_ _08430_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__nand2_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _06676_ _06611_ _06616_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__nand3_1
XFILLER_0_181_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17281_ _10298_ _10297_ vssd1 vssd1 vccd1 vccd1 _10300_ sky130_fd_sc_hd__and2b_1
X_10725_ net7117 net2907 _04097_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _07620_ _07663_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19020_ net4031 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
X_16232_ _08992_ _09083_ _09208_ _09324_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__a31oi_4
X_13444_ _06441_ _06549_ _06614_ _06550_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10656_ net6918 net2155 _04138_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ _09253_ _09255_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10587_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__buf_4
X_13375_ net559 _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__nor2_2
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15114_ _08179_ _08174_ _08173_ _08172_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__a2bb2o_1
X_12326_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _04912_ vssd1 vssd1 vccd1 vccd1 _05512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16094_ _09185_ _09187_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__xor2_2
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ net8261 _08119_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__nand2_2
XFILLER_0_142_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19922_ net2802 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
X_12257_ rbzero.tex_g1\[57\] rbzero.tex_g1\[56\] _04837_ vssd1 vssd1 vccd1 vccd1 _05444_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ net2608 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__clkbuf_1
X_19853_ net3078 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
X_12188_ _05040_ _04691_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20606__337 clknet_1_0__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__inv_2
X_18804_ net1878 net3083 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__nand2_1
X_11139_ net2280 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__clkbuf_1
X_16996_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10017_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15947_ _09039_ _09041_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__xor2_2
X_18735_ _02853_ _02871_ _02846_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18666_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _08947_ _08953_ _08955_ _08938_ _08972_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17617_ _01855_ _01856_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__nor2_1
X_14829_ _07983_ _07984_ _07985_ _07987_ _07913_ net7785 vssd1 vssd1 vccd1 vccd1 _07988_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_176_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18597_ net4635 net4879 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17548_ _01786_ _01787_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ _01718_ _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20652__379 clknet_1_0__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__inv_2
X_19218_ net5436 _03167_ _03197_ _03189_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6105 rbzero.tex_g0\[5\] vssd1 vssd1 vccd1 vccd1 net6632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6116 net1652 vssd1 vssd1 vccd1 vccd1 net6643 sky130_fd_sc_hd__dlygate4sd3_1
X_20351__107 clknet_1_0__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__inv_2
X_19149_ net2066 _03147_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__or2_1
Xhold6127 rbzero.tex_g0\[6\] vssd1 vssd1 vccd1 vccd1 net6654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6138 net1613 vssd1 vssd1 vccd1 vccd1 net6665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6149 rbzero.spi_registers.new_texadd\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net6676
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5404 rbzero.spi_registers.got_new_floor vssd1 vssd1 vccd1 vccd1 net5931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5415 rbzero.spi_registers.got_new_other vssd1 vssd1 vccd1 vccd1 net5942 sky130_fd_sc_hd__dlygate4sd3_1
X_22160_ clknet_leaf_96_i_clk net5035 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5426 _02708_ vssd1 vssd1 vccd1 vccd1 net5953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5437 gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 net5964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4703 net853 vssd1 vssd1 vccd1 vccd1 net5230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5448 _06145_ vssd1 vssd1 vccd1 vccd1 net5975 sky130_fd_sc_hd__dlygate4sd3_1
X_21111_ clknet_leaf_94_i_clk net3636 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold5459 net3338 vssd1 vssd1 vccd1 vccd1 net5986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4714 _00791_ vssd1 vssd1 vccd1 vccd1 net5241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4725 net866 vssd1 vssd1 vccd1 vccd1 net5252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22091_ net153 net2231 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4736 rbzero.spi_registers.texadd1\[0\] vssd1 vssd1 vccd1 vccd1 net5263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4747 net983 vssd1 vssd1 vccd1 vccd1 net5274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4758 _00823_ vssd1 vssd1 vccd1 vccd1 net5285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21042_ clknet_leaf_64_i_clk _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4769 net902 vssd1 vssd1 vccd1 vccd1 net5296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20546__284 clknet_1_0__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__inv_2
XFILLER_0_158_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21944_ net386 net2517 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03511_ clknet_0__03511_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03511_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ net317 net2112 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ net3871 net3976 net4083 _03988_ _06237_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a41o_1
XFILLER_0_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20757_ net984 net5448 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ net2561 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ _04679_ net3552 net3990 _04465_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20688_ _03352_ net920 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7340 net4382 vssd1 vssd1 vccd1 vccd1 net7867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7351 net3426 vssd1 vssd1 vccd1 vccd1 net7878 sky130_fd_sc_hd__dlygate4sd3_1
X_10441_ net7710 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7362 net1023 vssd1 vssd1 vccd1 vccd1 net7889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7373 net4218 vssd1 vssd1 vccd1 vccd1 net7900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7395 net4297 vssd1 vssd1 vccd1 vccd1 net7922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6650 rbzero.pov.spi_buffer\[44\] vssd1 vssd1 vccd1 vccd1 net7177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6661 net791 vssd1 vssd1 vccd1 vccd1 net7188 sky130_fd_sc_hd__dlygate4sd3_1
X_13160_ _06276_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__xnor2_2
Xhold6672 rbzero.tex_r0\[51\] vssd1 vssd1 vccd1 vccd1 net7199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6683 net2459 vssd1 vssd1 vccd1 vccd1 net7210 sky130_fd_sc_hd__dlygate4sd3_1
X_12111_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _04951_ vssd1 vssd1 vccd1 vccd1 _05299_
+ sky130_fd_sc_hd__mux2_1
Xhold6694 rbzero.tex_r0\[26\] vssd1 vssd1 vccd1 vccd1 net7221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5960 rbzero.tex_r0\[19\] vssd1 vssd1 vccd1 vccd1 net6487 sky130_fd_sc_hd__dlygate4sd3_1
X_13091_ _06241_ _06261_ _06262_ _06242_ net5408 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21309_ clknet_leaf_5_i_clk net5374 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5971 net1577 vssd1 vssd1 vccd1 vccd1 net6498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5982 rbzero.spi_registers.new_texadd\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net6509
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12042_ _05206_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__or2_1
Xhold5993 net1811 vssd1 vssd1 vccd1 vccd1 net6520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold290 net4596 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
X_16850_ _09873_ net4665 net4649 vssd1 vssd1 vccd1 vccd1 _09874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _08868_ _08873_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__xnor2_1
X_16781_ _09811_ net3945 _09769_ vssd1 vssd1 vccd1 vccd1 _09812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13993_ _06857_ _07124_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__and2b_1
XFILLER_0_172_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18520_ _02627_ net4828 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__or2_1
X_15732_ _08797_ _08802_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__xor2_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12944_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ net4603 net3509 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15663_ _08704_ _08707_ _08757_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__o21a_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12875_ net3807 net3447 _06028_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__o21a_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19793__71 clknet_1_1__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17402_ _10292_ _10301_ _10299_ vssd1 vssd1 vccd1 vccd1 _10420_ sky130_fd_sc_hd__a21oi_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _07506_ _07559_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__nor2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ net3781 _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__and2_1
X_18382_ net3661 _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _08676_ _08688_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__and2_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17333_ _10106_ _10351_ vssd1 vssd1 vccd1 vccd1 _10352_ sky130_fd_sc_hd__xnor2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14545_ _07489_ _07198_ _07713_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__or3_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _04829_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__buf_4
XFILLER_0_166_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ _10281_ _10282_ vssd1 vssd1 vccd1 vccd1 _10283_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ net2661 net7035 _04160_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ _07628_ _07645_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11688_ _04871_ _04877_ _04868_ net4057 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a22o_1
X_19003_ net5766 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
X_16215_ _09185_ _09187_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ _06531_ _06533_ _06447_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__a21o_1
X_10639_ net7019 net6822 _04127_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__mux2_1
X_17195_ _09272_ _09403_ vssd1 vssd1 vccd1 vccd1 _10215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _09228_ _09238_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _06491_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__xnor2_4
X_12309_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _05239_ vssd1 vssd1 vccd1 vccd1 _05495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16077_ _08458_ _09170_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ _06346_ _06404_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__and2_1
Xhold3309 net7970 vssd1 vssd1 vccd1 vccd1 net3836 sky130_fd_sc_hd__dlygate4sd3_1
X_19905_ net3214 net7534 _03561_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__mux2_1
X_15028_ _08122_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__buf_4
Xhold2608 _03569_ vssd1 vssd1 vccd1 vccd1 net3135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2619 _03529_ vssd1 vssd1 vccd1 vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19836_ net3027 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
Xhold1907 _01447_ vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1918 _04120_ vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1929 net6986 vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16979_ _09596_ _09703_ _09702_ _09701_ vssd1 vssd1 vccd1 vccd1 _10001_ sky130_fd_sc_hd__o2bb2a_1
Xinput3 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_4
XFILLER_0_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18718_ net4709 net3575 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__and2_1
X_19698_ net6623 net3674 _03468_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18649_ net3619 _02805_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21660_ clknet_leaf_24_i_clk net1167 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21591_ net225 net1821 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5201 net2754 vssd1 vssd1 vccd1 vccd1 net5728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5212 net3189 vssd1 vssd1 vccd1 vccd1 net5739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5223 net1906 vssd1 vssd1 vccd1 vccd1 net5750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5234 _03705_ vssd1 vssd1 vccd1 vccd1 net5761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5245 _03678_ vssd1 vssd1 vccd1 vccd1 net5772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4500 net718 vssd1 vssd1 vccd1 vccd1 net5027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5256 net4441 vssd1 vssd1 vccd1 vccd1 net5783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4511 _00828_ vssd1 vssd1 vccd1 vccd1 net5038 sky130_fd_sc_hd__dlygate4sd3_1
X_22143_ clknet_leaf_44_i_clk _01630_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold4522 net691 vssd1 vssd1 vccd1 vccd1 net5049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5278 net3524 vssd1 vssd1 vccd1 vccd1 net5805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4533 rbzero.spi_registers.texadd1\[9\] vssd1 vssd1 vccd1 vccd1 net5060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5289 net1535 vssd1 vssd1 vccd1 vccd1 net5816 sky130_fd_sc_hd__buf_1
Xhold4544 net708 vssd1 vssd1 vccd1 vccd1 net5071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3810 net745 vssd1 vssd1 vccd1 vccd1 net4337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4555 _00787_ vssd1 vssd1 vccd1 vccd1 net5082 sky130_fd_sc_hd__dlygate4sd3_1
X_22074_ net516 net2154 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold3821 _00759_ vssd1 vssd1 vccd1 vccd1 net4348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4566 net723 vssd1 vssd1 vccd1 vccd1 net5093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3832 net838 vssd1 vssd1 vccd1 vccd1 net4359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4577 rbzero.spi_registers.texadd3\[8\] vssd1 vssd1 vccd1 vccd1 net5104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4588 net770 vssd1 vssd1 vccd1 vccd1 net5115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3843 _00768_ vssd1 vssd1 vccd1 vccd1 net4370 sky130_fd_sc_hd__dlygate4sd3_1
X_21025_ clknet_leaf_53_i_clk net4222 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3854 net7871 vssd1 vssd1 vccd1 vccd1 net4381 sky130_fd_sc_hd__buf_1
Xhold4599 _00809_ vssd1 vssd1 vccd1 vccd1 net5126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3865 net7942 vssd1 vssd1 vccd1 vccd1 net4392 sky130_fd_sc_hd__buf_1
Xhold3876 net8325 vssd1 vssd1 vccd1 vccd1 net4403 sky130_fd_sc_hd__buf_1
Xhold3887 net8036 vssd1 vssd1 vccd1 vccd1 net4414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3898 net8098 vssd1 vssd1 vccd1 vccd1 net4425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10990_ net5642 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21927_ net369 net2967 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ net55 _05818_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a21o_1
X_21858_ net300 net2118 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _04781_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20809_ net991 net5739 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nor2_1
X_12591_ net43 _05744_ _05764_ net44 _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21789_ clknet_leaf_21_i_clk net1221 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _07482_ _07499_ _07500_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a21oi_1
X_11542_ net4384 net4393 net4366 net2587 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _07429_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__or2b_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ net3857 net3641 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__nand2_1
Xhold7170 rbzero.spi_registers.spi_buffer\[9\] vssd1 vssd1 vccd1 vccd1 net7697 sky130_fd_sc_hd__dlygate4sd3_1
X_16000_ net5929 net4168 _04511_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13212_ net8035 net8051 _04491_ _06263_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a211o_4
Xhold7181 net3857 vssd1 vssd1 vccd1 vccd1 net7708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7192 net3644 vssd1 vssd1 vccd1 vccd1 net7719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14192_ _07240_ _07305_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6480 net2849 vssd1 vssd1 vccd1 vccd1 net7007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6491 rbzero.tex_r0\[40\] vssd1 vssd1 vccd1 vccd1 net7018 sky130_fd_sc_hd__dlygate4sd3_1
X_13143_ _06311_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__xnor2_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5790 net1362 vssd1 vssd1 vccd1 vccd1 net6317 sky130_fd_sc_hd__dlygate4sd3_1
X_17951_ _02186_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__nand2_1
X_13074_ net5428 _06244_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__nor2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16902_ _09921_ _09922_ vssd1 vssd1 vccd1 vccd1 _09924_ sky130_fd_sc_hd__and2_1
X_12025_ _05204_ _05210_ _05212_ _05213_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__o211a_1
X_17882_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19621_ net1545 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
X_16833_ _09850_ _09851_ _09852_ vssd1 vssd1 vccd1 vccd1 _09858_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16764_ net4506 net4535 vssd1 vssd1 vccd1 vccd1 _09796_ sky130_fd_sc_hd__or2_1
X_19552_ net3978 _03139_ net1777 _03386_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a22o_1
X_13976_ _07143_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15715_ _08763_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__nor2_1
X_18503_ net3614 _09736_ _02679_ _04490_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ net3983 _04743_ _06060_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__a21oi_1
X_16695_ net8120 _09743_ _09744_ net4917 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
X_19483_ net1396 net6050 _03354_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15646_ _08720_ _08722_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__xor2_2
X_18434_ _04490_ _02614_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ _06032_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nor2_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _04976_ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _02541_ _02542_ _02543_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15577_ _08667_ _08671_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12789_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__nor2_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _10333_ _10334_ vssd1 vssd1 vccd1 vccd1 _10335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _07306_ _07327_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__nor2_1
X_18296_ net1457 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _10250_ _10252_ vssd1 vssd1 vccd1 vccd1 _10266_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14459_ _07629_ _07620_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17178_ _10195_ _10196_ vssd1 vssd1 vccd1 vccd1 _10198_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ _09150_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3106 _00744_ vssd1 vssd1 vccd1 vccd1 net3633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3117 net7718 vssd1 vssd1 vccd1 vccd1 net3644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3128 net7948 vssd1 vssd1 vccd1 vccd1 net3655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3139 _02388_ vssd1 vssd1 vccd1 vccd1 net3666 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2405 _01281_ vssd1 vssd1 vccd1 vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
X_20463__208 clknet_1_0__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__inv_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2416 net7408 vssd1 vssd1 vccd1 vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2427 net7525 vssd1 vssd1 vccd1 vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2438 net7042 vssd1 vssd1 vccd1 vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1704 _01578_ vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 _01130_ vssd1 vssd1 vccd1 vccd1 net2976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1715 net7594 vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1726 net7239 vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
X_19819_ net7312 net3329 _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_1
Xhold1737 _01093_ vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1748 net6949 vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1759 net5575 vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21712_ clknet_leaf_103_i_clk net4475 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20658__385 clknet_1_1__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__inv_2
XFILLER_0_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19772__52 clknet_1_0__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20357__113 clknet_1_1__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__inv_2
X_21643_ clknet_leaf_116_i_clk net2976 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21574_ net208 net1054 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_30 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_41 net4694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 rbzero.wall_tracer.visualWallDist\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_74 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_85 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_96 _04942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5020 rbzero.tex_r1\[28\] vssd1 vssd1 vccd1 vccd1 net5547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5031 net1275 vssd1 vssd1 vccd1 vccd1 net5558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5042 rbzero.spi_registers.new_other\[10\] vssd1 vssd1 vccd1 vccd1 net5569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5053 rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 net5580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5064 net2215 vssd1 vssd1 vccd1 vccd1 net5591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5075 _04174_ vssd1 vssd1 vccd1 vccd1 net5602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4330 _02908_ vssd1 vssd1 vccd1 vccd1 net4857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4341 _02670_ vssd1 vssd1 vccd1 vccd1 net4868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22126_ clknet_leaf_53_i_clk net5490 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold5086 net2104 vssd1 vssd1 vccd1 vccd1 net5613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5097 net2475 vssd1 vssd1 vccd1 vccd1 net5624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4352 net942 vssd1 vssd1 vccd1 vccd1 net4879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4363 net4331 vssd1 vssd1 vccd1 vccd1 net4890 sky130_fd_sc_hd__clkbuf_1
Xhold4374 net2426 vssd1 vssd1 vccd1 vccd1 net4901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4385 net4674 vssd1 vssd1 vccd1 vccd1 net4912 sky130_fd_sc_hd__buf_1
Xhold3640 net8250 vssd1 vssd1 vccd1 vccd1 net4167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4396 _01598_ vssd1 vssd1 vccd1 vccd1 net4923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3651 _05043_ vssd1 vssd1 vccd1 vccd1 net4178 sky130_fd_sc_hd__dlygate4sd3_1
X_22057_ net499 net1117 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold3662 _09712_ vssd1 vssd1 vccd1 vccd1 net4189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3673 net599 vssd1 vssd1 vccd1 vccd1 net4200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3684 net7889 vssd1 vssd1 vccd1 vccd1 net4211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3695 net865 vssd1 vssd1 vccd1 vccd1 net4222 sky130_fd_sc_hd__dlygate4sd3_1
X_21008_ clknet_leaf_38_i_clk net4261 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2950 net4662 vssd1 vssd1 vccd1 vccd1 net3477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2961 net8319 vssd1 vssd1 vccd1 vccd1 net3488 sky130_fd_sc_hd__clkbuf_2
Xhold2972 net5795 vssd1 vssd1 vccd1 vccd1 net3499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2983 _03757_ vssd1 vssd1 vccd1 vccd1 net3510 sky130_fd_sc_hd__dlygate4sd3_1
X_13830_ _06813_ _07000_ _06708_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__mux2_1
Xhold2994 _03362_ vssd1 vssd1 vccd1 vccd1 net3521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13761_ net556 _06931_ _06727_ _06758_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10973_ net6502 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ _08567_ _08594_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__xor2_2
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap76 _07692_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
Xmax_cap87 _04850_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_2
X_12712_ net4111 _05673_ net4071 net4092 net28 net30 vssd1 vssd1 vccd1 vccd1 _05890_
+ sky130_fd_sc_hd__mux4_1
X_16480_ _09436_ _09438_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__nor2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _06851_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ _08524_ _08525_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12643_ net51 net41 net40 _05203_ _05797_ _05802_ vssd1 vssd1 vccd1 vccd1 _05822_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_182_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ _02372_ _02375_ _09845_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a21o_1
X_15362_ net4168 _08162_ net8400 vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__o21ai_2
X_12574_ _05750_ _05752_ _05753_ net20 vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a2bb2o_1
X_17101_ _10120_ _10121_ vssd1 vssd1 vccd1 vccd1 _10122_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14313_ _07412_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__xnor2_4
X_18081_ net3749 net4381 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__nand2_1
X_11525_ _04709_ _04710_ _04711_ _04713_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15293_ _08385_ _08387_ _08377_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20676__21 clknet_1_0__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_0_68_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17032_ _10051_ _10052_ vssd1 vssd1 vccd1 vccd1 _10053_ sky130_fd_sc_hd__nor2_1
X_14244_ _07413_ _07360_ _07414_ net5902 vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ _04600_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ _07242_ net569 vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__nor2_1
X_11387_ _04566_ rbzero.spi_registers.texadd3\[23\] vssd1 vssd1 vccd1 vccd1 _04579_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ net3719 net3614 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ net1536 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _02168_ _02169_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__or2_1
X_13057_ _06193_ _06195_ _06231_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__o211a_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12008_ _05194_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nand2_1
X_17865_ _10190_ _09612_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19604_ net4842 _03139_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__nand2_1
Xnet99_2 clknet_leaf_67_i_clk vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
X_16816_ _09841_ _09842_ vssd1 vssd1 vccd1 vccd1 _09843_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17796_ _02012_ _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19535_ net5943 _03139_ _03344_ net3084 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__o2bb2a_1
X_16747_ net5722 _09769_ _09768_ _09781_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a22o_1
X_13959_ _07128_ _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16678_ net4335 _09741_ _09742_ net744 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a22o_1
X_19466_ net1734 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18417_ net3494 net4501 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__xor2_2
X_15629_ _08692_ _08693_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__xor2_2
X_19397_ net3217 _03141_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18348_ _04480_ _09734_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__nand2_1
Xhold7917 net7795 vssd1 vssd1 vccd1 vccd1 net8444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18279_ net2204 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20310_ net1201 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_8
XFILLER_0_47_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21290_ clknet_leaf_26_i_clk net4359 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03868_ clknet_0__03868_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03868_
+ sky130_fd_sc_hd__clkbuf_16
Xhold801 net6300 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold812 _00992_ vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 _03470_ vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
X_20241_ net4024 _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__nand2_1
Xhold834 net8307 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_1
Xhold845 net6385 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 net6553 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _00956_ vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_19809__86 clknet_1_0__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__inv_2
X_20172_ _03728_ net7646 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_1
Xhold878 net6387 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 net6418 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2202 _04158_ vssd1 vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2213 _01415_ vssd1 vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 net7080 vssd1 vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2235 net7036 vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1501 _01594_ vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 _01099_ vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1512 net5542 vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2257 _04229_ vssd1 vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2268 _01471_ vssd1 vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 net6797 vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2279 _01065_ vssd1 vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 net6008 vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 net6931 vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1556 _04389_ vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 net7016 vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1578 _03408_ vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 net6873 vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21626_ clknet_leaf_127_i_clk net1232 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21557_ net191 net2856 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ net3641 vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12290_ _05474_ _05475_ _05206_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21488_ clknet_leaf_12_i_clk net1630 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ net6215 net2072 _04445_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__mux2_1
X_20439_ clknet_1_0__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__buf_1
XFILLER_0_28_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20411__162 clknet_1_1__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__inv_2
X_11172_ net2655 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
Xhold4160 _03775_ vssd1 vssd1 vccd1 vccd1 net4687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22109_ net147 net3069 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold4171 rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 net4698 sky130_fd_sc_hd__buf_2
X_15980_ _09073_ _09074_ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__xor2_2
Xhold4182 rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 net4709 sky130_fd_sc_hd__buf_2
Xhold4193 _00430_ vssd1 vssd1 vccd1 vccd1 net4720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3470 net6045 vssd1 vssd1 vccd1 vccd1 net3997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3481 _06131_ vssd1 vssd1 vccd1 vccd1 net4008 sky130_fd_sc_hd__dlygate4sd3_1
X_14931_ net3913 _08050_ _08052_ net3820 net4706 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3492 rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1 net4019 sky130_fd_sc_hd__buf_2
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2780 _01166_ vssd1 vssd1 vccd1 vccd1 net3307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nand2_1
Xhold2791 net4364 vssd1 vssd1 vccd1 vccd1 net3318 sky130_fd_sc_hd__dlygate4sd3_1
X_14862_ _06505_ _08016_ _07869_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__a21o_2
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _09688_ _09689_ _09663_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__a21oi_1
X_13813_ _06960_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__nor2_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _01691_ _01699_ _01697_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_203_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14793_ _07949_ _07951_ _07956_ net7824 net4704 vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__a221o_1
X_16532_ _09504_ _09616_ _09620_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__and3_1
X_19320_ net1371 _03251_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13744_ _06706_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__nor2_1
X_10956_ net6506 net1920 _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16463_ _09551_ _09553_ vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__xor2_2
X_19251_ _03205_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_183_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ _06842_ _06843_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10887_ net6884 net1964 _04253_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
X_19751__33 clknet_1_0__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_15414_ _08266_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__clkbuf_4
X_18202_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12626_ _05802_ net7571 net26 _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a211o_1
X_19182_ net6297 _03170_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__or2_1
X_16394_ _09483_ _09484_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18133_ net8039 _02360_ _09845_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15345_ _05985_ _06416_ net4180 vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12557_ _05726_ _05737_ net14 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18064_ _10062_ _09974_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__nor2_1
X_11508_ net3457 net3641 vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__xor2_1
X_15276_ _08113_ net8498 vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12488_ net4147 _05643_ _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a211o_1
Xhold108 _01041_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17015_ _10034_ _10035_ vssd1 vssd1 vccd1 vccd1 _10036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold119 net4562 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ _07283_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__or2_1
X_11439_ rbzero.spi_registers.texadd0\[1\] rbzero.spi_registers.texadd0\[0\] _04020_
+ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _06696_ _07198_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _06693_ _06698_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__or2_1
X_18966_ net2875 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _02150_ _02153_ _02154_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__o21a_1
X_18897_ net2365 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17848_ _02022_ _02023_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17779_ _02016_ _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__xnor2_1
X_20575__309 clknet_1_0__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__inv_2
XFILLER_0_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19518_ net1737 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20790_ _03954_ _03956_ _03955_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_53_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19449_ net4312 _03334_ net1034 _03299_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7703 _01617_ vssd1 vssd1 vccd1 vccd1 net8230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7714 rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 net8241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21411_ clknet_leaf_38_i_clk net5516 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7725 rbzero.debug_overlay.vplaneY\[-9\] vssd1 vssd1 vccd1 vccd1 net8252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7736 net8018 vssd1 vssd1 vccd1 vccd1 net8263 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7747 net4761 vssd1 vssd1 vccd1 vccd1 net8274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7769 rbzero.row_render.size\[10\] vssd1 vssd1 vccd1 vccd1 net8296 sky130_fd_sc_hd__dlygate4sd3_1
X_21342_ clknet_leaf_20_i_clk net5370 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20469__214 clknet_1_1__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__inv_2
XFILLER_0_170_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 _00695_ vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
X_21273_ clknet_leaf_25_i_clk net5573 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold631 net6248 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 net6232 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 net6224 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20224_ _04459_ net3576 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__or2_1
Xhold664 net6242 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold675 _01266_ vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
X_20670__16 clknet_1_0__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold686 _00968_ vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold697 _00670_ vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
X_20155_ rbzero.debug_overlay.facingY\[-8\] _03711_ vssd1 vssd1 vccd1 vccd1 _03731_
+ sky130_fd_sc_hd__or2_1
Xhold2010 _04381_ vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 net7120 vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2032 _01295_ vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2043 net7181 vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
X_20086_ net2396 _03631_ _03659_ _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o211a_1
Xhold2054 net7368 vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _01496_ vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2065 net7251 vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _01095_ vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2076 _01287_ vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1342 net7509 vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2087 _04018_ vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2098 net7221 vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1353 _02473_ vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1364 net6632 vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 _01380_ vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _04079_ vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1397 _03443_ vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20441__188 clknet_1_1__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__inv_2
X_10810_ net7171 net7250 _04216_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _04979_ vssd1 vssd1 vccd1 vccd1 _04980_
+ sky130_fd_sc_hd__mux2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20988_ clknet_leaf_112_i_clk net3920 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ net2701 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ _06547_ _06630_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ _04104_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _04922_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21609_ clknet_leaf_132_i_clk net3147 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ _06392_ _06558_ _06561_ _06491_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15130_ _08118_ _08223_ _08224_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _05258_ vssd1 vssd1 vccd1 vccd1 _05528_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15061_ _06370_ _08150_ net8412 _08155_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__a31o_4
X_12273_ net4140 _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__nand2_1
X_14012_ _07149_ _07150_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__a21oi_2
X_11224_ net7387 net6768 _04434_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ net3935 _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__xnor2_1
X_11155_ net7363 net6103 _04401_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18751_ _02899_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__xnor2_1
X_15963_ _08562_ _08540_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__or2b_1
X_11086_ net7306 net7530 _04364_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17702_ _01743_ _01834_ _01941_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a21oi_1
X_14914_ net8021 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__o21a_1
X_15894_ _08761_ _08812_ _08986_ _08988_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__a22o_4
X_18682_ net4764 _02825_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__and2_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _01784_ _01760_ _01783_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__or3_1
X_14845_ _07934_ _08001_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__nand2_1
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17564_ _01781_ _01804_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__xnor2_1
X_14776_ net7833 net8354 vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11988_ net4126 net4057 _04462_ net4160 vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a2bb2o_1
X_19303_ net5073 _03236_ _03248_ _03246_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__o211a_1
X_16515_ _09599_ _09601_ _09604_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__and3_1
X_13727_ net551 _06879_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__xor2_1
X_10939_ net6723 net2217 _04287_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17495_ _01734_ _01735_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19234_ net6504 _03203_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or2_1
X_16446_ _08417_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__clkbuf_4
X_13658_ _06577_ _06726_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _05747_ _05749_ _05787_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a31o_1
X_16377_ _08543_ _09225_ _09347_ vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19165_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__buf_2
X_20418__168 clknet_1_1__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__inv_2
X_13589_ _06757_ _06758_ _06759_ _06577_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__a22o_1
Xhold6309 net1976 vssd1 vssd1 vccd1 vccd1 net6836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18116_ net3732 _02343_ _02344_ _06057_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15328_ _07991_ _08404_ vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__nor2_2
X_19096_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5608 rbzero.spi_registers.new_texadd\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net6135
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5619 net1065 vssd1 vssd1 vccd1 vccd1 net6146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ _08353_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__inv_2
X_18047_ _02281_ _02282_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__xnor2_1
Xhold4907 net1025 vssd1 vssd1 vccd1 vccd1 net5434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4918 _00806_ vssd1 vssd1 vccd1 vccd1 net5445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4929 net1118 vssd1 vssd1 vccd1 vccd1 net5456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19998_ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18949_ net2759 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21960_ net402 net2434 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20911_ clknet_leaf_80_i_clk _00398_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_21891_ net333 net2606 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _09721_ clknet_1_0__leaf__05847_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__and2_2
XFILLER_0_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20773_ _03942_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7500 _02803_ vssd1 vssd1 vccd1 vccd1 net8027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7511 net3508 vssd1 vssd1 vccd1 vccd1 net8038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7522 _02564_ vssd1 vssd1 vccd1 vccd1 net8049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7533 _02879_ vssd1 vssd1 vccd1 vccd1 net8060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7544 net7999 vssd1 vssd1 vccd1 vccd1 net8071 sky130_fd_sc_hd__buf_1
Xhold6810 rbzero.tex_b1\[53\] vssd1 vssd1 vccd1 vccd1 net7337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7555 net4538 vssd1 vssd1 vccd1 vccd1 net8082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6821 net2728 vssd1 vssd1 vccd1 vccd1 net7348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7566 _02824_ vssd1 vssd1 vccd1 vccd1 net8093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6832 net3128 vssd1 vssd1 vccd1 vccd1 net7359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7577 rbzero.wall_tracer.rayAddendX\[-8\] vssd1 vssd1 vccd1 vccd1 net8104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6843 _04124_ vssd1 vssd1 vccd1 vccd1 net7370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7588 rbzero.spi_registers.texadd2\[19\] vssd1 vssd1 vccd1 vccd1 net8115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6854 net2533 vssd1 vssd1 vccd1 vccd1 net7381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7599 net960 vssd1 vssd1 vccd1 vccd1 net8126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6865 rbzero.tex_b0\[42\] vssd1 vssd1 vccd1 vccd1 net7392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21325_ clknet_leaf_45_i_clk net5143 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6876 net2959 vssd1 vssd1 vccd1 vccd1 net7403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6887 rbzero.tex_r0\[61\] vssd1 vssd1 vccd1 vccd1 net7414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6898 net2889 vssd1 vssd1 vccd1 vccd1 net7425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _01563_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
X_21256_ clknet_leaf_2_i_clk net3585 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold461 net4208 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _01323_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold483 net8014 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
X_20207_ net7188 _03743_ net4604 _03732_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__o211a_1
Xhold494 _03426_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
X_21187_ clknet_leaf_127_i_clk net3197 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20138_ rbzero.debug_overlay.facingX\[-3\] net1932 _03710_ vssd1 vssd1 vccd1 vccd1
+ _03720_ sky130_fd_sc_hd__mux2_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _08190_ _03610_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nor2_1
X_12960_ net3960 _06061_ _06135_ net4034 vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a22o_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 net6584 vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20523__263 clknet_1_0__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__inv_2
Xhold1161 net6648 vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ _05079_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and2b_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _01007_ vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 net5813 vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ net4748 vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__inv_2
Xhold1194 net6779 vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _07451_ _07799_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__nor2_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _04828_ _04930_ _05026_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14561_ _07696_ _07731_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__xnor2_2
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _04961_ _04962_ _04915_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__mux2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _08391_ _08411_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__nor2_1
X_13512_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__buf_6
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _10297_ _10298_ vssd1 vssd1 vccd1 vccd1 _10299_ sky130_fd_sc_hd__and2b_1
X_10724_ net2908 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__clkbuf_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _07618_ _07619_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__nor2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16231_ _09109_ _09081_ _09207_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13443_ _06531_ _06533_ _06438_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__a21o_1
X_10655_ net6653 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _09133_ _09254_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__nand2_1
X_13374_ _06540_ _06541_ _06542_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__o21a_2
XFILLER_0_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10586_ _04102_ _04021_ _04027_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__or3b_4
XFILLER_0_140_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15113_ _08200_ _08207_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__nor2_1
X_12325_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _05249_ vssd1 vssd1 vccd1 vccd1 _05511_
+ sky130_fd_sc_hd__mux2_1
X_16093_ _09030_ _09042_ _09186_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__a21oi_2
X_15044_ _08133_ _08135_ _08138_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__o21ai_4
X_19921_ net2801 net3227 _03561_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__mux2_1
X_12256_ _05441_ _05442_ _04910_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__mux2_1
X_11207_ net7202 net6673 _04423_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19852_ net3077 net7540 _03528_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__mux2_1
X_12187_ net7723 _05374_ net7570 vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__mux2_2
XFILLER_0_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18803_ net4814 net3940 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__and2b_1
X_11138_ net6973 net6746 _04390_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16995_ _10013_ _10014_ _09884_ net8383 vssd1 vssd1 vccd1 vccd1 _10016_ sky130_fd_sc_hd__o211ai_1
X_18734_ _02882_ net4807 net8061 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__o21ai_1
X_11069_ net2239 net5592 _04353_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__mux2_1
X_15946_ _08444_ net8033 _09040_ _08452_ _08434_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__o32a_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18665_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__nand2_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _08954_ _08971_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__and2_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _01777_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__and3_1
X_20498__240 clknet_1_0__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__inv_2
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14828_ _07839_ _07986_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__nor2_1
X_18596_ _02753_ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ _01786_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14759_ _07860_ _07849_ _07925_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_175_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17478_ _10144_ _10373_ _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19217_ net1432 _03169_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__or2_1
X_16429_ _09398_ _09501_ _09518_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__nand3_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6106 net1891 vssd1 vssd1 vccd1 vccd1 net6633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6117 _04220_ vssd1 vssd1 vccd1 vccd1 net6644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19148_ net4393 _03145_ net1831 _03149_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__o211a_1
Xhold6128 net1973 vssd1 vssd1 vccd1 vccd1 net6655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6139 _03597_ vssd1 vssd1 vccd1 vccd1 net6666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5405 rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 net5932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5416 net3623 vssd1 vssd1 vccd1 vccd1 net5943 sky130_fd_sc_hd__dlygate4sd3_1
X_19079_ net2436 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__clkbuf_1
Xhold5427 net3779 vssd1 vssd1 vccd1 vccd1 net5954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5438 net4065 vssd1 vssd1 vccd1 vccd1 net5965 sky130_fd_sc_hd__buf_2
Xhold4704 rbzero.spi_registers.texadd0\[15\] vssd1 vssd1 vccd1 vccd1 net5231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5449 _06159_ vssd1 vssd1 vccd1 vccd1 net5976 sky130_fd_sc_hd__dlygate4sd3_1
X_21110_ clknet_leaf_93_i_clk net3143 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4715 net800 vssd1 vssd1 vccd1 vccd1 net5242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4726 _01606_ vssd1 vssd1 vccd1 vccd1 net5253 sky130_fd_sc_hd__dlygate4sd3_1
X_22090_ net152 net2501 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4737 net860 vssd1 vssd1 vccd1 vccd1 net5264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4748 rbzero.spi_registers.texadd2\[17\] vssd1 vssd1 vccd1 vccd1 net5275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4759 net879 vssd1 vssd1 vccd1 vccd1 net5286 sky130_fd_sc_hd__dlygate4sd3_1
X_21041_ clknet_leaf_64_i_clk _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_106_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19779__58 clknet_1_0__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
XFILLER_0_198_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21943_ net385 net1654 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03510_ clknet_0__03510_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03510_
+ sky130_fd_sc_hd__clkbuf_16
X_21874_ net316 net2267 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _04485_ net4122 vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20756_ net984 net5448 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20687_ net6058 net4922 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__xnor2_1
Xhold7330 rbzero.wall_tracer.stepDistX\[-10\] vssd1 vssd1 vccd1 vccd1 net7857 sky130_fd_sc_hd__dlygate4sd3_1
X_20553__289 clknet_1_0__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__inv_2
X_10440_ net6039 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__clkbuf_8
Xhold7341 net3459 vssd1 vssd1 vccd1 vccd1 net7868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7352 rbzero.wall_tracer.stepDistY\[4\] vssd1 vssd1 vccd1 vccd1 net7879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7363 rbzero.traced_texVinit\[1\] vssd1 vssd1 vccd1 vccd1 net7890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7374 net1101 vssd1 vssd1 vccd1 vccd1 net7901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6640 net2282 vssd1 vssd1 vccd1 vccd1 net7167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7385 _00500_ vssd1 vssd1 vccd1 vccd1 net7912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7396 net968 vssd1 vssd1 vccd1 vccd1 net7923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6651 net2069 vssd1 vssd1 vccd1 vccd1 net7178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6662 rbzero.tex_g0\[33\] vssd1 vssd1 vccd1 vccd1 net7189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6673 net2444 vssd1 vssd1 vccd1 vccd1 net7200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6684 rbzero.tex_g0\[2\] vssd1 vssd1 vccd1 vccd1 net7211 sky130_fd_sc_hd__dlygate4sd3_1
X_12110_ net4964 net7722 _04845_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__mux2_1
Xhold5950 rbzero.tex_g1\[18\] vssd1 vssd1 vccd1 vccd1 net6477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21308_ clknet_leaf_8_i_clk net5246 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6695 net2625 vssd1 vssd1 vccd1 vccd1 net7222 sky130_fd_sc_hd__dlygate4sd3_1
X_13090_ _06244_ _06260_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__or2_1
Xhold5961 net1520 vssd1 vssd1 vccd1 vccd1 net6488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5972 rbzero.tex_g0\[10\] vssd1 vssd1 vccd1 vccd1 net6499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5983 net1459 vssd1 vssd1 vccd1 vccd1 net6510 sky130_fd_sc_hd__dlygate4sd3_1
X_12041_ rbzero.tex_r1\[19\] rbzero.tex_r1\[18\] _04979_ vssd1 vssd1 vccd1 vccd1 _05230_
+ sky130_fd_sc_hd__mux2_1
Xhold5994 _03447_ vssd1 vssd1 vccd1 vccd1 net6521 sky130_fd_sc_hd__dlygate4sd3_1
X_21239_ clknet_leaf_45_i_clk net4042 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold280 net5245 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 net5247 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15800_ _08885_ _08888_ _08889_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__a21o_1
X_20447__194 clknet_1_0__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_70_i_clk clknet_4_13__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16780_ _06058_ _09808_ _09810_ vssd1 vssd1 vccd1 vccd1 _09811_ sky130_fd_sc_hd__o21ai_1
X_13992_ _07114_ _07162_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__xnor2_1
X_15731_ _08824_ _08825_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12943_ _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__clkbuf_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ net4603 net3509 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__nor2_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _08657_ _08703_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__or2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _06034_ _06047_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__o21a_1
XFILLER_0_201_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _10407_ _10418_ vssd1 vssd1 vccd1 vccd1 _10419_ sky130_fd_sc_hd__xnor2_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11825_ net3648 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__inv_2
X_14613_ _07558_ _07606_ _07608_ _07780_ _07783_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__a32o_2
XFILLER_0_201_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15593_ _08676_ _08677_ _08687_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__nand3_1
X_18381_ net4501 net4733 _05155_ _02524_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__o31a_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17332_ _10347_ _10350_ vssd1 vssd1 vccd1 vccd1 _10351_ sky130_fd_sc_hd__xnor2_2
X_14544_ _07713_ _07714_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _04930_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ net2662 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__clkbuf_1
X_17263_ _10279_ _10280_ vssd1 vssd1 vccd1 vccd1 _10282_ sky130_fd_sc_hd__nor2_1
X_14475_ _07628_ _07645_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__xor2_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ net3405 net3954 _04870_ _04462_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19002_ net5764 net4454 _02992_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16214_ _09285_ _09306_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13426_ _06450_ net82 _06525_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__or3_1
X_10638_ net6916 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__clkbuf_1
X_17194_ _10212_ _10213_ vssd1 vssd1 vccd1 vccd1 _10214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _09236_ _09237_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13357_ net82 _06525_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nor2_2
XFILLER_0_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10569_ net2525 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _05239_ vssd1 vssd1 vccd1 vccd1 _05494_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16076_ _08181_ _08450_ _09169_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_23_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13288_ _06456_ _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xor2_4
X_19904_ net3321 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
X_15027_ net4083 net3627 _06117_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__and3_1
X_12239_ _05424_ _05425_ _04847_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2609 _01133_ vssd1 vssd1 vccd1 vccd1 net3136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19835_ net3026 net3019 _03517_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
Xhold1908 net7276 vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1919 _01520_ vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_38_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19766_ clknet_1_1__leaf__03506_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__buf_1
XFILLER_0_194_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16978_ _09893_ _09999_ vssd1 vssd1 vccd1 vccd1 _10000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
X_18717_ net4709 net3575 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nor2_1
X_15929_ _09016_ _09023_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19697_ net6349 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18648_ net4528 net4635 _05164_ _02767_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__o31a_1
XFILLER_0_189_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18579_ net7702 net3999 net4648 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21590_ net224 net2514 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20472_ clknet_1_0__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5202 rbzero.tex_r1\[16\] vssd1 vssd1 vccd1 vccd1 net5729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5213 _01619_ vssd1 vssd1 vccd1 vccd1 net5740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5224 _03670_ vssd1 vssd1 vccd1 vccd1 net5751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5235 net3470 vssd1 vssd1 vccd1 vccd1 net5762 sky130_fd_sc_hd__dlygate4sd3_1
X_22142_ clknet_leaf_40_i_clk _01629_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold4501 rbzero.spi_registers.texadd1\[7\] vssd1 vssd1 vccd1 vccd1 net5028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5246 _01189_ vssd1 vssd1 vccd1 vccd1 net5773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5257 net7691 vssd1 vssd1 vccd1 vccd1 net5784 sky130_fd_sc_hd__buf_1
Xhold4512 net704 vssd1 vssd1 vccd1 vccd1 net5039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4523 _00889_ vssd1 vssd1 vccd1 vccd1 net5050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5268 _02819_ vssd1 vssd1 vccd1 vccd1 net5795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5279 _00627_ vssd1 vssd1 vccd1 vccd1 net5806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4534 net826 vssd1 vssd1 vccd1 vccd1 net5061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3800 rbzero.pov.ready_buffer\[50\] vssd1 vssd1 vccd1 vccd1 net4327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4545 rbzero.spi_registers.texadd2\[8\] vssd1 vssd1 vccd1 vccd1 net5072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3811 net3715 vssd1 vssd1 vccd1 vccd1 net4338 sky130_fd_sc_hd__dlygate4sd3_1
X_22073_ net515 net2983 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4556 net712 vssd1 vssd1 vccd1 vccd1 net5083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3822 net891 vssd1 vssd1 vccd1 vccd1 net4349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4567 _00783_ vssd1 vssd1 vccd1 vccd1 net5094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3833 net3686 vssd1 vssd1 vccd1 vccd1 net4360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4578 net795 vssd1 vssd1 vccd1 vccd1 net5105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3844 net1178 vssd1 vssd1 vccd1 vccd1 net4371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4589 rbzero.spi_registers.texadd2\[6\] vssd1 vssd1 vccd1 vccd1 net5116 sky130_fd_sc_hd__dlygate4sd3_1
X_21024_ clknet_leaf_63_i_clk net4301 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3855 net7866 vssd1 vssd1 vccd1 vccd1 net4382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3866 net8169 vssd1 vssd1 vccd1 vccd1 net4393 sky130_fd_sc_hd__clkbuf_2
Xhold3877 net7902 vssd1 vssd1 vccd1 vccd1 net4404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3888 net8038 vssd1 vssd1 vccd1 vccd1 net4415 sky130_fd_sc_hd__buf_1
Xhold3899 net653 vssd1 vssd1 vccd1 vccd1 net4426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21926_ net368 net632 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21857_ net299 net2859 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _04787_ _04796_ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o21a_1
X_20808_ _03969_ _03970_ _03971_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__o21a_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ net46 _05763_ _05745_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a21bo_1
X_21788_ clknet_leaf_20_i_clk net1592 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_20635__364 clknet_1_0__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__inv_2
X_11541_ net2587 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__inv_2
X_20739_ net896 net5376 vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14260_ _07395_ _07408_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o21ai_1
X_11472_ net3995 net4065 net4091 net3 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__or4b_1
XFILLER_0_163_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ _06303_ _06304_ _06306_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__a21o_1
Xhold7160 net3959 vssd1 vssd1 vccd1 vccd1 net7687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7171 net2953 vssd1 vssd1 vccd1 vccd1 net7698 sky130_fd_sc_hd__dlymetal6s2s_1
X_14191_ _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__nand2_1
Xhold7182 gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 net7709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7193 _05464_ vssd1 vssd1 vccd1 vccd1 net7720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6470 net2168 vssd1 vssd1 vccd1 vccd1 net6997 sky130_fd_sc_hd__dlygate4sd3_1
X_13142_ _06281_ _06312_ _06279_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a21o_1
Xhold6481 rbzero.tex_r0\[53\] vssd1 vssd1 vccd1 vccd1 net7008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6492 net2043 vssd1 vssd1 vccd1 vccd1 net7019 sky130_fd_sc_hd__dlygate4sd3_1
X_17950_ _02068_ _02092_ _02185_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__nand3_1
X_13073_ net5428 _06244_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__and2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5780 net1435 vssd1 vssd1 vccd1 vccd1 net6307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5791 _03834_ vssd1 vssd1 vccd1 vccd1 net6318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16901_ _09921_ _09922_ vssd1 vssd1 vccd1 vccd1 _09923_ sky130_fd_sc_hd__nor2_1
X_12024_ _04829_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__buf_4
X_17881_ _10432_ _09114_ _02117_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19620_ net6448 net4016 _03430_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
X_16832_ _09857_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__clkbuf_1
X_20380__134 clknet_1_1__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__inv_2
X_19551_ net2224 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
X_19758__39 clknet_1_0__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
X_16763_ _09795_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13975_ _07144_ _07145_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18502_ _02677_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__xnor2_1
X_15714_ _08805_ _08808_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__and2_2
X_19482_ net1481 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
X_12926_ net4779 net4643 _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__and3_1
X_16694_ net984 _09743_ _09744_ net8029 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18433_ _02601_ _02613_ _02612_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _08735_ _08739_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__nand2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ net7776 vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__inv_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _04978_ vssd1 vssd1 vccd1 vccd1 _04998_
+ sky130_fd_sc_hd__mux2_1
X_18364_ net4501 _02540_ _04480_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a21oi_1
X_15576_ _08669_ _08670_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _05961_ _05962_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _10314_ _10315_ _10332_ vssd1 vssd1 vccd1 vccd1 _10334_ sky130_fd_sc_hd__nand3_1
X_11739_ _04922_ _04925_ _04927_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14527_ _07665_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18295_ net6407 net3596 _02493_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17246_ _10262_ _10263_ _10136_ _10140_ vssd1 vssd1 vccd1 vccd1 _10265_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _07621_ _07617_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ _06531_ _06533_ _06450_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a21oi_1
X_17177_ _10195_ _10196_ vssd1 vssd1 vccd1 vccd1 _10197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14389_ _07531_ _07553_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16128_ _09152_ _09130_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _09130_ _09152_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__xnor2_1
Xhold3118 _03330_ vssd1 vssd1 vccd1 vccd1 net3645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3129 net7729 vssd1 vssd1 vccd1 vccd1 net3656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2406 rbzero.pov.spi_buffer\[38\] vssd1 vssd1 vccd1 vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2417 net7410 vssd1 vssd1 vccd1 vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2428 _00933_ vssd1 vssd1 vccd1 vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2439 _04237_ vssd1 vssd1 vccd1 vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1705 net6023 vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
X_19818_ net2312 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__clkbuf_4
Xhold1716 net4478 vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1727 _04328_ vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 net6935 vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 _01300_ vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21711_ clknet_leaf_109_i_clk net4479 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21642_ clknet_leaf_116_i_clk net3262 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21573_ net207 net1931 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_20 rbzero.wall_tracer.visualWallDist\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_42 net4751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_75 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_86 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5010 _00765_ vssd1 vssd1 vccd1 vccd1 net5537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5021 _04071_ vssd1 vssd1 vccd1 vccd1 net5548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5032 _04101_ vssd1 vssd1 vccd1 vccd1 net5559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5043 net1764 vssd1 vssd1 vccd1 vccd1 net5570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5054 net1616 vssd1 vssd1 vccd1 vccd1 net5581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5065 rbzero.tex_b1\[28\] vssd1 vssd1 vccd1 vccd1 net5592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4320 rbzero.wall_tracer.rayAddendY\[-6\] vssd1 vssd1 vccd1 vccd1 net4847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5076 net2794 vssd1 vssd1 vccd1 vccd1 net5603 sky130_fd_sc_hd__dlygate4sd3_1
X_22125_ clknet_leaf_54_i_clk net5494 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold4331 _02909_ vssd1 vssd1 vccd1 vccd1 net4858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4342 _02671_ vssd1 vssd1 vccd1 vccd1 net4869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5087 _03155_ vssd1 vssd1 vccd1 vccd1 net5614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5098 rbzero.tex_b0\[2\] vssd1 vssd1 vccd1 vccd1 net5625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4353 _01653_ vssd1 vssd1 vccd1 vccd1 net4880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4364 net7817 vssd1 vssd1 vccd1 vccd1 net4891 sky130_fd_sc_hd__clkbuf_2
Xhold3630 _08094_ vssd1 vssd1 vccd1 vccd1 net4157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4375 _03685_ vssd1 vssd1 vccd1 vccd1 net4902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4386 _09343_ vssd1 vssd1 vccd1 vccd1 net4913 sky130_fd_sc_hd__clkbuf_2
X_22056_ net498 net1066 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold3641 net3386 vssd1 vssd1 vccd1 vccd1 net4168 sky130_fd_sc_hd__buf_4
Xhold4397 net603 vssd1 vssd1 vccd1 vccd1 net4924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3652 _03804_ vssd1 vssd1 vccd1 vccd1 net4179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3663 _09713_ vssd1 vssd1 vccd1 vccd1 net4190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3674 net7884 vssd1 vssd1 vccd1 vccd1 net4201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2940 net8382 vssd1 vssd1 vccd1 vccd1 net3467 sky130_fd_sc_hd__dlygate4sd3_1
X_21007_ clknet_leaf_37_i_clk net4323 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3685 net7896 vssd1 vssd1 vccd1 vccd1 net4212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3696 net7908 vssd1 vssd1 vccd1 vccd1 net4223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2951 net7578 vssd1 vssd1 vccd1 vccd1 net3478 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2962 net8219 vssd1 vssd1 vccd1 vccd1 net3489 sky130_fd_sc_hd__clkbuf_4
Xhold2973 net5797 vssd1 vssd1 vccd1 vccd1 net3500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2984 _03758_ vssd1 vssd1 vccd1 vccd1 net3511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2995 _00917_ vssd1 vssd1 vccd1 vccd1 net3522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ _06702_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__inv_2
X_10972_ net6500 net2670 _04298_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21909_ net351 net2925 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap77 _06722_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_2
X_12711_ net32 net33 _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__and3b_1
XFILLER_0_168_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap88 _04846_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_2
X_13691_ _06852_ _06861_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15430_ _08280_ _08323_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ net4066 _05798_ _05817_ net71 _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20559__295 clknet_1_1__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__inv_2
XFILLER_0_155_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _08454_ _08444_ net8033 _08427_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__or4b_4
X_12573_ net4149 net4141 net4164 net7727 _05749_ net19 vssd1 vssd1 vccd1 vccd1 _05753_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ _09930_ _09996_ _09994_ vssd1 vssd1 vccd1 vccd1 _10121_ sky130_fd_sc_hd__a21oi_2
X_14312_ _07424_ _07423_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__and2b_1
X_11524_ _04464_ net4152 net4306 _04682_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a2bb2o_1
X_15292_ _08161_ _08368_ _08386_ _08180_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__a2bb2o_1
X_18080_ _02315_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17031_ _10049_ _10050_ vssd1 vssd1 vccd1 vccd1 _10052_ sky130_fd_sc_hd__and2_1
X_14243_ _07310_ _07344_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11455_ _04629_ _04646_ _04494_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14174_ _07343_ _07344_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11386_ rbzero.spi_registers.texadd0\[23\] vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__inv_2
X_13125_ _06278_ _06292_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18982_ net6239 net5816 _03058_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _02168_ _02169_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__nand2_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _06197_ _06199_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ net4138 _04460_ _05191_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__o211a_1
X_17864_ _02100_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19603_ net1031 net4835 _03312_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__a21oi_1
X_16815_ net4508 net4383 vssd1 vssd1 vccd1 vccd1 _09842_ sky130_fd_sc_hd__nand2_1
X_17795_ _02013_ _02033_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19534_ net1765 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
X_16746_ _09779_ _09780_ vssd1 vssd1 vccd1 vccd1 _09781_ sky130_fd_sc_hd__xnor2_1
X_13958_ _07117_ _07127_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19465_ net1622 net5994 _03345_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
X_12909_ _06084_ net3884 net2379 net2006 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a211o_1
XFILLER_0_186_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16677_ net4259 _09741_ _09742_ net1154 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13889_ _07057_ _07059_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18416_ _02596_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__xnor2_1
X_15628_ _08720_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__nand2_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18347_ _02526_ _02527_ _02528_ _02533_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a32o_1
X_15559_ _08625_ _08649_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7907 _08149_ vssd1 vssd1 vccd1 vccd1 net8434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ net1242 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17229_ _10246_ _10248_ vssd1 vssd1 vccd1 vccd1 _10249_ sky130_fd_sc_hd__xor2_4
Xinput40 i_mode[0] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_6
XFILLER_0_25_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput51 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_8
Xclkbuf_1_1__f__03867_ clknet_0__03867_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03867_
+ sky130_fd_sc_hd__clkbuf_16
Xhold802 net6302 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20240_ net3996 net4128 _05050_ _05730_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__and4bb_1
Xhold813 net6274 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold824 _01001_ vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 net6316 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _00588_ vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 net6555 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20171_ rbzero.debug_overlay.facingY\[-2\] net3711 _03723_ vssd1 vssd1 vccd1 vccd1
+ _03741_ sky130_fd_sc_hd__mux2_1
Xhold868 net4027 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _03445_ vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2203 _01485_ vssd1 vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 net5729 vssd1 vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2225 _01450_ vssd1 vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2236 _01475_ vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1502 net6749 vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2247 net7294 vssd1 vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2258 _01422_ vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 net2789 vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 net7349 vssd1 vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 _01465_ vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _00909_ vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1546 net6933 vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _01084_ vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1568 _04139_ vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1579 _00949_ vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21625_ clknet_leaf_128_i_clk net1690 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21556_ net190 net2481 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21487_ clknet_leaf_47_i_clk net1280 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11240_ net2893 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20438_ clknet_1_0__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11171_ net7417 net7393 _04401_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__mux2_1
Xhold4150 net3381 vssd1 vssd1 vccd1 vccd1 net4677 sky130_fd_sc_hd__dlygate4sd3_1
X_22108_ net146 net2550 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4161 _01236_ vssd1 vssd1 vccd1 vccd1 net4688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4172 _03759_ vssd1 vssd1 vccd1 vccd1 net4699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4183 _03779_ vssd1 vssd1 vccd1 vccd1 net4710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4194 net627 vssd1 vssd1 vccd1 vccd1 net4721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3460 _08105_ vssd1 vssd1 vccd1 vccd1 net3987 sky130_fd_sc_hd__dlygate4sd3_1
X_22039_ net481 net2203 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
Xhold3471 rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 net3998 sky130_fd_sc_hd__dlygate4sd3_1
X_14930_ net8467 _06237_ _04482_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__o21a_1
Xhold3482 _06132_ vssd1 vssd1 vccd1 vccd1 net4009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3493 net7692 vssd1 vssd1 vccd1 vccd1 net4020 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2770 rbzero.pov.spi_buffer\[35\] vssd1 vssd1 vccd1 vccd1 net3297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2781 net5924 vssd1 vssd1 vccd1 vccd1 net3308 sky130_fd_sc_hd__dlygate4sd3_1
X_14861_ _06545_ _07960_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__a21o_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2792 rbzero.pov.spi_buffer\[39\] vssd1 vssd1 vccd1 vccd1 net3319 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _09663_ _09688_ _09689_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__and3_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13812_ _06954_ _06958_ _06959_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__nor3_1
X_17580_ _01819_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__nand2_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _07954_ _07955_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ _09504_ _09616_ _09620_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__a21oi_1
X_10955_ _04264_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__clkbuf_4
X_13743_ net571 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19250_ net6417 _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__or2_1
X_16462_ _08446_ _09552_ _09420_ _09421_ _09412_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ net2576 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__clkbuf_1
X_13674_ _06729_ _06721_ _06839_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18201_ net3669 net4459 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20492__235 clknet_1_0__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__inv_2
X_15413_ _08186_ _08244_ _08246_ _08243_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ net25 vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__inv_2
X_19181_ net5185 _03168_ _03177_ _03176_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__o211a_1
X_16393_ _09480_ _09482_ _09479_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18132_ net8039 _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12556_ _05729_ _05736_ net11 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__mux2_1
X_15344_ _07991_ _07998_ _08004_ _08404_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__or4_4
XFILLER_0_108_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11507_ net4102 _04692_ _04695_ _04495_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a221o_1
X_18063_ _01784_ _09666_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ net8497 _06364_ net4181 vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__mux2_1
X_12487_ net43 _05646_ _05642_ net46 vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a22o_1
X_17014_ _08543_ _09472_ _09899_ _09897_ vssd1 vssd1 vccd1 vccd1 _10035_ sky130_fd_sc_hd__o31a_1
Xhold109 net6815 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ _07241_ _07282_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__and2_1
X_11438_ rbzero.spi_registers.texadd0\[3\] rbzero.spi_registers.texadd0\[2\] _04020_
+ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _06696_ _07323_ _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11369_ _04558_ _04559_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13108_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__and2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _06695_ _06729_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__and2b_1
X_18965_ net3052 net7567 net2874 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17916_ _02150_ _02153_ net90 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a21oi_1
X_13039_ _06212_ net3669 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ net6125 net2364 _03014_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__mux2_1
X_17847_ _02083_ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _01784_ _09181_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19517_ net1396 net5540 net3086 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16729_ net4647 _08035_ vssd1 vssd1 vccd1 vccd1 _09767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ net1033 _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ net5153 _03283_ _03292_ _03288_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21410_ clknet_leaf_38_i_clk net4314 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7704 rbzero.traced_texa\[-8\] vssd1 vssd1 vccd1 vccd1 net8231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7715 _02904_ vssd1 vssd1 vccd1 vccd1 net8242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7726 rbzero.debug_overlay.vplaneX\[-7\] vssd1 vssd1 vccd1 vccd1 net8253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7737 net7832 vssd1 vssd1 vccd1 vccd1 net8264 sky130_fd_sc_hd__clkbuf_2
Xhold7748 net8088 vssd1 vssd1 vccd1 vccd1 net8275 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21341_ clknet_leaf_20_i_clk net5039 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold610 net5461 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
X_21272_ clknet_leaf_24_i_clk net4349 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold621 net6214 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 net6250 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20223_ net3575 net1970 _03709_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__mux2_1
Xhold643 _00660_ vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold654 _01410_ vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold665 net6244 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 net6596 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold687 net6264 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 net6270 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ net3688 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
Xhold2000 net7106 vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2011 _01284_ vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2022 _04034_ vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2033 net6998 vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2044 _01441_ vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
X_20085_ _08301_ _03631_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 net5567 vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2055 net5578 vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 net6668 vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2066 _04170_ vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2077 net7422 vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1332 net6557 vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1343 net6666 vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2088 _01660_ vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1354 _03397_ vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2099 _04147_ vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1365 net6634 vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1376 net6726 vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1387 _01554_ vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1398 _00977_ vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20987_ clknet_leaf_113_i_clk net3958 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10740_ net6615 net6910 _04182_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ net2092 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ rbzero.tex_b1\[47\] rbzero.tex_b1\[46\] _04924_ vssd1 vssd1 vccd1 vccd1 _05595_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21608_ clknet_leaf_132_i_clk net1858 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _06394_ net82 _06525_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__or3_1
X_12341_ _04922_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21539_ net173 net1945 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ _06416_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12272_ _05040_ _05455_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_209_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14011_ _07179_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__xnor2_1
X_11223_ net7127 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__clkbuf_1
X_11154_ net7206 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18750_ _02869_ _02887_ _02889_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
X_15962_ _08561_ _08541_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__or2b_1
X_11085_ net6848 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17701_ _01831_ _01833_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3290 _03087_ vssd1 vssd1 vccd1 vccd1 net3817 sky130_fd_sc_hd__dlygate4sd3_1
X_14913_ _08035_ vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__clkbuf_4
X_18681_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__xor2_1
X_15893_ _08761_ _08987_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__xnor2_4
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _10190_ _09116_ _01765_ _01763_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__o31ai_2
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ _07839_ _07986_ net7846 vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__o21ai_2
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17563_ _01802_ _01803_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14775_ _07899_ _07900_ net7813 vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ net4154 _04747_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__nand2_1
X_20500__242 clknet_1_0__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__inv_2
X_19302_ net1508 _03238_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__or2_1
X_16514_ _09479_ _09603_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13726_ _06885_ _06896_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__xnor2_2
X_10938_ net2723 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
X_17494_ _10385_ _10386_ _10383_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19233_ net5125 _03201_ _03208_ _03206_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__o211a_1
X_16445_ _09534_ _09535_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__nand2_1
X_10869_ net7133 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__clkbuf_1
X_13657_ _06807_ _06821_ _06805_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19164_ net3842 _03140_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__and2_1
X_12608_ _05746_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__inv_2
X_16376_ _09372_ _09388_ _09466_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__a21bo_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13588_ net78 _06634_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_186_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18115_ _02343_ _02344_ net3732 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15327_ _07989_ _07937_ _07997_ _07868_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_147_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19095_ net3623 _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__and2_1
X_12539_ _05708_ _05717_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5609 net1399 vssd1 vssd1 vccd1 vccd1 net6136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18046_ _09040_ _09114_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15258_ _08144_ _08352_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4908 rbzero.spi_registers.texadd0\[22\] vssd1 vssd1 vccd1 vccd1 net5435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4919 net1068 vssd1 vssd1 vccd1 vccd1 net5446 sky130_fd_sc_hd__dlygate4sd3_1
X_14209_ _07370_ _07379_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nor2_1
X_15189_ _08269_ _08283_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__or2b_1
X_19997_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__buf_2
X_18948_ net7178 net3440 _03036_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
X_18879_ net2869 net7409 _03003_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20910_ clknet_leaf_81_i_clk _00397_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21890_ net332 net2565 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20841_ _03997_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20772_ _03937_ _03940_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7501 _00628_ vssd1 vssd1 vccd1 vccd1 net8028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7512 _02357_ vssd1 vssd1 vccd1 vccd1 net8039 sky130_fd_sc_hd__buf_1
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7523 _00600_ vssd1 vssd1 vccd1 vccd1 net8050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7534 _02881_ vssd1 vssd1 vccd1 vccd1 net8061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6800 rbzero.tex_r1\[49\] vssd1 vssd1 vccd1 vccd1 net7327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7545 _08140_ vssd1 vssd1 vccd1 vccd1 net8072 sky130_fd_sc_hd__buf_1
Xhold6811 net2545 vssd1 vssd1 vccd1 vccd1 net7338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6822 rbzero.tex_r1\[30\] vssd1 vssd1 vccd1 vccd1 net7349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7567 _02825_ vssd1 vssd1 vccd1 vccd1 net8094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6833 rbzero.tex_g0\[23\] vssd1 vssd1 vccd1 vccd1 net7360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7578 net693 vssd1 vssd1 vccd1 vccd1 net8105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6844 net2611 vssd1 vssd1 vccd1 vccd1 net7371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7589 net4195 vssd1 vssd1 vccd1 vccd1 net8116 sky130_fd_sc_hd__dlygate4sd3_1
X_21324_ clknet_leaf_45_i_clk net5099 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6855 rbzero.tex_b1\[18\] vssd1 vssd1 vccd1 vccd1 net7382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6866 net2813 vssd1 vssd1 vccd1 vccd1 net7393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6877 rbzero.tex_b0\[54\] vssd1 vssd1 vccd1 vccd1 net7404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6888 net2914 vssd1 vssd1 vccd1 vccd1 net7415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6899 rbzero.tex_g1\[53\] vssd1 vssd1 vccd1 vccd1 net7426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 net8234 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_1
X_21255_ clknet_leaf_3_i_clk net3483 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold451 net5351 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 net5411 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
X_20206_ net4603 _03744_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or2_1
Xhold473 net5343 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 net5387 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
X_21186_ clknet_leaf_102_i_clk net1917 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold495 net4817 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20137_ net3692 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ net5859 _03660_ _03668_ _03628_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__o211a_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 _01009_ vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 _02497_ vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 _03546_ vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net4105 _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nor2_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1173 net5534 vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ net3682 net4007 _06043_ net4436 _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a221o_1
Xhold1184 _00713_ vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 net6781 vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _05028_ _05030_ net4321 vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a21oi_2
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _04923_ vssd1 vssd1 vccd1 vccd1 _04962_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14560_ _07691_ _07698_ _07730_ _07694_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__and4_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10723_ net2907 net50 _04097_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
X_13511_ _06663_ _06673_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a21bo_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ _07660_ _07661_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__nand2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _09321_ _09322_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__nand2_4
XFILLER_0_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ net6651 net2405 _04138_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__mux2_1
X_13442_ net561 net560 _06406_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _08535_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13373_ net7833 _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nor2_2
X_10585_ _04028_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__inv_6
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15112_ _08206_ vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__buf_2
X_12324_ _05508_ _05509_ _04984_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__mux2_1
X_16092_ _09039_ _09041_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12255_ rbzero.tex_g1\[63\] rbzero.tex_g1\[62\] _04933_ vssd1 vssd1 vccd1 vccd1 _05442_
+ sky130_fd_sc_hd__mux2_1
X_15043_ net4381 _08119_ _08137_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19920_ net1886 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ net2963 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19851_ net2808 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
X_12186_ _04909_ _05333_ _05368_ _05373_ _05017_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__a32o_1
XFILLER_0_208_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11137_ net6028 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
X_18802_ net5863 net7496 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__and2b_2
X_16994_ _09884_ net8383 _10013_ _10014_ vssd1 vssd1 vccd1 vccd1 _10015_ sky130_fd_sc_hd__a211o_1
X_18733_ net8061 _02882_ net4807 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__or3_1
X_11068_ net5651 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
X_15945_ _08181_ _08450_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__nand2_4
XFILLER_0_204_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18664_ net5796 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__clkbuf_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _08951_ _08956_ _08970_ _08969_ _08968_ vssd1 vssd1 vccd1 vccd1 _08971_ sky130_fd_sc_hd__a32o_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _01777_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14827_ _07860_ _07837_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__nor2_1
X_18595_ net4424 net4599 _02753_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nand3b_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17546_ _10316_ _08616_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14758_ _07818_ _07861_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13709_ _06878_ _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17477_ _10371_ _10372_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14689_ _07818_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19216_ net5348 _03167_ _03196_ _03189_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__o211a_1
X_16428_ _09398_ _09501_ _09518_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6107 _04313_ vssd1 vssd1 vccd1 vccd1 net6634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19147_ net1830 _03147_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16359_ net8207 net8214 _08111_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__mux2_1
Xhold6118 net1653 vssd1 vssd1 vccd1 vccd1 net6645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6129 rbzero.tex_b1\[25\] vssd1 vssd1 vccd1 vccd1 net6656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5406 net3848 vssd1 vssd1 vccd1 vccd1 net5933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19078_ net43 net7277 _03109_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
Xhold5417 _03385_ vssd1 vssd1 vccd1 vccd1 net5944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5428 net3611 vssd1 vssd1 vccd1 vccd1 net5955 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5439 _05730_ vssd1 vssd1 vccd1 vccd1 net5966 sky130_fd_sc_hd__buf_1
X_18029_ _02160_ _02184_ _02161_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4705 net870 vssd1 vssd1 vccd1 vccd1 net5232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4716 rbzero.spi_registers.texadd0\[12\] vssd1 vssd1 vccd1 vccd1 net5243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4727 net867 vssd1 vssd1 vccd1 vccd1 net5254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4738 _00807_ vssd1 vssd1 vccd1 vccd1 net5265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21040_ clknet_leaf_56_i_clk net5330 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4749 net898 vssd1 vssd1 vccd1 vccd1 net5276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20507__248 clknet_1_1__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__inv_2
XFILLER_0_119_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21942_ net384 net2998 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21873_ net315 net1741 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20824_ net4083 net3452 _04485_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_210_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20755_ _03878_ _03928_ net8197 _03883_ net4980 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20686_ net4922 net63 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__nor2_1
Xhold7320 rbzero.wall_tracer.stepDistY\[6\] vssd1 vssd1 vccd1 vccd1 net7847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7331 net4534 vssd1 vssd1 vccd1 vccd1 net7858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7342 rbzero.wall_tracer.stepDistY\[-11\] vssd1 vssd1 vccd1 vccd1 net7869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7353 net4458 vssd1 vssd1 vccd1 vccd1 net7880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7364 net4205 vssd1 vssd1 vccd1 vccd1 net7891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6630 net2208 vssd1 vssd1 vccd1 vccd1 net7157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7375 rbzero.wall_tracer.stepDistX\[3\] vssd1 vssd1 vccd1 vccd1 net7902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6641 _04273_ vssd1 vssd1 vccd1 vccd1 net7168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7386 net4243 vssd1 vssd1 vccd1 vccd1 net7913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6652 rbzero.tex_g1\[36\] vssd1 vssd1 vccd1 vccd1 net7179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6663 net2616 vssd1 vssd1 vccd1 vccd1 net7190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6674 rbzero.tex_b0\[26\] vssd1 vssd1 vccd1 vccd1 net7201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21307_ clknet_leaf_10_i_clk net5294 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6685 net655 vssd1 vssd1 vccd1 vccd1 net7212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5940 _04191_ vssd1 vssd1 vccd1 vccd1 net6467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold5951 net1257 vssd1 vssd1 vccd1 vccd1 net6478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6696 rbzero.tex_r0\[30\] vssd1 vssd1 vccd1 vccd1 net7223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5962 _04155_ vssd1 vssd1 vccd1 vccd1 net6489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5973 net1272 vssd1 vssd1 vccd1 vccd1 net6500 sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ rbzero.tex_r1\[17\] rbzero.tex_r1\[16\] _04838_ vssd1 vssd1 vccd1 vccd1 _05229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21238_ clknet_leaf_45_i_clk net4018 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5984 rbzero.pov.spi_buffer\[23\] vssd1 vssd1 vccd1 vccd1 net6511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold270 net5108 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5995 net1812 vssd1 vssd1 vccd1 vccd1 net6522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 net5172 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 net5249 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
X_21169_ clknet_leaf_132_i_clk net2958 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13991_ _07160_ _07161_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__or2_1
X_15730_ _08326_ _08691_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__nor2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _04485_ _06117_ net3773 vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__and3b_2
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _08653_ _08755_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__nand2_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _06048_ _06028_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _10416_ _10417_ vssd1 vssd1 vccd1 vccd1 _10418_ sky130_fd_sc_hd__nor2_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__inv_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ net4080 vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__inv_2
X_18380_ net8047 net4784 _02560_ _02554_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a211o_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08683_ _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__xnor2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _10348_ _10349_ vssd1 vssd1 vccd1 vccd1 _10350_ sky130_fd_sc_hd__nand2_2
XFILLER_0_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07489_ _07198_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__nor2_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11755_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _04923_ vssd1 vssd1 vccd1 vccd1 _04945_
+ sky130_fd_sc_hd__mux2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17262_ _10279_ _10280_ vssd1 vssd1 vccd1 vccd1 _10281_ sky130_fd_sc_hd__and2_1
X_10706_ net7285 net2661 _04160_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ _07630_ _07643_ _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11686_ _04855_ _04872_ _04873_ _04875_ net3954 vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__o32a_1
X_19001_ net5793 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16213_ _09303_ _09305_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__xnor2_2
X_13425_ _06592_ _06595_ _06557_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ net6914 net2043 _04127_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__mux2_1
X_17193_ _10211_ _09664_ _10096_ _08918_ vssd1 vssd1 vccd1 vccd1 _10213_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20612__343 clknet_1_1__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__inv_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _09134_ _09229_ _09235_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__nand3_1
X_10568_ net6607 net7266 _04086_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _06516_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _04930_ _05492_ net86 vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__o21a_1
X_16075_ net3726 _08128_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__and2_1
X_10499_ net5788 net7063 _04053_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__mux2_1
X_13287_ _06457_ _06385_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nor2_2
X_19903_ net3320 net3214 _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__mux2_1
X_15026_ _07892_ net8403 _08114_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__mux2_2
X_12238_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _04968_ vssd1 vssd1 vccd1 vccd1 _05425_
+ sky130_fd_sc_hd__mux2_1
X_12169_ _04910_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__or2_1
X_19834_ net2263 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
Xhold1909 _03112_ vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
X_16977_ _09997_ _09998_ vssd1 vssd1 vccd1 vccd1 _09999_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
X_15928_ _09017_ _09022_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18716_ _02864_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__xnor2_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19696_ net6347 net3556 _03468_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18647_ _02801_ net8025 net4771 _02794_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _08947_ _08953_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18578_ net7701 _02741_ _02245_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17529_ _01768_ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5203 net2741 vssd1 vssd1 vccd1 vccd1 net5730 sky130_fd_sc_hd__dlygate4sd3_1
X_20587__320 clknet_1_0__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__inv_2
Xhold5214 net3190 vssd1 vssd1 vccd1 vccd1 net5741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5225 _01185_ vssd1 vssd1 vccd1 vccd1 net5752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22141_ clknet_leaf_40_i_clk _01628_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5236 rbzero.pov.spi_buffer\[70\] vssd1 vssd1 vccd1 vccd1 net5763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5247 net3446 vssd1 vssd1 vccd1 vccd1 net5774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4502 net699 vssd1 vssd1 vccd1 vccd1 net5029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4513 rbzero.spi_registers.texadd3\[1\] vssd1 vssd1 vccd1 vccd1 net5040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5258 _03073_ vssd1 vssd1 vccd1 vccd1 net5785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4524 net692 vssd1 vssd1 vccd1 vccd1 net5051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5269 net3499 vssd1 vssd1 vccd1 vccd1 net5796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4535 _00816_ vssd1 vssd1 vccd1 vccd1 net5062 sky130_fd_sc_hd__dlygate4sd3_1
X_22072_ net514 net1940 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold3801 _03676_ vssd1 vssd1 vccd1 vccd1 net4328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4546 net725 vssd1 vssd1 vccd1 vccd1 net5073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4557 rbzero.spi_registers.texadd2\[11\] vssd1 vssd1 vccd1 vccd1 net5084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3812 net3405 vssd1 vssd1 vccd1 vccd1 net4339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3823 net7876 vssd1 vssd1 vccd1 vccd1 net4350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4568 net724 vssd1 vssd1 vccd1 vccd1 net5095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21023_ clknet_leaf_63_i_clk net4276 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3834 net3423 vssd1 vssd1 vccd1 vccd1 net4361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4579 _00863_ vssd1 vssd1 vccd1 vccd1 net5106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3845 net8373 vssd1 vssd1 vccd1 vccd1 net4372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3856 net7868 vssd1 vssd1 vccd1 vccd1 net4383 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3867 _00775_ vssd1 vssd1 vccd1 vccd1 net4394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3878 net7904 vssd1 vssd1 vccd1 vccd1 net4405 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3889 rbzero.debug_overlay.facingY\[-1\] vssd1 vssd1 vccd1 vccd1 net4416 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21925_ net367 net2025 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21856_ net298 net657 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ net5726 _03877_ _03874_ _03973_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21787_ clknet_leaf_4_i_clk net1401 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ net4138 _04728_ net4393 _04657_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20738_ net896 net5376 vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11471_ _04659_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__or2b_1
XFILLER_0_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7150 net7743 vssd1 vssd1 vccd1 vccd1 net7677 sky130_fd_sc_hd__dlygate4sd3_1
X_13210_ _06306_ _06370_ _06378_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__o211a_1
Xhold7161 _02732_ vssd1 vssd1 vccd1 vccd1 net7688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7172 rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 net7699 sky130_fd_sc_hd__dlygate4sd3_1
X_14190_ _07314_ _07346_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7183 net4115 vssd1 vssd1 vccd1 vccd1 net7710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7194 rbzero.color_floor\[2\] vssd1 vssd1 vccd1 vccd1 net7721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6460 net2456 vssd1 vssd1 vccd1 vccd1 net6987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6471 rbzero.tex_r1\[36\] vssd1 vssd1 vccd1 vccd1 net6998 sky130_fd_sc_hd__dlygate4sd3_1
X_13141_ _06288_ _06278_ _06291_ _06293_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__a31o_1
Xhold6482 net2247 vssd1 vssd1 vccd1 vccd1 net7009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6493 rbzero.pov.ready_buffer\[15\] vssd1 vssd1 vccd1 vccd1 net7020 sky130_fd_sc_hd__dlygate4sd3_1
X_13072_ net5531 _06242_ _06241_ _06246_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a22o_1
Xhold5770 net1295 vssd1 vssd1 vccd1 vccd1 net6297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5781 rbzero.spi_registers.new_texadd\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net6308
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5792 net1363 vssd1 vssd1 vccd1 vccd1 net6319 sky130_fd_sc_hd__dlygate4sd3_1
X_16900_ _09615_ _09623_ _09621_ vssd1 vssd1 vccd1 vccd1 _09922_ sky130_fd_sc_hd__a21oi_1
X_12023_ _05206_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__or2_1
X_17880_ _10432_ _09114_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16831_ _09856_ net4500 net4649 vssd1 vssd1 vccd1 vccd1 _09857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19550_ net6960 net2205 _03388_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
X_16762_ _09794_ net4667 _09769_ vssd1 vssd1 vccd1 vccd1 _09795_ sky130_fd_sc_hd__mux2_1
X_13974_ net535 _07089_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__xnor2_4
X_18501_ _02658_ _02661_ _02659_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a21bo_1
X_15713_ _08806_ _08805_ _08807_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__nand3_1
XFILLER_0_38_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19481_ net1622 net6019 _03354_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__mux2_1
X_12925_ _06098_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__nor2_1
X_16693_ net822 _09743_ _09744_ net8021 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__a22o_1
X_18432_ _02593_ _02599_ _02587_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__o21ai_1
X_15644_ _08735_ _08737_ _08738_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__nand3_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12856_ net4043 vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__inv_2
XFILLER_0_180_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _04979_ vssd1 vssd1 vccd1 vccd1 _04997_
+ sky130_fd_sc_hd__mux2_1
X_18363_ net4501 net4733 _05155_ net3565 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _08180_ _08204_ _08205_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__xor2_1
X_17314_ _10314_ _10315_ _10332_ vssd1 vssd1 vccd1 vccd1 _10333_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_105_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _07688_ _07687_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__and2b_1
X_11738_ net86 vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__buf_4
X_18294_ net1860 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ _10136_ _10140_ _10262_ _10263_ vssd1 vssd1 vccd1 vccd1 _10264_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14457_ _07585_ _07597_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ net3014 _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13408_ _06462_ _06558_ _06578_ _06491_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__a211o_1
X_17176_ _09262_ _09025_ vssd1 vssd1 vccd1 vccd1 _10196_ sky130_fd_sc_hd__nor2_1
X_14388_ _07556_ _07558_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ _09129_ _09198_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13339_ _06505_ _06506_ _06509_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16058_ _09150_ _09151_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__nand2_1
Xhold3108 net5822 vssd1 vssd1 vccd1 vccd1 net3635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3119 _03331_ vssd1 vssd1 vccd1 vccd1 net3646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15009_ net3988 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__clkbuf_1
Xhold2407 net1102 vssd1 vssd1 vccd1 vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2418 _00658_ vssd1 vssd1 vccd1 vccd1 net2945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2429 net3144 vssd1 vssd1 vccd1 vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1706 _03359_ vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_19817_ net2311 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__clkbuf_1
Xhold1717 rbzero.tex_g1\[57\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 _01332_ vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _04296_ vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_205_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19679_ net6399 net3402 _03457_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21710_ clknet_leaf_109_i_clk net4628 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20619__349 clknet_1_0__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__inv_2
X_21641_ clknet_leaf_116_i_clk net3168 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21572_ net206 net2383 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_10 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 rbzero.wall_tracer.visualWallDist\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net6143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_54 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_98 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5000 _03133_ vssd1 vssd1 vccd1 vccd1 net5527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5011 net1804 vssd1 vssd1 vccd1 vccd1 net5538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5022 net2153 vssd1 vssd1 vccd1 vccd1 net5549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5033 net1276 vssd1 vssd1 vccd1 vccd1 net5560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5044 _03132_ vssd1 vssd1 vccd1 vccd1 net5571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5055 net8210 vssd1 vssd1 vccd1 vccd1 net5582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4310 net1032 vssd1 vssd1 vccd1 vccd1 net4837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5066 _04358_ vssd1 vssd1 vccd1 vccd1 net5593 sky130_fd_sc_hd__dlygate4sd3_1
X_22124_ clknet_leaf_54_i_clk net5450 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold4321 net892 vssd1 vssd1 vccd1 vccd1 net4848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4332 _00636_ vssd1 vssd1 vccd1 vccd1 net4859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5077 rbzero.wall_tracer.mapY\[6\] vssd1 vssd1 vccd1 vccd1 net5604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4343 _00608_ vssd1 vssd1 vccd1 vccd1 net4870 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_84_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold5088 _00773_ vssd1 vssd1 vccd1 vccd1 net5615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5099 net2835 vssd1 vssd1 vccd1 vccd1 net5626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4354 net943 vssd1 vssd1 vccd1 vccd1 net4881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3620 net4121 vssd1 vssd1 vccd1 vccd1 net4147 sky130_fd_sc_hd__buf_4
X_22055_ net497 net2372 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold4376 _01191_ vssd1 vssd1 vccd1 vccd1 net4903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3631 _00457_ vssd1 vssd1 vccd1 vccd1 net4158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4387 _10027_ vssd1 vssd1 vccd1 vccd1 net4914 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3642 _05112_ vssd1 vssd1 vccd1 vccd1 net4169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3653 rbzero.side_hot vssd1 vssd1 vccd1 vccd1 net4180 sky130_fd_sc_hd__buf_2
Xhold4398 rbzero.wall_tracer.trackDistY\[-8\] vssd1 vssd1 vccd1 vccd1 net4925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3664 net7861 vssd1 vssd1 vccd1 vccd1 net4191 sky130_fd_sc_hd__dlygate4sd3_1
X_21006_ clknet_leaf_81_i_clk _00493_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20364__119 clknet_1_0__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__inv_2
Xhold3675 net7886 vssd1 vssd1 vccd1 vccd1 net4202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2930 net8213 vssd1 vssd1 vccd1 vccd1 net3457 sky130_fd_sc_hd__buf_2
Xhold3686 net7898 vssd1 vssd1 vccd1 vccd1 net4213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2941 net8057 vssd1 vssd1 vccd1 vccd1 net3468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3697 net7910 vssd1 vssd1 vccd1 vccd1 net4224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2952 _03100_ vssd1 vssd1 vccd1 vccd1 net3479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2963 net4619 vssd1 vssd1 vccd1 vccd1 net3490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2974 net8358 vssd1 vssd1 vccd1 vccd1 net3501 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_99_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2985 _01224_ vssd1 vssd1 vccd1 vccd1 net3512 sky130_fd_sc_hd__dlygate4sd3_1
X_10971_ net1716 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _05850_ _05851_ net4147 _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a31o_1
X_21908_ net350 net2693 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap78 _06722_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13690_ _06854_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_22_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xmax_cap89 net91 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_2
XFILLER_0_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ net49 _05818_ _05819_ _05814_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a211o_1
X_21839_ net281 net2992 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15360_ rbzero.wall_tracer.visualWallDist\[-11\] _08117_ vssd1 vssd1 vccd1 vccd1
+ _08455_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ _05749_ net4068 net20 _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ _07461_ _07481_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ net4127 net2038 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nand2_1
X_15291_ _08374_ _08375_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_37_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17030_ _10049_ _10050_ vssd1 vssd1 vccd1 vccd1 _10051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ _06755_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11454_ _04630_ _04631_ _04638_ _04645_ _04495_ _04545_ vssd1 vssd1 vccd1 vccd1 _04646_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14173_ _07284_ _07305_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__nor2_1
X_11385_ _04569_ _04575_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6290 rbzero.tex_g1\[61\] vssd1 vssd1 vccd1 vccd1 net6817 sky130_fd_sc_hd__dlygate4sd3_1
X_13124_ _06279_ _06283_ _06284_ _06293_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a221o_1
X_18981_ net3099 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ net8008 _09410_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__nor2_1
X_13055_ _06230_ _06200_ _06197_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__nand3b_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ net4177 _04462_ _04684_ _04682_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__o22a_1
XFILLER_0_206_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17863_ _10163_ net4913 _02099_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19602_ net4815 net4834 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16814_ net4508 net4383 vssd1 vssd1 vccd1 vccd1 _09841_ sky130_fd_sc_hd__nor2_1
X_17794_ _02031_ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ net5472 _09103_ _09778_ vssd1 vssd1 vccd1 vccd1 _09780_ sky130_fd_sc_hd__a21bo_1
X_19533_ net3838 net5570 net3086 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__mux2_1
X_13957_ _07117_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19464_ _04458_ _02954_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or3_4
X_12908_ net4019 vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__inv_2
X_16676_ net4321 _09741_ _09742_ net672 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ _07056_ _07049_ _07054_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15627_ _08715_ _08721_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__and2_1
X_18415_ net4725 _02586_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__and2_1
X_19395_ net3217 _03123_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and2_1
X_12839_ _05967_ _06014_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__xnor2_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _02529_ _02532_ _04489_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a21oi_1
X_15558_ _08650_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__nand2_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14509_ _07675_ _07678_ _07679_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__a21bo_1
Xhold7919 rbzero.wall_tracer.stepDistX\[-3\] vssd1 vssd1 vccd1 vccd1 net8446 sky130_fd_sc_hd__dlygate4sd3_1
X_18277_ net6299 net4016 _02477_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
X_15489_ _08570_ _08577_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17228_ _10023_ _10122_ _10247_ vssd1 vssd1 vccd1 vccd1 _10248_ sky130_fd_sc_hd__a21oi_2
Xinput30 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03866_ clknet_0__03866_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03866_
+ sky130_fd_sc_hd__clkbuf_16
Xinput41 i_mode[1] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_8
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput52 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_8
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold803 _00982_ vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ _10079_ _10148_ _10178_ vssd1 vssd1 vccd1 vccd1 _10179_ sky130_fd_sc_hd__a21o_1
Xhold814 _03815_ vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 net6441 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold836 net6318 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 net6366 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _01537_ vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
X_20170_ net7544 _03707_ net4487 _03732_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold869 net4029 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__buf_4
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2204 net7233 vssd1 vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2215 net5731 vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2226 net5725 vssd1 vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 net7553 vssd1 vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1503 _04231_ vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2248 _04065_ vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 net7286 vssd1 vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1514 net5599 vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 net6755 vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1536 net6893 vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _01030_ vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1558 net6773 vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1569 _01503_ vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21624_ clknet_leaf_101_i_clk net3175 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21555_ net189 net1826 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21486_ clknet_leaf_48_i_clk net1670 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11170_ net2805 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4140 net3382 vssd1 vssd1 vccd1 vccd1 net4667 sky130_fd_sc_hd__clkbuf_2
X_22107_ net145 net2028 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4162 net747 vssd1 vssd1 vccd1 vccd1 net4689 sky130_fd_sc_hd__dlygate4sd3_1
X_20299_ net1442 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
Xhold4173 _01225_ vssd1 vssd1 vccd1 vccd1 net4700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4184 _01239_ vssd1 vssd1 vccd1 vccd1 net4711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4195 net8005 vssd1 vssd1 vccd1 vccd1 net4722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3450 _01624_ vssd1 vssd1 vccd1 vccd1 net3977 sky130_fd_sc_hd__dlygate4sd3_1
X_22038_ net480 net2329 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
Xhold3461 _08106_ vssd1 vssd1 vccd1 vccd1 net3988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3472 _06109_ vssd1 vssd1 vccd1 vccd1 net3999 sky130_fd_sc_hd__clkbuf_4
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3483 _08107_ vssd1 vssd1 vccd1 vccd1 net4010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3494 _03658_ vssd1 vssd1 vccd1 vccd1 net4021 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2760 _03586_ vssd1 vssd1 vccd1 vccd1 net3287 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2771 net1646 vssd1 vssd1 vccd1 vccd1 net3298 sky130_fd_sc_hd__dlygate4sd3_1
X_14860_ _07934_ _08012_ _08013_ _08014_ _06543_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__o311a_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2782 net5926 vssd1 vssd1 vccd1 vccd1 net3309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2793 net1151 vssd1 vssd1 vccd1 vccd1 net3320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ net578 net534 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__xnor2_2
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _07913_ _07914_ _07934_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__a21oi_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _09481_ _09619_ vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ net546 _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__xnor2_1
X_10954_ net1740 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _09548_ _09417_ _06124_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ _06729_ _06721_ net540 _06719_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__o2bb2a_1
X_10885_ net7291 net6884 _04253_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18200_ net3669 net4459 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__nand2_1
X_15412_ _08483_ _08487_ _08506_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__o21ai_2
X_12624_ _05802_ net4156 vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__nor2_1
X_19180_ net6367 _03170_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__or2_1
X_16392_ _09479_ _09480_ _09482_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18131_ _02358_ _02359_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__or2b_1
XFILLER_0_171_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15343_ _08436_ _08422_ _08360_ _08437_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__a31o_1
X_12555_ net13 _05732_ _05735_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18062_ _01794_ _01693_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ net4110 net4188 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15274_ _07968_ _07975_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12486_ net44 _05644_ _05641_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a21bo_1
X_17013_ _10032_ _10033_ vssd1 vssd1 vccd1 vccd1 _10034_ sky130_fd_sc_hd__xnor2_1
X_14225_ _07284_ _07310_ _07281_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11437_ _04624_ _04626_ _04627_ _04628_ _04503_ _04496_ vssd1 vssd1 vccd1 vccd1 _04629_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ _07326_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ rbzero.spi_registers.texadd3\[18\] rbzero.spi_registers.texadd1\[18\] rbzero.spi_registers.texadd0\[18\]
+ rbzero.spi_registers.texadd2\[18\] _04554_ _04555_ vssd1 vssd1 vccd1 vccd1 _04560_
+ sky130_fd_sc_hd__mux4_2
X_13107_ _06270_ _06276_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _07212_ _07213_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__or2_1
X_18964_ net3324 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__clkbuf_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _01949_ _01951_ _02049_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__o31ai_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _06212_ net3669 _06213_ net3811 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a22o_1
X_18895_ _02992_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _01794_ _10220_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nor2_1
X_17777_ _10062_ _09410_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__nor2_1
X_14989_ _08092_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19516_ net1641 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ _09750_ _09764_ vssd1 vssd1 vccd1 vccd1 _09766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19447_ net3978 _03123_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ _04478_ _09734_ vssd1 vssd1 vccd1 vccd1 _09738_ sky130_fd_sc_hd__nor2_4
XFILLER_0_53_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19378_ net6496 _03284_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7705 _03893_ vssd1 vssd1 vccd1 vccd1 net8232 sky130_fd_sc_hd__dlygate4sd3_1
X_18329_ net4501 net4852 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__nand2_1
Xhold7716 _02910_ vssd1 vssd1 vccd1 vccd1 net8243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7727 rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 net8254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7738 net8009 vssd1 vssd1 vccd1 vccd1 net8265 sky130_fd_sc_hd__clkbuf_2
Xhold7749 rbzero.spi_registers.new_texadd\[0\]\[22\] vssd1 vssd1 vccd1 vccd1 net8276
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21340_ clknet_leaf_4_i_clk net5059 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21271_ clknet_leaf_27_i_clk net4317 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03849_ clknet_0__03849_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03849_
+ sky130_fd_sc_hd__clkbuf_16
Xhold600 net6202 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold611 net7855 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_1
Xhold622 net6216 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _01329_ vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
X_20222_ net3621 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
Xhold644 net4590 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold655 net6246 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold666 _01451_ vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold677 _03151_ vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
X_20153_ _03728_ net7640 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__or2_1
Xhold688 _03823_ vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 net6272 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2001 net7108 vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2012 net7362 vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2023 _01595_ vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
X_20084_ net3445 _03660_ net5772 _03679_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__o211a_1
Xhold2034 _04062_ vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 net7243 vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 net6636 vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _01022_ vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2056 _01517_ vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1322 net6670 vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2067 _01474_ vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2078 _04278_ vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1333 _02495_ vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2089 net7189 vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1344 _01159_ vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1355 _03398_ vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 _01346_ vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1377 net6728 vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1388 net7142 vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 net6833 vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ clknet_leaf_30_i_clk net3860 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10670_ net6703 net6084 _04138_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21607_ clknet_leaf_131_i_clk net3028 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _05249_ vssd1 vssd1 vccd1 vccd1 _05526_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21538_ net172 net2166 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12271_ _05189_ _05456_ _05457_ _04707_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21469_ clknet_leaf_21_i_clk net1394 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14010_ _07118_ _07126_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__o21a_1
X_11222_ net7125 net2917 _04434_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__mux2_1
X_11153_ net7204 net2539 _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15961_ _09054_ _09055_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__and2b_1
X_11084_ net3243 net6846 _04364_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
Xhold3280 net7668 vssd1 vssd1 vccd1 vccd1 net3807 sky130_fd_sc_hd__buf_2
X_17700_ _01857_ _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__xnor2_1
X_14912_ net4665 _08050_ _08036_ net4567 net4551 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__o221a_1
Xhold3291 _00729_ vssd1 vssd1 vccd1 vccd1 net3818 sky130_fd_sc_hd__dlygate4sd3_1
X_15892_ _08754_ _08812_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__nor2_2
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18680_ _02559_ net4765 net8094 net3915 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2590 net7503 vssd1 vssd1 vccd1 vccd1 net3117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _01869_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__xor2_2
X_14843_ _07959_ _07972_ _07913_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__mux2_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03869_ clknet_0__03869_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03869_
+ sky130_fd_sc_hd__clkbuf_16
X_17562_ _01688_ _01782_ _01801_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__nand3_1
X_14774_ _07939_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _04664_ _05058_ net4171 net4140 vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__a211o_1
X_16513_ _09133_ net4909 vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__and2_1
X_19301_ net5296 _03236_ _03247_ _03246_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__o211a_1
X_13725_ _06893_ _06895_ _06891_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10937_ net7232 net6723 _04287_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17493_ _01732_ _01733_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16444_ _08916_ _09403_ _09411_ _08948_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__o22ai_1
X_19232_ net6341 _03203_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__or2_1
X_13656_ _06823_ _06825_ _06826_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10868_ net7131 net2685 _04171_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ net6041 _05745_ _05783_ net54 vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
X_19163_ net5392 _03144_ _03165_ _03160_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__o211a_1
X_16375_ _09389_ _09371_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__or2b_1
XFILLER_0_183_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13587_ _06701_ _06705_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_171_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _04193_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__clkbuf_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18114_ net3731 _02336_ _02337_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ net3453 vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__buf_4
XFILLER_0_186_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19094_ _03122_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__buf_6
X_12538_ clknet_1_1__leaf__05645_ _05712_ _05697_ net6100 _05718_ vssd1 vssd1 vccd1
+ vccd1 _05719_ sky130_fd_sc_hd__o221a_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18045_ _01760_ _09114_ _02206_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15257_ _08285_ _08336_ _08351_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__a21oi_1
X_12469_ net52 _05646_ _05642_ net53 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4909 net1087 vssd1 vssd1 vccd1 vccd1 net5436 sky130_fd_sc_hd__dlygate4sd3_1
X_14208_ _07372_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__o21ba_1
X_15188_ _08273_ _08281_ _08282_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ _07307_ _07309_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__xnor2_4
X_20581__315 clknet_1_1__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__inv_2
X_19996_ _03122_ _03483_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18947_ net2089 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18878_ net3112 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
X_17829_ _01818_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20840_ _03320_ clknet_1_0__leaf__05794_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__and2_2
X_20771_ net864 net5488 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7502 net4584 vssd1 vssd1 vccd1 vccd1 net8029 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7524 net4811 vssd1 vssd1 vccd1 vccd1 net8051 sky130_fd_sc_hd__clkbuf_4
Xhold7535 _02885_ vssd1 vssd1 vccd1 vccd1 net8062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6801 net2438 vssd1 vssd1 vccd1 vccd1 net7328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6812 rbzero.tex_g1\[17\] vssd1 vssd1 vccd1 vccd1 net7339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7557 _02640_ vssd1 vssd1 vccd1 vccd1 net8084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6823 rbzero.tex_g1\[3\] vssd1 vssd1 vccd1 vccd1 net7350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7568 _00630_ vssd1 vssd1 vccd1 vccd1 net8095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6834 net2482 vssd1 vssd1 vccd1 vccd1 net7361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7579 _01648_ vssd1 vssd1 vccd1 vccd1 net8106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6845 rbzero.tex_g1\[29\] vssd1 vssd1 vccd1 vccd1 net7372 sky130_fd_sc_hd__dlygate4sd3_1
X_20333__91 clknet_1_0__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__inv_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21323_ clknet_leaf_12_i_clk net5354 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6856 net2557 vssd1 vssd1 vccd1 vccd1 net7383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6867 rbzero.spi_registers.new_mapd\[3\] vssd1 vssd1 vccd1 vccd1 net7394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6878 net2987 vssd1 vssd1 vccd1 vccd1 net7405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6889 rbzero.tex_b0\[43\] vssd1 vssd1 vccd1 vccd1 net7416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21254_ clknet_leaf_2_i_clk net3480 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold430 net7302 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 net7922 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 net5353 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold463 net5413 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20205_ net2364 _03743_ net4555 _03732_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__o211a_1
X_21185_ clknet_leaf_102_i_clk net2487 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold474 net5345 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold485 net5389 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 net7888 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
X_20136_ _03689_ net7663 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or2_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ _03661_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__or2_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _00958_ vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 net6541 vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 _00585_ vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _01112_ vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 _03379_ vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 net6537 vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _01036_ vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ net1822 net4271 _04851_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or4_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _04923_ vssd1 vssd1 vccd1 vccd1 _04961_
+ sky130_fd_sc_hd__mux2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ clknet_leaf_88_i_clk _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _06546_ _06675_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__a21o_1
X_10722_ net6361 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _07284_ _07390_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__nor2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _06392_ net82 _06525_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__or3_1
X_10653_ net2095 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16160_ _09251_ _09252_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _06540_ _06541_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__o21ai_4
X_10584_ net5560 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__clkbuf_1
X_15111_ _08204_ _08205_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__nand2_1
X_12323_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _05237_ vssd1 vssd1 vccd1 vccd1 _05509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16091_ _09168_ _09184_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20530__269 clknet_1_1__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__inv_2
X_15042_ _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__buf_4
X_12254_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _04933_ vssd1 vssd1 vccd1 vccd1 _05441_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11205_ net7459 net7202 _04423_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19850_ net6247 net3077 _03528_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__mux2_1
X_12185_ _05033_ _05035_ _05371_ _05372_ net3781 vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18801_ net5957 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
X_11136_ net6026 net2279 _04390_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__mux2_1
X_16993_ net4589 net4483 vssd1 vssd1 vccd1 vccd1 _10014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18732_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _02856_
+ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__o21a_1
X_11067_ net5592 net5649 _04353_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__mux2_1
X_15944_ _09032_ _09038_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15875_ _08967_ _08968_ _08969_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__or3_1
X_18663_ rbzero.wall_tracer.rayAddendY\[0\] _02818_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02819_ sky130_fd_sc_hd__mux2_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20424__174 clknet_1_0__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__inv_2
X_17614_ _01756_ _01757_ _01754_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14826_ _07821_ _07830_ _07971_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__a21oi_1
X_18594_ net4598 net681 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__or2_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _01783_ _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__xnor2_1
X_14757_ net7845 _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ _05155_ _05113_ _05156_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a211o_1
X_13708_ _06871_ _06866_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__xnor2_2
X_17476_ _10273_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14688_ net7812 vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19215_ net1649 _03169_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__or2_1
X_16427_ _09507_ _09517_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__xnor2_1
X_13639_ _06735_ _06738_ _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ _09335_ _09449_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19146_ net4366 _03145_ net958 _03149_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6108 net1892 vssd1 vssd1 vccd1 vccd1 net6635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6119 rbzero.spi_registers.new_texadd\[0\]\[11\] vssd1 vssd1 vccd1 vccd1 net6646
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15309_ _07968_ _07975_ _07981_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__o21a_4
X_16289_ _08308_ _08418_ _09380_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19077_ net2047 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__clkbuf_1
Xhold5407 _02718_ vssd1 vssd1 vccd1 vccd1 net5934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5418 gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 net5945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5429 _02946_ vssd1 vssd1 vccd1 vccd1 net5956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ _02260_ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__xnor2_1
Xhold4706 _00798_ vssd1 vssd1 vccd1 vccd1 net5233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4717 net806 vssd1 vssd1 vccd1 vccd1 net5244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4728 rbzero.spi_registers.texadd0\[7\] vssd1 vssd1 vccd1 vccd1 net5255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4739 net861 vssd1 vssd1 vccd1 vccd1 net5266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19979_ net7506 net3199 _08092_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21941_ net383 net2653 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21872_ net314 net1271 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20399__151 clknet_1_1__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__inv_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _03985_ _03986_ net5609 net63 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20754_ _03924_ _03925_ _03926_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_4__f_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7310 net7821 vssd1 vssd1 vccd1 vccd1 net7837 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7321 net4427 vssd1 vssd1 vccd1 vccd1 net7848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7343 net4380 vssd1 vssd1 vccd1 vccd1 net7870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7354 rbzero.traced_texVinit\[10\] vssd1 vssd1 vccd1 vccd1 net7881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6620 net2841 vssd1 vssd1 vccd1 vccd1 net7147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7365 net1008 vssd1 vssd1 vccd1 vccd1 net7892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6631 _04329_ vssd1 vssd1 vccd1 vccd1 net7158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7376 net4404 vssd1 vssd1 vccd1 vccd1 net7903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6642 net2283 vssd1 vssd1 vccd1 vccd1 net7169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7387 net757 vssd1 vssd1 vccd1 vccd1 net7914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6653 net2569 vssd1 vssd1 vccd1 vccd1 net7180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7398 _00502_ vssd1 vssd1 vccd1 vccd1 net7925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6664 rbzero.tex_r1\[24\] vssd1 vssd1 vccd1 vccd1 net7191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6675 net2607 vssd1 vssd1 vccd1 vccd1 net7202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5930 _04211_ vssd1 vssd1 vccd1 vccd1 net6457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21306_ clknet_leaf_10_i_clk net5214 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5941 net1451 vssd1 vssd1 vccd1 vccd1 net6468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6686 _04315_ vssd1 vssd1 vccd1 vccd1 net7213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5952 _04228_ vssd1 vssd1 vccd1 vccd1 net6479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6697 net2390 vssd1 vssd1 vccd1 vccd1 net7224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5963 net1521 vssd1 vssd1 vccd1 vccd1 net6490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5974 _04307_ vssd1 vssd1 vccd1 vccd1 net6501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5985 net1222 vssd1 vssd1 vccd1 vccd1 net6512 sky130_fd_sc_hd__dlygate4sd3_1
X_21237_ clknet_leaf_13_i_clk net4078 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold260 net5136 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5996 rbzero.tex_b1\[35\] vssd1 vssd1 vccd1 vccd1 net6523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 net5110 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net5174 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 net5223 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
X_20683__4 clknet_1_0__leaf__03506_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
X_21168_ clknet_leaf_98_i_clk net3021 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_20119_ _03706_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__clkbuf_4
X_13990_ _07104_ _06832_ _07159_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__o21a_1
X_21099_ clknet_leaf_9_i_clk net1382 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12941_ net5922 net3975 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__and2b_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _08650_ _08652_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__or2_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ net3807 vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__inv_2
XANTENNA_100 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _07558_ _07781_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__xnor2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11823_ net5968 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__clkbuf_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15591_ _08684_ _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__xor2_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _08948_ _08916_ _09970_ vssd1 vssd1 vccd1 vccd1 _10349_ sky130_fd_sc_hd__a21oi_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _07072_ _07194_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__or2_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _04924_ vssd1 vssd1 vccd1 vccd1 _04944_
+ sky130_fd_sc_hd__mux2_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _08226_ _09472_ vssd1 vssd1 vccd1 vccd1 _10280_ sky130_fd_sc_hd__nor2_1
X_10705_ net6965 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__clkbuf_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14473_ _07631_ _07642_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11685_ _04856_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16212_ _09300_ _09304_ _09183_ _09184_ _09168_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__a32o_1
XFILLER_0_148_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19000_ net3237 net5791 _02992_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ _06550_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__or3_1
X_10636_ net6671 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__clkbuf_1
X_17192_ _08880_ _10211_ _09411_ _10096_ vssd1 vssd1 vccd1 vccd1 _10212_ sky130_fd_sc_hd__or4_2
XFILLER_0_64_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _09134_ _09229_ _09235_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ _06489_ _06525_ net82 vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10567_ net2371 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _04912_ vssd1 vssd1 vccd1 vccd1 _05492_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16074_ _09163_ _09167_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__xor2_2
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13286_ _06346_ _06350_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10498_ net7065 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__clkbuf_1
X_19902_ net2312 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__clkbuf_4
X_15025_ rbzero.wall_tracer.rayAddendY\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] net4181
+ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__mux2_1
X_12237_ rbzero.tex_g1\[41\] rbzero.tex_g1\[40\] _04968_ vssd1 vssd1 vccd1 vccd1 _05424_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19833_ net7310 net3026 _03517_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
X_12168_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _04916_ vssd1 vssd1 vccd1 vccd1 _05356_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11119_ net5684 net7342 _04375_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16976_ _09633_ _09700_ _09698_ vssd1 vssd1 vccd1 vccd1 _09998_ sky130_fd_sc_hd__a21o_1
X_12099_ net1822 _04991_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__nor2_1
X_18715_ _02866_ rbzero.wall_tracer.rayAddendY\[3\] _02862_ vssd1 vssd1 vccd1 vccd1
+ _02867_ sky130_fd_sc_hd__a21oi_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _09020_ _09021_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__xnor2_2
Xinput6 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19695_ net6424 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18646_ net8026 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__inv_2
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _08939_ _08952_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__xor2_1
X_19784__63 clknet_1_1__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
X_14809_ net7813 _07899_ _07900_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__and3_1
X_18577_ _09760_ _02740_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15789_ _08878_ _08883_ _08876_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17528_ _01761_ _10437_ _01767_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17459_ _10352_ _10353_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19129_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5204 _04084_ vssd1 vssd1 vccd1 vccd1 net5731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5215 rbzero.pov.ready_buffer\[49\] vssd1 vssd1 vccd1 vccd1 net5742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5226 net3373 vssd1 vssd1 vccd1 vccd1 net5753 sky130_fd_sc_hd__dlygate4sd3_1
X_22140_ clknet_leaf_24_i_clk _01627_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold5237 net1979 vssd1 vssd1 vccd1 vccd1 net5764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4503 _00814_ vssd1 vssd1 vccd1 vccd1 net5030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5259 net1614 vssd1 vssd1 vccd1 vccd1 net5786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4514 net709 vssd1 vssd1 vccd1 vccd1 net5041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4525 rbzero.spi_registers.texadd0\[1\] vssd1 vssd1 vccd1 vccd1 net5052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4536 net827 vssd1 vssd1 vccd1 vccd1 net5063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22071_ net513 net2721 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3802 _01188_ vssd1 vssd1 vccd1 vccd1 net4329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4547 _00839_ vssd1 vssd1 vccd1 vccd1 net5074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4558 net695 vssd1 vssd1 vccd1 vccd1 net5085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3813 net8312 vssd1 vssd1 vccd1 vccd1 net4340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3824 net7878 vssd1 vssd1 vccd1 vccd1 net4351 sky130_fd_sc_hd__buf_1
XFILLER_0_125_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4569 rbzero.spi_registers.texadd1\[4\] vssd1 vssd1 vccd1 vccd1 net5096 sky130_fd_sc_hd__dlygate4sd3_1
X_21022_ clknet_leaf_63_i_clk net4258 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3835 net5742 vssd1 vssd1 vccd1 vccd1 net4362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3846 net3430 vssd1 vssd1 vccd1 vccd1 net4373 sky130_fd_sc_hd__buf_1
Xhold3857 net8168 vssd1 vssd1 vccd1 vccd1 net4384 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3868 net1832 vssd1 vssd1 vccd1 vccd1 net4395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3879 net8318 vssd1 vssd1 vccd1 vccd1 net4406 sky130_fd_sc_hd__dlygate4sd3_1
X_21924_ net366 net2401 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ net297 net2699 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20806_ _03969_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21786_ clknet_leaf_1_i_clk net2222 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20737_ _03909_ _03910_ _03911_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ net4110 net4023 net4102 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__nor3_2
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7140 net3782 vssd1 vssd1 vccd1 vccd1 net7667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7151 net3954 vssd1 vssd1 vccd1 vccd1 net7678 sky130_fd_sc_hd__buf_2
XFILLER_0_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7162 rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 net7689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7173 rbzero.debug_overlay.playerX\[3\] vssd1 vssd1 vccd1 vccd1 net7700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7184 rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 net7711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6450 net2230 vssd1 vssd1 vccd1 vccd1 net6977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7195 net3547 vssd1 vssd1 vccd1 vccd1 net7722 sky130_fd_sc_hd__dlygate4sd3_1
X_13140_ _06282_ _06283_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6461 rbzero.tex_r0\[20\] vssd1 vssd1 vccd1 vccd1 net6988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6472 net2560 vssd1 vssd1 vccd1 vccd1 net6999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6483 _04118_ vssd1 vssd1 vccd1 vccd1 net7010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6494 net2161 vssd1 vssd1 vccd1 vccd1 net7021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5760 net1292 vssd1 vssd1 vccd1 vccd1 net6287 sky130_fd_sc_hd__dlygate4sd3_1
X_13071_ _06243_ _06245_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5771 rbzero.spi_registers.new_texadd\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net6298
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5782 net1322 vssd1 vssd1 vccd1 vccd1 net6309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5793 rbzero.spi_registers.new_texadd\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 net6320
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12022_ rbzero.tex_r1\[3\] rbzero.tex_r1\[2\] _04979_ vssd1 vssd1 vccd1 vccd1 _05211_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16830_ _06058_ _09854_ _09855_ vssd1 vssd1 vccd1 vccd1 _09856_ sky130_fd_sc_hd__o21ai_1
X_16761_ _09788_ net3805 _09790_ _09793_ vssd1 vssd1 vccd1 vccd1 _09794_ sky130_fd_sc_hd__a31o_1
X_13973_ net3498 _07093_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18500_ _02675_ _02676_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__nand2_1
X_15712_ _08749_ _08764_ _08804_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__a21o_1
X_12924_ net4366 net4642 _06048_ net4357 _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16692_ net834 _09743_ _09744_ net8018 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__a22o_1
X_19480_ net1879 _02472_ _04458_ _03344_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__or4_4
X_18431_ _02610_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15643_ _08729_ _08731_ _08734_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__a21o_1
X_12855_ _06030_ _06028_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__xnor2_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _04977_ _04993_ _04995_ _04829_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o211a_1
X_15574_ net3637 _08162_ net7836 _08185_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18362_ net5823 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__clkbuf_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__or2_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _10330_ _10331_ vssd1 vssd1 vccd1 vccd1 _10332_ sky130_fd_sc_hd__nand2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _07656_ net76 vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__xor2_2
X_11737_ _04910_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__or2_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ net6558 net3745 _02493_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20536__275 clknet_1_0__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__inv_2
X_17244_ net4610 net4405 vssd1 vssd1 vccd1 vccd1 _10263_ sky130_fd_sc_hd__nor2_1
X_14456_ _07624_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__nor2_1
X_11668_ net3151 net3488 _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ net561 net560 _06453_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ net2677 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__clkbuf_1
X_17175_ _10193_ _10194_ vssd1 vssd1 vccd1 vccd1 _10195_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14387_ _07506_ _07557_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__nor2_1
X_11599_ net2474 _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16126_ _09195_ _09197_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__or2_1
X_13338_ _06467_ net574 _06507_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16057_ _09131_ _09132_ _09149_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__nand3_1
XFILLER_0_110_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _06354_ _06319_ _06404_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_122_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3109 net5824 vssd1 vssd1 vccd1 vccd1 net3636 sky130_fd_sc_hd__dlygate4sd3_1
X_15008_ _08038_ net3987 vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__and2_1
Xhold2408 _03559_ vssd1 vssd1 vccd1 vccd1 net2935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2419 rbzero.tex_r0\[63\] vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
X_19816_ net2310 net7273 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__nand2_1
Xhold1707 _00915_ vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1718 net6911 vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 net6843 vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16959_ _09968_ _09979_ _09980_ vssd1 vssd1 vccd1 vccd1 _09981_ sky130_fd_sc_hd__nand3_1
XFILLER_0_155_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19678_ net1801 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18629_ rbzero.wall_tracer.rayAddendY\[-3\] _02787_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21640_ clknet_leaf_127_i_clk net3216 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21571_ net205 net2213 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_22 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 net6714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_55 _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_66 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_77 net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 net2094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_99 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5001 _00761_ vssd1 vssd1 vccd1 vccd1 net5528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5012 rbzero.spi_registers.new_other\[1\] vssd1 vssd1 vccd1 vccd1 net5539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5023 rbzero.tex_r1\[1\] vssd1 vssd1 vccd1 vccd1 net5550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5034 rbzero.spi_registers.new_vshift\[2\] vssd1 vssd1 vccd1 vccd1 net5561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4300 net1942 vssd1 vssd1 vccd1 vccd1 net4827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5045 _00760_ vssd1 vssd1 vccd1 vccd1 net5572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5056 net1617 vssd1 vssd1 vccd1 vccd1 net5583 sky130_fd_sc_hd__dlygate4sd3_1
X_22123_ clknet_leaf_54_i_clk net4982 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
Xhold4311 net3455 vssd1 vssd1 vccd1 vccd1 net4838 sky130_fd_sc_hd__clkbuf_2
Xhold5067 net1989 vssd1 vssd1 vccd1 vccd1 net5594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4322 _01654_ vssd1 vssd1 vccd1 vccd1 net4849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5078 net2277 vssd1 vssd1 vccd1 vccd1 net5605 sky130_fd_sc_hd__buf_1
Xhold4333 net3763 vssd1 vssd1 vccd1 vccd1 net4860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4344 net3616 vssd1 vssd1 vccd1 vccd1 net4871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5089 net2588 vssd1 vssd1 vccd1 vccd1 net5616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4355 rbzero.wall_tracer.rayAddendX\[-5\] vssd1 vssd1 vccd1 vccd1 net4882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3610 net7738 vssd1 vssd1 vccd1 vccd1 net4137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3621 _05052_ vssd1 vssd1 vccd1 vccd1 net4148 sky130_fd_sc_hd__dlygate4sd3_1
X_22054_ net496 net2526 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold4366 net8364 vssd1 vssd1 vccd1 vccd1 net4893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4377 net3327 vssd1 vssd1 vccd1 vccd1 net4904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3632 gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 net4159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3643 _05119_ vssd1 vssd1 vccd1 vccd1 net4170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4388 rbzero.wall_tracer.trackDistY\[-5\] vssd1 vssd1 vccd1 vccd1 net4915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4399 net3786 vssd1 vssd1 vccd1 vccd1 net4926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3654 _04510_ vssd1 vssd1 vccd1 vccd1 net4181 sky130_fd_sc_hd__buf_2
Xhold3665 net7863 vssd1 vssd1 vccd1 vccd1 net4192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2920 net7574 vssd1 vssd1 vccd1 vccd1 net3447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21005_ clknet_leaf_81_i_clk _00492_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2931 net5852 vssd1 vssd1 vccd1 vccd1 net3458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3676 net7881 vssd1 vssd1 vccd1 vccd1 net4203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3687 net7893 vssd1 vssd1 vccd1 vccd1 net4214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2942 rbzero.debug_overlay.playerY\[5\] vssd1 vssd1 vccd1 vccd1 net3469 sky130_fd_sc_hd__buf_2
Xhold3698 rbzero.wall_tracer.visualWallDist\[7\] vssd1 vssd1 vccd1 vccd1 net4225 sky130_fd_sc_hd__buf_1
Xhold2953 _00741_ vssd1 vssd1 vccd1 vccd1 net3480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2964 net8324 vssd1 vssd1 vccd1 vccd1 net3491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2975 net1585 vssd1 vssd1 vccd1 vccd1 net3502 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2997 net5804 vssd1 vssd1 vccd1 vccd1 net3524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19748__30 clknet_1_1__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
X_10970_ net6641 net6500 _04298_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21907_ net349 net2054 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap79 _06643_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_6
XFILLER_0_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ net50 _05797_ _05802_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__and3_1
X_19763__44 clknet_1_1__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
X_21838_ net280 net2624 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ net19 vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__inv_2
X_21769_ clknet_leaf_11_i_clk net1370 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _07479_ _07480_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__nor2_2
X_11522_ net4126 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__buf_1
X_15290_ _08200_ _08384_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _07401_ _07407_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__xor2_4
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _04502_ _04639_ _04641_ _04642_ _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__o32a_1
XFILLER_0_190_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14172_ _06725_ _07342_ _07309_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11384_ _04021_ _04569_ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__and3_1
Xhold6280 rbzero.tex_g1\[20\] vssd1 vssd1 vccd1 vccd1 net6807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and2_1
Xhold6291 net2226 vssd1 vssd1 vccd1 vccd1 net6818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18980_ net7455 net5745 _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5590 rbzero.tex_b1\[46\] vssd1 vssd1 vccd1 vccd1 net6117 sky130_fd_sc_hd__dlygate4sd3_1
X_17931_ _02166_ _02167_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__xnor2_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _06220_ _06226_ _06229_ _06215_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__o2bb2a_1
X_12005_ _04657_ _04464_ _04600_ net4095 _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17862_ _10163_ net4913 _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19601_ net1030 _03139_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__nand2_1
X_16813_ net4632 _09833_ _09834_ vssd1 vssd1 vccd1 vccd1 _09840_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17793_ _02014_ _02015_ _02030_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19532_ net7526 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
X_16744_ net5722 _09103_ vssd1 vssd1 vccd1 vccd1 _09779_ sky130_fd_sc_hd__xnor2_1
X_13956_ _07118_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__xnor2_1
X_19463_ net3940 net5895 net3906 vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or3b_4
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ net3443 net3960 net4642 net4748 _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a221o_1
X_13887_ _07034_ _07039_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__xnor2_1
X_16675_ net4194 _09741_ _09742_ _07998_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__a22o_1
X_18414_ net4724 net3604 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__xor2_1
X_15626_ _08682_ _08714_ _08713_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12838_ _05949_ _05956_ _05960_ _05957_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__o31a_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ net4976 _03268_ _03300_ _03299_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18345_ _02529_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15557_ _08353_ _08651_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__and2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12769_ net7727 _05903_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7909 _08455_ vssd1 vssd1 vccd1 vccd1 net8436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14508_ _07489_ _07194_ _07676_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__or3_1
X_15488_ _08581_ _08582_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__xnor2_4
X_18276_ net4038 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__buf_1
X_20667__13 clknet_1_0__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17227_ _10120_ _10121_ vssd1 vssd1 vccd1 vccd1 _10247_ sky130_fd_sc_hd__nor2_1
Xinput20 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
Xinput31 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_4
X_14439_ _07580_ _07603_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_1_1__f__03865_ clknet_0__03865_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03865_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput42 i_mode[2] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_4
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput53 i_vec_csb vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_6
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17158_ _10161_ _10177_ vssd1 vssd1 vccd1 vccd1 _10178_ sky130_fd_sc_hd__xnor2_1
Xhold804 net6400 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold815 _01254_ vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 net6443 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 _01272_ vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _09201_ _09202_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold848 net6368 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17089_ _10108_ _10109_ vssd1 vssd1 vccd1 vccd1 _10110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold859 net6175 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2205 _04281_ vssd1 vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2216 _01549_ vssd1 vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2227 net5727 vssd1 vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2238 net7420 vssd1 vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1504 _01420_ vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _01567_ vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1515 _01571_ vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _04259_ vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1537 net6895 vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1548 net6067 vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _04230_ vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21623_ clknet_leaf_101_i_clk net2181 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21554_ net188 net635 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20505_ clknet_1_1__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__buf_1
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21485_ clknet_leaf_48_i_clk net1297 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4130 net3856 vssd1 vssd1 vccd1 vccd1 net4657 sky130_fd_sc_hd__clkbuf_2
X_22106_ net168 net1607 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold4141 net7977 vssd1 vssd1 vccd1 vccd1 net4668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4152 net8202 vssd1 vssd1 vccd1 vccd1 net4679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4163 net4220 vssd1 vssd1 vccd1 vccd1 net4690 sky130_fd_sc_hd__clkbuf_2
X_20298_ net6378 net3816 _03814_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__mux2_1
Xhold4174 net763 vssd1 vssd1 vccd1 vccd1 net4701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3440 _04492_ vssd1 vssd1 vccd1 vccd1 net3967 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4185 net677 vssd1 vssd1 vccd1 vccd1 net4712 sky130_fd_sc_hd__dlygate4sd3_1
X_22037_ net479 net2386 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
Xhold4196 net3913 vssd1 vssd1 vccd1 vccd1 net4723 sky130_fd_sc_hd__clkbuf_2
Xhold3451 net7745 vssd1 vssd1 vccd1 vccd1 net3978 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_104_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold3462 _00463_ vssd1 vssd1 vccd1 vccd1 net3989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3473 net7703 vssd1 vssd1 vccd1 vccd1 net4000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3484 _08108_ vssd1 vssd1 vccd1 vccd1 net4011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2750 _03028_ vssd1 vssd1 vccd1 vccd1 net3277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3495 _01181_ vssd1 vssd1 vccd1 vccd1 net4022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2761 _01148_ vssd1 vssd1 vccd1 vccd1 net3288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2772 _03556_ vssd1 vssd1 vccd1 vccd1 net3299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2783 _00625_ vssd1 vssd1 vccd1 vccd1 net3310 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2794 _03562_ vssd1 vssd1 vccd1 vccd1 net3321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _06940_ _06941_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__xor2_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ net7846 _07952_ _07953_ net7785 vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__o211a_1
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ _06873_ _06876_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_119_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10953_ net6591 net6506 _04287_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16460_ _09542_ _09550_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__xor2_2
X_13672_ _06729_ _06793_ _06799_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__and3_1
X_10884_ net6094 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15411_ _08499_ _08504_ _08505_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ net22 vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__clkbuf_4
X_16391_ _09352_ _09481_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ _07989_ _07946_ _08003_ _07868_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__a211oi_1
X_18130_ net3757 net4379 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ _05708_ _05733_ _05734_ _05718_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11505_ net3461 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__inv_2
X_15273_ _08181_ _08366_ _08367_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__a21boi_1
X_18061_ _02278_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__xnor2_1
X_12485_ _05649_ _05666_ net7 vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17012_ _08542_ _09472_ vssd1 vssd1 vccd1 vccd1 _10033_ sky130_fd_sc_hd__or2_1
X_14224_ _07328_ _07330_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__xor2_1
X_11436_ rbzero.spi_registers.texadd3\[5\] rbzero.spi_registers.texadd1\[5\] rbzero.spi_registers.texadd0\[5\]
+ rbzero.spi_registers.texadd2\[5\] _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04628_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14155_ _07325_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11367_ rbzero.spi_registers.texadd3\[17\] rbzero.spi_registers.texadd1\[17\] rbzero.spi_registers.texadd0\[17\]
+ rbzero.spi_registers.texadd2\[17\] _04554_ _04555_ vssd1 vssd1 vccd1 vccd1 _04559_
+ sky130_fd_sc_hd__mux4_2
X_13106_ net4462 net3604 vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nand2_1
X_20648__376 clknet_1_1__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__inv_2
X_14086_ _07168_ _07214_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__or2b_1
X_18963_ net7367 net5771 net2874 vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11298_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__clkbuf_4
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20347__104 clknet_1_1__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__inv_2
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _01947_ _02151_ _02048_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a21o_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ net4610 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__inv_2
X_18894_ net6709 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17845_ _02081_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17776_ _01924_ _01918_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__or2b_1
X_14988_ net92 vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19515_ net1622 net5526 net3086 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16727_ _09750_ _09764_ vssd1 vssd1 vccd1 vccd1 _09765_ sky130_fd_sc_hd__or2_1
X_13939_ _06727_ net541 _07109_ _06693_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19446_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__clkbuf_2
X_16658_ _09736_ vssd1 vssd1 vccd1 vccd1 _09737_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_83_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15609_ _08657_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_45_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19377_ net5224 _03283_ _03291_ _03288_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16589_ _09674_ _09675_ _09677_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20393__146 clknet_1_0__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__inv_2
X_18328_ _02510_ _02515_ _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__o21a_1
Xhold7706 rbzero.traced_texa\[5\] vssd1 vssd1 vccd1 vccd1 net8233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7717 rbzero.debug_overlay.vplaneX\[-8\] vssd1 vssd1 vccd1 vccd1 net8244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7728 _02523_ vssd1 vssd1 vccd1 vccd1 net8255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7739 _08058_ vssd1 vssd1 vccd1 vccd1 net8266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ net4832 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21270_ clknet_leaf_27_i_clk net4311 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03848_ clknet_0__03848_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03848_
+ sky130_fd_sc_hd__clkbuf_16
Xhold601 net6204 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 net6234 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold623 _01031_ vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
X_20221_ _04459_ net3620 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold634 net5471 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 net4592 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold656 _03533_ vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 net2770 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_21_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20152_ rbzero.debug_overlay.facingY\[-9\] net3182 _03723_ vssd1 vssd1 vccd1 vccd1
+ _03729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold678 net4421 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold689 _01262_ vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2002 _01049_ vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2013 _04403_ vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2024 net7136 vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _09725_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__clkbuf_4
Xhold2035 _01569_ vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 net7245 vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 net6638 vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 net6714 vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 net3213 vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2068 rbzero.tex_g1\[4\] vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 _01511_ vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2079 _01378_ vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _00583_ vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 net6704 vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1356 _03399_ vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 net2816 vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1378 _00984_ vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
X_20661__7 clknet_1_1__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
Xhold1389 _03022_ vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20985_ clknet_leaf_29_i_clk net4125 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21606_ clknet_leaf_131_i_clk net2264 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21537_ net171 net2897 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _04751_ _05198_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nor2_1
X_21468_ clknet_leaf_23_i_clk net1479 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ net6032 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21399_ clknet_leaf_41_i_clk net3572 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11152_ _04264_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15960_ _09051_ _09053_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__nand2_1
X_11083_ net3093 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3270 net4920 vssd1 vssd1 vccd1 vccd1 net3797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3281 net7670 vssd1 vssd1 vccd1 vccd1 net3808 sky130_fd_sc_hd__dlygate4sd3_1
X_14911_ net8018 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__o21a_1
XFILLER_0_179_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3292 net7991 vssd1 vssd1 vccd1 vccd1 net3819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _08811_ _08856_ _08983_ _08985_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__a22o_2
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2580 net7485 vssd1 vssd1 vccd1 vccd1 net3107 sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _09373_ _10289_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nor2_1
Xhold2591 _04407_ vssd1 vssd1 vccd1 vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _07999_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03868_ clknet_0__03868_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03868_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1890 net7028 vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
X_17561_ _01688_ _01782_ _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ net4139 vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__inv_2
X_14773_ net4415 _07938_ _07872_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19300_ net1631 _03238_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__or2_1
X_16512_ _06124_ net4908 vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__nor2_1
X_10936_ net3264 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
X_13724_ _06870_ _06894_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17492_ net4659 net4653 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19231_ net5332 _03201_ _03207_ _03206_ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__o211a_1
X_16443_ _08401_ _08916_ _09292_ _09411_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__or4_1
X_10867_ net2292 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__clkbuf_1
X_13655_ _06822_ _06791_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__or2b_1
XFILLER_0_183_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ net47 _05763_ _05764_ clknet_leaf_89_i_clk vssd1 vssd1 vccd1 vccd1 _05786_
+ sky130_fd_sc_hd__a22o_2
X_19162_ net1997 _03146_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or2_1
X_16374_ _09349_ _09367_ _09365_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _06495_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__buf_2
X_10798_ net3170 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__clkbuf_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ net4565 net4403 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15325_ _08416_ _08419_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12537_ net13 net12 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__nor2_1
X_19093_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18044_ _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15256_ _08337_ _08350_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__and2b_1
X_12468_ net7 _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14207_ _07374_ _07375_ _07376_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__and3_1
X_11419_ _04496_ _04547_ _04610_ _04021_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a31oi_1
X_15187_ _08270_ _08272_ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__or2_1
X_12399_ rbzero.tex_b1\[35\] rbzero.tex_b1\[34\] _05250_ vssd1 vssd1 vccd1 vccd1 _05584_
+ sky130_fd_sc_hd__mux2_1
X_14138_ _07308_ _07303_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19995_ net4168 _03607_ net5746 _03339_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ net543 vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__clkbuf_4
X_18946_ net2974 net7083 _03036_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18877_ net3111 net5045 _03003_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ _02004_ _02065_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__xor2_2
XFILLER_0_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17759_ _01914_ _01970_ _01996_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20770_ net864 net5488 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401__153 clknet_1_0__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__inv_2
XFILLER_0_130_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19429_ net3519 _03122_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nand2_2
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7503 _00510_ vssd1 vssd1 vccd1 vccd1 net8030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7514 _08445_ vssd1 vssd1 vccd1 vccd1 net8041 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7525 _00001_ vssd1 vssd1 vccd1 vccd1 net8052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7536 _00634_ vssd1 vssd1 vccd1 vccd1 net8063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6802 _04048_ vssd1 vssd1 vccd1 vccd1 net7329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7547 _02582_ vssd1 vssd1 vccd1 vccd1 net8074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6813 net2783 vssd1 vssd1 vccd1 vccd1 net7340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7558 _02642_ vssd1 vssd1 vccd1 vccd1 net8085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6824 net2462 vssd1 vssd1 vccd1 vccd1 net7351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7569 rbzero.wall_tracer.rayAddendY\[-9\] vssd1 vssd1 vccd1 vccd1 net8096 sky130_fd_sc_hd__dlygate4sd3_1
X_21322_ clknet_leaf_12_i_clk net5127 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6835 rbzero.tex_b0\[51\] vssd1 vssd1 vccd1 vccd1 net7362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6846 net3169 vssd1 vssd1 vccd1 vccd1 net7373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6857 _04369_ vssd1 vssd1 vccd1 vccd1 net7384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6868 net3002 vssd1 vssd1 vccd1 vccd1 net7395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6879 rbzero.tex_b1\[17\] vssd1 vssd1 vccd1 vccd1 net7406 sky130_fd_sc_hd__dlygate4sd3_1
X_21253_ clknet_leaf_1_i_clk net3868 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold420 net5369 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _03156_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 net8233 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20204_ net4554 _03744_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
Xhold453 net5371 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 net8199 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold475 net8128 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
X_21184_ clknet_leaf_101_i_clk net3291 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold486 net5419 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold497 net5431 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20135_ rbzero.debug_overlay.facingX\[-4\] net3690 _03710_ vssd1 vssd1 vccd1 vccd1
+ _03718_ sky130_fd_sc_hd__mux2_1
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ net3252 _08177_ _03614_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__mux2_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _03032_ vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 net8155 vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _03438_ vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 net4897 vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 net6598 vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 _00929_ vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 net6539 vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1197 net6002 vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11770_ _04847_ _04959_ _04829_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ clknet_leaf_69_i_clk _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10721_ net2793 net6359 _04171_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__mux2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20899_ clknet_leaf_32_i_clk net5607 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20376__130 clknet_1_1__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__inv_2
XFILLER_0_166_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ _06492_ _06608_ _06610_ _06564_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__a211o_1
X_10652_ net7017 net6651 _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13371_ _06466_ _06469_ _06471_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__nand3_2
XFILLER_0_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ net5558 net5550 _04097_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _05237_ vssd1 vssd1 vccd1 vccd1 _05508_
+ sky130_fd_sc_hd__mux2_1
X_15110_ net3459 _08136_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__or2_2
X_16090_ _09179_ _09183_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15041_ net3774 _04485_ _06117_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__or3b_4
X_12253_ _04947_ _05435_ _05437_ _05439_ _04942_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11204_ net7109 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__clkbuf_1
X_12184_ net4080 _05021_ _05015_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18800_ net5955 _02945_ _02536_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
X_11135_ net2649 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
X_16992_ net4589 net4483 vssd1 vssd1 vccd1 vccd1 _10013_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _02862_ _02864_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__and2_1
X_11066_ net1889 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
X_15943_ _09036_ _09037_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__xor2_2
X_18662_ _02812_ _02817_ _04480_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _08957_ _08963_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _01779_ _01744_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__or2b_1
XFILLER_0_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _07959_ vssd1 vssd1 vccd1 vccd1 _07984_ sky130_fd_sc_hd__inv_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18593_ net4423 net652 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__nand2_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20459__205 clknet_1_0__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__inv_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _01784_ _01760_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__nor2_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14756_ net7843 _07821_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11968_ rbzero.debug_overlay.vplaneX\[-6\] _05102_ _05090_ rbzero.debug_overlay.vplaneX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _06873_ _06876_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a21bo_1
X_17475_ _01714_ _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__xor2_1
X_10919_ net6856 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__buf_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ _05077_ net4118 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__nand2_2
X_14687_ _07841_ _07852_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__a21oi_1
X_19214_ net5336 _03167_ _03195_ _03189_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__o211a_1
X_16426_ _09515_ _09516_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13638_ _06715_ net544 _06739_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19145_ net957 _03147_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__or2_1
X_16357_ _09336_ _09448_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ _06733_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__xnor2_1
Xhold6109 rbzero.tex_b1\[9\] vssd1 vssd1 vccd1 vccd1 net6636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15308_ _08368_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19076_ net3793 net6611 _09725_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
X_16288_ _08306_ _08392_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5408 net3849 vssd1 vssd1 vccd1 vccd1 net5935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5419 net3917 vssd1 vssd1 vccd1 vccd1 net5946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18027_ _02261_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15239_ _08280_ _08326_ _08327_ _08333_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__o31a_2
Xhold4707 net871 vssd1 vssd1 vccd1 vccd1 net5234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4718 _00795_ vssd1 vssd1 vccd1 vccd1 net5245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4729 net922 vssd1 vssd1 vccd1 vccd1 net5256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19978_ net3200 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18929_ net3298 net7593 _03025_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21940_ net382 net2404 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21871_ net313 net1922 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20822_ _03980_ _03982_ _03984_ _09720_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a31o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20753_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7300 net4480 vssd1 vssd1 vccd1 vccd1 net7827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7344 net3460 vssd1 vssd1 vccd1 vccd1 net7871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7355 net4203 vssd1 vssd1 vccd1 vccd1 net7882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6610 net2551 vssd1 vssd1 vccd1 vccd1 net7137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7366 rbzero.traced_texVinit\[5\] vssd1 vssd1 vccd1 vccd1 net7893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6621 rbzero.tex_r0\[23\] vssd1 vssd1 vccd1 vccd1 net7148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6632 net2209 vssd1 vssd1 vccd1 vccd1 net7159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7377 net3492 vssd1 vssd1 vccd1 vccd1 net7904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6643 rbzero.tex_g1\[22\] vssd1 vssd1 vccd1 vccd1 net7170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7388 rbzero.wall_tracer.stepDistY\[-9\] vssd1 vssd1 vccd1 vccd1 net7915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6654 _04208_ vssd1 vssd1 vccd1 vccd1 net7181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7399 net4319 vssd1 vssd1 vccd1 vccd1 net7926 sky130_fd_sc_hd__dlygate4sd3_1
X_21305_ clknet_leaf_12_i_clk net5326 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6665 net2465 vssd1 vssd1 vccd1 vccd1 net7192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5920 rbzero.spi_registers.new_texadd\[0\]\[4\] vssd1 vssd1 vccd1 vccd1 net6447
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6676 rbzero.tex_b0\[52\] vssd1 vssd1 vccd1 vccd1 net7203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5931 net1314 vssd1 vssd1 vccd1 vccd1 net6458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6687 net2858 vssd1 vssd1 vccd1 vccd1 net7214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5942 rbzero.spi_registers.new_texadd\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net6469
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5953 net1258 vssd1 vssd1 vccd1 vccd1 net6480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6698 rbzero.tex_r1\[14\] vssd1 vssd1 vccd1 vccd1 net7225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5964 rbzero.spi_registers.new_texadd\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net6491
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 net8151 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21236_ clknet_leaf_13_i_clk net4032 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5975 net1273 vssd1 vssd1 vccd1 vccd1 net6502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold261 net5138 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5986 _03019_ vssd1 vssd1 vccd1 vccd1 net6513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5997 net1408 vssd1 vssd1 vccd1 vccd1 net6524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 net5239 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 net2363 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 net5225 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
X_21167_ clknet_leaf_132_i_clk net2470 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20118_ _03123_ _03605_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nand2_4
XFILLER_0_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21098_ clknet_leaf_5_i_clk net1679 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20408__159 clknet_1_1__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__inv_2
XFILLER_0_77_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20049_ _03651_ _03652_ _03653_ net3683 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o22a_1
X_12940_ _06056_ net4645 vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nor2_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _06036_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__and2_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 net4705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _07606_ _07608_ _07556_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__a21o_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11822_ _04909_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__and2_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _08273_ _08281_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__xnor2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _04847_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14541_ _07413_ _07327_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__nor2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ net6963 net2143 _04160_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__mux2_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17260_ _10150_ _10278_ vssd1 vssd1 vccd1 vccd1 _10279_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ _07631_ _07642_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__xor2_2
X_11684_ _04854_ _04855_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _09171_ _09178_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10635_ net6669 net2423 _04127_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__mux2_1
X_13423_ _06530_ _06532_ _06461_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ _08391_ vssd1 vssd1 vccd1 vccd1 _10211_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _09233_ _09234_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13354_ _06519_ _06521_ net554 _06524_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__or4bb_4
X_10566_ net7266 net7324 _04086_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12305_ _04976_ _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16073_ _09164_ _09166_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13285_ _06306_ _06338_ _06341_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__a21o_2
X_10497_ net7063 net2657 _04053_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12236_ _05204_ _05420_ _05422_ _04955_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__o211a_1
X_15024_ _08118_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__buf_4
X_19901_ net1152 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19832_ net6663 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
X_12167_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _05249_ vssd1 vssd1 vccd1 vccd1 _05355_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ net6958 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
X_16975_ _09930_ _09996_ vssd1 vssd1 vccd1 vccd1 _09997_ sky130_fd_sc_hd__xnor2_2
X_12098_ net1822 _04991_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18714_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__clkbuf_4
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net2707 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
X_15926_ _08389_ _08509_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19694_ net6422 net3592 _03468_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__mux2_1
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18645_ _02794_ net4771 net8025 _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08941_ _08945_ _08951_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__o21a_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14808_ _07969_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18576_ _09761_ _09753_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__nand2_1
X_15788_ _08879_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__xnor2_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17527_ _01761_ _10437_ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14739_ net7843 _07887_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17458_ _01691_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16409_ _09379_ _09387_ _09499_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__a21bo_1
X_17389_ _10295_ _10296_ _10294_ vssd1 vssd1 vccd1 vccd1 _10407_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19128_ net886 _03140_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__nand2_2
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20513__254 clknet_1_0__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__inv_2
Xhold5205 net2742 vssd1 vssd1 vccd1 vccd1 net5732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5216 net4362 vssd1 vssd1 vccd1 vccd1 net5743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19059_ net7581 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__clkbuf_1
Xhold5227 rbzero.map_overlay.i_otherx\[0\] vssd1 vssd1 vccd1 vccd1 net5754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5238 _03070_ vssd1 vssd1 vccd1 vccd1 net5765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4504 net700 vssd1 vssd1 vccd1 vccd1 net5031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5249 _02878_ vssd1 vssd1 vccd1 vccd1 net5776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4515 _00856_ vssd1 vssd1 vccd1 vccd1 net5042 sky130_fd_sc_hd__dlygate4sd3_1
X_22070_ net512 net2467 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold4526 net713 vssd1 vssd1 vccd1 vccd1 net5053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4537 rbzero.spi_registers.texadd0\[16\] vssd1 vssd1 vccd1 vccd1 net5064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3803 net3434 vssd1 vssd1 vccd1 vccd1 net4330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4548 net726 vssd1 vssd1 vccd1 vccd1 net5075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3814 net8314 vssd1 vssd1 vccd1 vccd1 net4341 sky130_fd_sc_hd__dlygate4sd3_1
X_21021_ clknet_leaf_54_i_clk net4241 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4559 _00842_ vssd1 vssd1 vccd1 vccd1 net5086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3825 net7937 vssd1 vssd1 vccd1 vccd1 net4352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3836 _03674_ vssd1 vssd1 vccd1 vccd1 net4363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3847 net5736 vssd1 vssd1 vccd1 vccd1 net4374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3858 _00776_ vssd1 vssd1 vccd1 vccd1 net4385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3869 net8381 vssd1 vssd1 vccd1 vccd1 net4396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21923_ net365 net1181 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21854_ net296 net2847 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _03970_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and2b_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21785_ clknet_leaf_1_i_clk net1364 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20736_ net5340 _03877_ _03874_ _03913_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7130 _03504_ vssd1 vssd1 vccd1 vccd1 net7657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7141 rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 net7668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7152 _04664_ vssd1 vssd1 vccd1 vccd1 net7679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7163 net3326 vssd1 vssd1 vccd1 vccd1 net7690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7174 net3431 vssd1 vssd1 vccd1 vccd1 net7701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6440 net2324 vssd1 vssd1 vccd1 vccd1 net6967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7185 net4033 vssd1 vssd1 vccd1 vccd1 net7712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6451 rbzero.tex_r0\[17\] vssd1 vssd1 vccd1 vccd1 net6978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7196 _05298_ vssd1 vssd1 vccd1 vccd1 net7723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6462 net2619 vssd1 vssd1 vccd1 vccd1 net6989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20488__231 clknet_1_1__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__inv_2
XFILLER_0_182_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6473 rbzero.tex_g1\[30\] vssd1 vssd1 vccd1 vccd1 net7000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6484 net2248 vssd1 vssd1 vccd1 vccd1 net7011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6495 rbzero.tex_b0\[6\] vssd1 vssd1 vccd1 vccd1 net7022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5750 net1206 vssd1 vssd1 vccd1 vccd1 net6277 sky130_fd_sc_hd__dlygate4sd3_1
X_13070_ net2277 _06244_ _06054_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5761 _03413_ vssd1 vssd1 vccd1 vccd1 net6288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5772 net1241 vssd1 vssd1 vccd1 vccd1 net6299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5783 _03824_ vssd1 vssd1 vccd1 vccd1 net6310 sky130_fd_sc_hd__dlygate4sd3_1
X_12021_ rbzero.tex_r1\[1\] rbzero.tex_r1\[0\] _04838_ vssd1 vssd1 vccd1 vccd1 _05210_
+ sky130_fd_sc_hd__mux2_1
X_21219_ clknet_leaf_120_i_clk net3100 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5794 net1266 vssd1 vssd1 vccd1 vccd1 net6321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16760_ _09791_ _08978_ _09792_ vssd1 vssd1 vccd1 vccd1 _09793_ sky130_fd_sc_hd__o21a_2
X_13972_ _07094_ _07097_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__xor2_1
X_15711_ _08692_ _08798_ _08800_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__and3_1
X_12923_ net4393 net3848 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xor2_1
X_16691_ net8123 _09743_ _09744_ net4293 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18430_ net3494 net4501 _02609_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15642_ _08736_ _08711_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__xnor2_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ net7575 vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11805_ _04832_ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__or2_1
X_18361_ rbzero.wall_tracer.rayAddendX\[-3\] _02547_ _02537_ vssd1 vssd1 vccd1 vccd1
+ _02548_ sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _08159_ _08157_ net7835 _08147_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__nand2_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _10321_ _10329_ vssd1 vssd1 vccd1 vccd1 _10331_ sky130_fd_sc_hd__or2_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _07691_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__nand2_1
X_11736_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _04912_ vssd1 vssd1 vccd1 vccd1 _04926_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ net1436 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17243_ net4610 net4405 vssd1 vssd1 vccd1 vccd1 _10262_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _07623_ _07622_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ net2910 _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or2_1
X_13406_ _06576_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__inv_2
X_10618_ net7184 net5706 _04116_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__mux2_1
X_17174_ _08326_ _09170_ vssd1 vssd1 vccd1 vccd1 _10194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11598_ _04785_ _04784_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__nand2_1
X_14386_ _07455_ _07505_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _08618_ _09066_ _09128_ _09126_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ net5730 net6872 _04075_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13337_ net570 _06470_ _06441_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ _09131_ _09132_ _09149_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13268_ net8217 _06314_ _06316_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__a21o_1
X_15007_ _04567_ net3986 _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__mux2_1
X_12219_ _04943_ _05403_ _05405_ _04947_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__o211a_1
X_13199_ _06368_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__xnor2_4
Xhold2409 _01124_ vssd1 vssd1 vccd1 vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1708 net7056 vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 _01462_ vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16958_ _09973_ _09977_ _09978_ vssd1 vssd1 vccd1 vccd1 _09980_ sky130_fd_sc_hd__a21o_1
XFILLER_0_205_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15909_ _09002_ _09003_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__nand2_1
X_19677_ net6532 net3816 _03457_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
X_16889_ _09617_ _09909_ vssd1 vssd1 vccd1 vccd1 _09911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18628_ _02526_ _02779_ _02780_ _02785_ _02786_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18559_ net3807 _06244_ _06050_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21570_ net204 net2843 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 _07903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 net8002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_56 _04911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_89 net2094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5002 net1818 vssd1 vssd1 vccd1 vccd1 net5529 sky130_fd_sc_hd__dlygate4sd3_1
X_20383_ clknet_1_1__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__buf_1
Xhold5013 net1736 vssd1 vssd1 vccd1 vccd1 net5540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5024 _04100_ vssd1 vssd1 vccd1 vccd1 net5551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5035 net1402 vssd1 vssd1 vccd1 vccd1 net5562 sky130_fd_sc_hd__dlygate4sd3_1
X_22122_ clknet_leaf_54_i_clk net4974 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
Xhold4301 net3529 vssd1 vssd1 vccd1 vccd1 net4828 sky130_fd_sc_hd__clkbuf_2
Xhold5046 net2186 vssd1 vssd1 vccd1 vccd1 net5573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5057 rbzero.wall_tracer.trackDistX\[6\] vssd1 vssd1 vccd1 vccd1 net5584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4312 _00638_ vssd1 vssd1 vccd1 vccd1 net4839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4323 net893 vssd1 vssd1 vccd1 vccd1 net4850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5068 rbzero.row_render.texu\[4\] vssd1 vssd1 vccd1 vccd1 net5595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5079 _00386_ vssd1 vssd1 vccd1 vccd1 net5606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4334 net5958 vssd1 vssd1 vccd1 vccd1 net4861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4345 rbzero.wall_tracer.trackDistX\[-9\] vssd1 vssd1 vccd1 vccd1 net4872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3600 _04712_ vssd1 vssd1 vccd1 vccd1 net4127 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22053_ net495 net1757 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold4356 net917 vssd1 vssd1 vccd1 vccd1 net4883 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3611 net4070 vssd1 vssd1 vccd1 vccd1 net4138 sky130_fd_sc_hd__clkbuf_4
Xhold3622 _05379_ vssd1 vssd1 vccd1 vccd1 net4149 sky130_fd_sc_hd__clkbuf_4
Xhold3633 net4094 vssd1 vssd1 vccd1 vccd1 net4160 sky130_fd_sc_hd__clkbuf_4
Xhold4378 rbzero.wall_tracer.trackDistY\[-4\] vssd1 vssd1 vccd1 vccd1 net4905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3644 _05173_ vssd1 vssd1 vccd1 vccd1 net4171 sky130_fd_sc_hd__dlygate4sd3_1
X_21004_ clknet_leaf_85_i_clk _00491_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4389 net3756 vssd1 vssd1 vccd1 vccd1 net4916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2910 _03717_ vssd1 vssd1 vccd1 vccd1 net3437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3655 _04511_ vssd1 vssd1 vccd1 vccd1 net4182 sky130_fd_sc_hd__buf_1
Xhold2921 net7576 vssd1 vssd1 vccd1 vccd1 net3448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3666 net8296 vssd1 vssd1 vccd1 vccd1 net4193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3677 net7883 vssd1 vssd1 vccd1 vccd1 net4204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2932 net7867 vssd1 vssd1 vccd1 vccd1 net3459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3688 net7895 vssd1 vssd1 vccd1 vccd1 net4215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2943 net5761 vssd1 vssd1 vccd1 vccd1 net3470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2954 net7596 vssd1 vssd1 vccd1 vccd1 net3481 sky130_fd_sc_hd__clkbuf_2
Xhold3699 net8069 vssd1 vssd1 vccd1 vccd1 net4226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2965 net7903 vssd1 vssd1 vccd1 vccd1 net3492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2987 _02569_ vssd1 vssd1 vccd1 vccd1 net3514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2998 net5806 vssd1 vssd1 vccd1 vccd1 net3525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21906_ net348 net805 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21837_ net279 net2737 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12570_ _05749_ net4156 vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21768_ clknet_leaf_10_i_clk net1557 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20719_ _03894_ _03895_ _03896_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ net4126 net2038 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21699_ clknet_leaf_116_i_clk net4346 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _07374_ _07375_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ rbzero.spi_registers.texadd1\[1\] _04548_ _04643_ vssd1 vssd1 vccd1 vccd1
+ _04644_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14171_ net5902 _07304_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__and2_4
XFILLER_0_151_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11383_ rbzero.spi_registers.texadd0\[22\] _04545_ _04574_ vssd1 vssd1 vccd1 vccd1
+ _04575_ sky130_fd_sc_hd__o21ai_1
Xhold6270 _04180_ vssd1 vssd1 vccd1 vccd1 net6797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6281 net1961 vssd1 vssd1 vccd1 vccd1 net6808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _06286_ _06289_ _06287_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__o21ba_1
Xhold6292 _04179_ vssd1 vssd1 vccd1 vccd1 net6819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5580 net924 vssd1 vssd1 vccd1 vccd1 net6107 sky130_fd_sc_hd__dlygate4sd3_1
X_17930_ _01784_ _09540_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__nor2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _06218_ _06228_ _06214_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a21oi_1
Xhold5591 net997 vssd1 vssd1 vccd1 vccd1 net6118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12004_ net4095 _04600_ _04467_ net4127 vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__o2bb2a_1
X_17861_ _08472_ _09225_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4890 _00780_ vssd1 vssd1 vccd1 vccd1 net5417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16812_ _09839_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__clkbuf_1
X_19600_ net3844 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17792_ _02014_ _02015_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19531_ net2953 net7524 net3086 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
X_16743_ _09768_ _09777_ _09778_ _09769_ net5472 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13955_ _07120_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__xnor2_2
X_20542__280 clknet_1_1__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__inv_2
X_19462_ net3907 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
X_12906_ net3326 _06061_ _06032_ net3473 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a22o_1
X_16674_ net4341 _09741_ _09742_ _07991_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a22o_1
X_13886_ _07049_ _07054_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18413_ _02559_ net4726 net8076 net3639 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a31o_1
X_15625_ _08716_ _08719_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12837_ _05999_ _06002_ _06006_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__or4_1
X_19393_ net1386 _03270_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _02530_ _02531_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15556_ _08144_ _08352_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ net39 _05911_ _05920_ _05900_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__o221a_2
XFILLER_0_167_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _07676_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__xnor2_1
X_11719_ net42 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__inv_2
X_18275_ net1282 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__clkbuf_1
X_15487_ _08211_ _08200_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ net32 _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17226_ _10146_ _10245_ vssd1 vssd1 vccd1 vccd1 _10246_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_2
X_14438_ _07560_ _07605_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__xor2_4
Xclkbuf_1_1__f__03864_ clknet_0__03864_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03864_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
Xinput32 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_2
Xinput43 i_reg_csb vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_6
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_6
XFILLER_0_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17157_ _10175_ _10176_ vssd1 vssd1 vccd1 vccd1 _10177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _07413_ _07280_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__nor2_1
Xhold805 net6402 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 net6190 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ _09199_ _09200_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__nand2_1
Xhold827 _01321_ vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 net2097 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _09979_ _09981_ _10107_ vssd1 vssd1 vccd1 vccd1 _10109_ sky130_fd_sc_hd__and3_1
Xhold849 _00971_ vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16039_ _08253_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2206 _01375_ vssd1 vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2217 net7269 vssd1 vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2228 net7237 vssd1 vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20625__355 clknet_1_0__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__inv_2
Xhold2239 _00649_ vssd1 vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1505 net7128 vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1516 net7018 vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _01394_ vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 _01328_ vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 net6069 vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19729_ net7673 net5496 _03489_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21622_ clknet_leaf_128_i_clk net3024 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ net187 net2681 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21484_ clknet_leaf_44_i_clk net1376 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20370__125 clknet_1_1__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__inv_2
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4120 _06161_ vssd1 vssd1 vccd1 vccd1 net4647 sky130_fd_sc_hd__dlygate4sd3_1
X_22105_ net167 net2350 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
Xhold4131 net7979 vssd1 vssd1 vccd1 vccd1 net4658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4142 net3869 vssd1 vssd1 vccd1 vccd1 net4669 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4153 _00414_ vssd1 vssd1 vccd1 vccd1 net4680 sky130_fd_sc_hd__dlygate4sd3_1
X_20297_ net1264 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
Xhold4164 _08056_ vssd1 vssd1 vccd1 vccd1 net4691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3430 _09726_ vssd1 vssd1 vccd1 vccd1 net3957 sky130_fd_sc_hd__dlygate4sd3_1
X_22036_ net478 net1144 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
Xhold4186 net8244 vssd1 vssd1 vccd1 vccd1 net4713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3441 net5780 vssd1 vssd1 vccd1 vccd1 net3968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4197 rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 net4724 sky130_fd_sc_hd__clkbuf_2
Xhold3452 _03395_ vssd1 vssd1 vccd1 vccd1 net3979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3463 rbzero.debug_overlay.playerX\[1\] vssd1 vssd1 vccd1 vccd1 net3990 sky130_fd_sc_hd__buf_2
Xhold3474 _00621_ vssd1 vssd1 vccd1 vccd1 net4001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2740 _03065_ vssd1 vssd1 vccd1 vccd1 net3267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3485 _08109_ vssd1 vssd1 vccd1 vccd1 net4012 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2751 _00678_ vssd1 vssd1 vccd1 vccd1 net3278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3496 net5980 vssd1 vssd1 vccd1 vccd1 net4023 sky130_fd_sc_hd__buf_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2762 net7547 vssd1 vssd1 vccd1 vccd1 net3289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2773 _01121_ vssd1 vssd1 vccd1 vccd1 net3300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2784 rbzero.pov.spi_buffer\[56\] vssd1 vssd1 vccd1 vccd1 net3311 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2795 _01126_ vssd1 vssd1 vccd1 vccd1 net3322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13740_ _06865_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10952_ net2266 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13671_ _06797_ _06798_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883_ net6092 net2575 _04253_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15410_ _08488_ _08490_ _08498_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__nand3_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ net27 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__inv_2
X_16390_ _08864_ _09354_ vssd1 vssd1 vccd1 vccd1 _09481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15341_ _06632_ _07988_ _07990_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__o21ba_1
X_12553_ _04468_ _04023_ _05691_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18060_ _02294_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__xnor2_1
X_11504_ net4102 _04692_ net8193 net3955 _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o221a_1
X_15272_ net4373 _06120_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12484_ net51 _05646_ _05642_ net40 _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17011_ _10029_ _10031_ vssd1 vssd1 vccd1 vccd1 _10032_ sky130_fd_sc_hd__nand2_1
X_14223_ net8355 _07387_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_62_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ rbzero.spi_registers.texadd3\[4\] rbzero.spi_registers.texadd1\[4\] rbzero.spi_registers.texadd0\[4\]
+ rbzero.spi_registers.texadd2\[4\] _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04627_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14154_ _07147_ _07324_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__or2_1
X_11366_ _04553_ _04556_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ _06273_ _06274_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__o21a_2
Xclkbuf_leaf_2_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14085_ _07254_ _07255_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__or2_1
X_18962_ net5712 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
X_11297_ _04023_ _04469_ _04026_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__o21ai_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _01962_ _01963_ _02046_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a21o_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ net4651 vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__inv_2
X_18893_ net3155 net6707 _03003_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
X_17844_ _10327_ _01693_ _10346_ _08799_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_156_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17775_ _01807_ _01923_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nand2_1
X_14987_ _08091_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
X_19514_ net3085 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16726_ _09751_ _09752_ _09762_ _09763_ vssd1 vssd1 vccd1 vccd1 _09764_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13938_ net3533 vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19445_ net3978 _03123_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16657_ _09735_ vssd1 vssd1 vccd1 vccd1 _09736_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13869_ _07034_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15608_ _08690_ _08701_ _08702_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_174_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19376_ net6570 _03284_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
X_16588_ _09674_ _09675_ _09677_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__nand3_1
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18327_ net4733 net4887 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15539_ _08631_ _08632_ _08633_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7707 rbzero.traced_texa\[-9\] vssd1 vssd1 vccd1 vccd1 net8234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7718 rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 net8245 sky130_fd_sc_hd__dlygate4sd3_1
X_18258_ net3770 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17209_ _10226_ _10227_ _10228_ vssd1 vssd1 vccd1 vccd1 _10229_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03847_ clknet_0__03847_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03847_
+ sky130_fd_sc_hd__clkbuf_16
X_18189_ _02401_ _02409_ _02407_ _02408_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 _01453_ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 net6236 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20220_ net3619 net1573 _03709_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 net3319 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 net5473 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 net6210 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _01100_ vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold668 _03007_ vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
X_20151_ _04458_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__clkbuf_4
Xhold679 net6276 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2003 net6982 vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
X_20082_ net5771 _03485_ _03662_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2014 _01072_ vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _04200_ vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2036 net6853 vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2047 _01070_ vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _01286_ vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19805__82 clknet_1_0__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__inv_2
Xhold1313 net6716 vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _03038_ vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2069 net7352 vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 net8147 vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__buf_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1335 net6680 vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 _04304_ vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1357 _00943_ vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1368 _04126_ vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1379 net5749 vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ clknet_leaf_30_i_clk _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_178_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21605_ clknet_leaf_130_i_clk net1581 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21536_ net170 net2837 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21467_ clknet_leaf_18_i_clk net1294 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11220_ net6030 net2679 _04434_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21398_ clknet_leaf_41_i_clk net5358 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11151_ net6997 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11082_ net6846 net7322 _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux2_1
Xhold3260 net3354 vssd1 vssd1 vccd1 vccd1 net3787 sky130_fd_sc_hd__clkbuf_2
X_22019_ net461 net2952 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
X_14910_ _06239_ vssd1 vssd1 vccd1 vccd1 _08050_ sky130_fd_sc_hd__clkbuf_4
Xhold3271 _09860_ vssd1 vssd1 vccd1 vccd1 net3798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3282 _00616_ vssd1 vssd1 vccd1 vccd1 net3809 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _08811_ _08984_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__xnor2_4
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3293 net3421 vssd1 vssd1 vccd1 vccd1 net3820 sky130_fd_sc_hd__clkbuf_2
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2570 _01122_ vssd1 vssd1 vccd1 vccd1 net3097 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2581 net7487 vssd1 vssd1 vccd1 vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
X_14841_ net4481 _07998_ _07976_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__mux2_1
Xhold2592 _01068_ vssd1 vssd1 vccd1 vccd1 net3119 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03867_ clknet_0__03867_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03867_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1880 _01501_ vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
X_17560_ _01790_ _01800_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1891 net7030 vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
X_14772_ _07931_ _07933_ _07937_ net7824 net4704 vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__a221o_2
X_11984_ _05097_ net4170 _05120_ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16511_ _09224_ _08542_ _09133_ _09600_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__a2bb2o_1
X_13723_ _06867_ _06869_ _06868_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__a21bo_1
X_10935_ net7484 net7232 _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__mux2_1
X_17491_ net4659 net4653 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19230_ net6313 _03203_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__or2_1
X_16442_ _09523_ _09532_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13654_ _06712_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__xnor2_1
X_10866_ net7145 net7131 _04171_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12605_ net55 _05764_ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19161_ net5420 _03144_ _03164_ _03160_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__o211a_1
X_16373_ _09342_ _09368_ _09463_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__a21bo_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20654__381 clknet_1_0__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__inv_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ net83 _06576_ _06754_ _06755_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__or4_2
X_10797_ net6168 net7373 _04205_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ net4565 net4403 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15324_ _08417_ _08418_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__nor2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ net53 _05699_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a21o_1
X_19092_ net3996 _05730_ net4097 _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__and4b_1
XFILLER_0_164_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18043_ _01784_ _09540_ _02166_ _02170_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__o31a_1
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15255_ _08339_ _08348_ _08349_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__a21o_2
XFILLER_0_48_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12467_ net6 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14206_ _07374_ _07375_ _07376_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__a21oi_1
X_11418_ _04513_ _04543_ _04546_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15186_ _08266_ _08280_ vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__or2_2
XFILLER_0_151_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _05250_ vssd1 vssd1 vccd1 vccd1 _05583_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14137_ _06796_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__clkbuf_4
X_11349_ _04511_ _04512_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__nor2_1
X_19994_ net5745 _03485_ _03609_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18945_ net2331 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
X_14068_ _07237_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ net4655 _06192_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18876_ net2957 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _09272_ _01922_ _01920_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17758_ _01914_ _01970_ _01996_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ net7667 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__clkbuf_1
X_17689_ _01927_ _01928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19428_ net3653 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19359_ net6265 _03271_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__or2_1
Xhold7504 net4275 vssd1 vssd1 vccd1 vccd1 net8031 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_103_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_190_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7515 _08446_ vssd1 vssd1 vccd1 vccd1 net8042 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_165_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7526 net4812 vssd1 vssd1 vccd1 vccd1 net8053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6803 net2439 vssd1 vssd1 vccd1 vccd1 net7330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7548 _02585_ vssd1 vssd1 vccd1 vccd1 net8075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6814 rbzero.tex_b1\[4\] vssd1 vssd1 vccd1 vccd1 net7341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7559 _02646_ vssd1 vssd1 vccd1 vccd1 net8086 sky130_fd_sc_hd__dlygate4sd3_1
X_21321_ clknet_leaf_14_i_clk net5334 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6825 _04243_ vssd1 vssd1 vccd1 vccd1 net7352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6836 net2539 vssd1 vssd1 vccd1 vccd1 net7363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6847 rbzero.tex_b0\[3\] vssd1 vssd1 vccd1 vccd1 net7374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6858 net2558 vssd1 vssd1 vccd1 vccd1 net7385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6869 rbzero.tex_g0\[40\] vssd1 vssd1 vccd1 vccd1 net7396 sky130_fd_sc_hd__dlygate4sd3_1
X_21252_ clknet_leaf_0_i_clk net3676 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold410 net5237 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold421 net8119 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_118_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold432 net4367 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 net8017 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
X_20203_ net3496 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
Xhold454 net5373 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21183_ clknet_leaf_127_i_clk net1224 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold465 net8090 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 net4532 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 net5421 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
X_20134_ net3437 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
Xhold498 net5433 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20482__226 clknet_1_1__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__inv_2
XFILLER_0_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20065_ net3489 _03660_ net4618 _03628_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__o211a_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 net6573 vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _00682_ vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 net5515 vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 _00973_ vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1154 net4759 vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 _03464_ vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 net5825 vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _01055_ vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _03349_ vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ clknet_leaf_69_i_clk _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10720_ net5603 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20898_ clknet_4_7__leaf_i_clk net4813 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ _04104_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ net5552 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__clkbuf_1
X_13370_ _06516_ net562 vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__and2_1
X_12321_ _05233_ _05502_ _05506_ _04942_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21519_ clknet_leaf_7_i_clk net1327 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ _07870_ net8365 _08114_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__mux2_2
X_12252_ _04977_ _05438_ net87 vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11203_ net7107 net2962 _04423_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12183_ _05031_ _05370_ net4080 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ net2648 net6026 _04390_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__mux2_1
X_16991_ _10012_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__clkbuf_1
X_11065_ net5649 net6866 _04353_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__mux2_1
X_15942_ _08450_ _08464_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__nand2_1
X_18730_ net8060 _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__and2_1
Xhold3090 net8327 vssd1 vssd1 vccd1 vccd1 net3617 sky130_fd_sc_hd__dlygate4sd3_1
X_18661_ _02813_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _08965_ _08966_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__and2_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _01849_ _01850_ _09845_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a21o_1
X_14824_ _07944_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _05164_ net681 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_97_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _08140_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _07920_ _07921_ net7839 vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__mux2_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ net3493 _05080_ _05103_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1
+ vccd1 _05156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _06708_ _06815_ _06874_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__or3_4
X_17474_ _10275_ _10370_ _01715_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a21oi_1
X_10918_ net6854 net3176 _04276_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14686_ net7811 _07856_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__and2_1
X_11898_ net4117 _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16425_ _09513_ _09514_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19213_ net1331 _03169_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__or2_1
X_13637_ _06732_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__buf_6
X_10849_ net6225 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19144_ net2587 _03145_ net5614 _03149_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__o211a_1
X_16356_ _09446_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__xnor2_4
X_13568_ _06735_ _06738_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15307_ net8414 vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19075_ net1728 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12519_ net10 net11 vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__and2b_2
X_16287_ _09377_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_35_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ _06493_ _06608_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5409 rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 net5936 sky130_fd_sc_hd__dlygate4sd3_1
X_18026_ _02188_ _02217_ _02218_ _02186_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ _08330_ _08332_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4708 rbzero.spi_registers.texadd0\[2\] vssd1 vssd1 vccd1 vccd1 net5235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4719 net807 vssd1 vssd1 vccd1 vccd1 net5246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15169_ _08156_ _08263_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19977_ net53 net3199 _03109_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18928_ net3274 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18859_ net3352 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21870_ net312 net2019 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20821_ _03980_ _03982_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a21oi_1
X_20752_ _03924_ _03925_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7312 _06606_ vssd1 vssd1 vccd1 vccd1 net7839 sky130_fd_sc_hd__clkbuf_2
Xhold7323 _06557_ vssd1 vssd1 vccd1 vccd1 net7850 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold7334 rbzero.traced_texVinit\[0\] vssd1 vssd1 vccd1 vccd1 net7861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6600 net2680 vssd1 vssd1 vccd1 vccd1 net7127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7345 rbzero.wall_tracer.stepDistX\[-11\] vssd1 vssd1 vccd1 vccd1 net7872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6611 _04199_ vssd1 vssd1 vccd1 vccd1 net7138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7356 net941 vssd1 vssd1 vccd1 vccd1 net7883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7367 net4214 vssd1 vssd1 vccd1 vccd1 net7894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6622 net2294 vssd1 vssd1 vccd1 vccd1 net7149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6633 rbzero.tex_r1\[43\] vssd1 vssd1 vccd1 vccd1 net7160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7378 rbzero.row_render.size\[1\] vssd1 vssd1 vccd1 vccd1 net7905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6644 net2402 vssd1 vssd1 vccd1 vccd1 net7171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7389 net4398 vssd1 vssd1 vccd1 vccd1 net7916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6655 net2570 vssd1 vssd1 vccd1 vccd1 net7182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5910 _03030_ vssd1 vssd1 vccd1 vccd1 net6437 sky130_fd_sc_hd__dlygate4sd3_1
X_21304_ clknet_leaf_47_i_clk net5242 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6666 rbzero.tex_g0\[14\] vssd1 vssd1 vccd1 vccd1 net7193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5921 net1544 vssd1 vssd1 vccd1 vccd1 net6448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5932 rbzero.tex_b0\[46\] vssd1 vssd1 vccd1 vccd1 net6459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6677 net2387 vssd1 vssd1 vccd1 vccd1 net7204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6688 rbzero.tex_g0\[58\] vssd1 vssd1 vccd1 vccd1 net7215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5943 net1502 vssd1 vssd1 vccd1 vccd1 net6470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6699 net2342 vssd1 vssd1 vccd1 vccd1 net7226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5954 rbzero.spi_registers.new_mapd\[10\] vssd1 vssd1 vccd1 vccd1 net6481 sky130_fd_sc_hd__dlygate4sd3_1
X_21235_ clknet_leaf_14_i_clk _00722_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold240 net6085 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5965 net1538 vssd1 vssd1 vccd1 vccd1 net6492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 net7934 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5976 rbzero.spi_registers.new_texadd\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net6503
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 net4886 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5987 net1223 vssd1 vssd1 vccd1 vccd1 net6514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 net5241 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5998 _04350_ vssd1 vssd1 vccd1 vccd1 net6525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold284 net4556 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
X_21166_ clknet_leaf_131_i_clk net1684 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold295 net8196 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_106_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20117_ _03352_ net5762 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__nor2_1
X_21097_ clknet_leaf_8_i_clk net1458 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ _03483_ _03646_ _03608_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ net3848 _06028_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a21o_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _04821_ _04966_ _04992_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a2bb2o_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21999_ net441 net2341 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _07675_ _07678_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__xnor2_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ net84 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__buf_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ net5546 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__clkbuf_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _07633_ _07640_ _07641_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__a21boi_2
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ net3406 net1361 net3641 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16210_ _09291_ _09302_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13422_ _06459_ _06463_ _06532_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__and3_1
X_10634_ net2994 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__clkbuf_1
X_17190_ _10097_ _10100_ _10209_ vssd1 vssd1 vccd1 vccd1 _10210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_181_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ _08127_ _09116_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13353_ _06435_ _06442_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__or3_1
XFILLER_0_183_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ net6146 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04916_ vssd1 vssd1 vccd1 vccd1 _05490_
+ sky130_fd_sc_hd__mux2_1
X_16072_ _08401_ _09165_ _08180_ _08430_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _06435_ _06442_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__or3_4
X_10496_ net7163 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__clkbuf_1
X_15023_ _08117_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__buf_4
X_19900_ net2934 net3320 _03550_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__mux2_1
X_12235_ _04921_ _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__or2_1
X_19831_ net6661 net1682 _03517_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__mux2_1
X_12166_ _04911_ _05351_ _05353_ _04919_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__o211a_1
X_20465__210 clknet_1_0__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__inv_2
XFILLER_0_120_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11117_ net2930 net6956 _04375_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16974_ _09994_ _09995_ vssd1 vssd1 vccd1 vccd1 _09996_ sky130_fd_sc_hd__nor2_2
X_12097_ _05014_ _05023_ _05285_ _05035_ _05016_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18713_ _02856_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__buf_2
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ net7099 net7346 _04342_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
X_15925_ _09018_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ net1335 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__clkbuf_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _08946_ _08950_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__nand2_1
X_18644_ net4560 rbzero.wall_tracer.rayAddendY\[-1\] vssd1 vssd1 vccd1 vccd1 _02801_
+ sky130_fd_sc_hd__or2_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14807_ net4461 _07968_ _07872_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__mux2_1
X_15787_ _08822_ _08881_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__or2_1
X_18575_ net3965 _09769_ net5918 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ net4518 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__inv_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17526_ _01765_ _01766_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _07860_ _07830_ _07875_ net7843 vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__a211o_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17457_ _01697_ _01698_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14669_ net7842 vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16408_ _09385_ _09386_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17388_ _10404_ _10405_ vssd1 vssd1 vccd1 vccd1 _10406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16339_ _09303_ _09305_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19127_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5206 net5758 vssd1 vssd1 vccd1 vccd1 net5733 sky130_fd_sc_hd__dlygate4sd3_1
X_19058_ net7579 net3481 net3397 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5217 rbzero.pov.ready_buffer\[59\] vssd1 vssd1 vccd1 vccd1 net5744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5228 net4152 vssd1 vssd1 vccd1 vccd1 net5755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5239 net1980 vssd1 vssd1 vccd1 vccd1 net5766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4505 rbzero.wall_tracer.rayAddendX\[-9\] vssd1 vssd1 vccd1 vccd1 net5032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4516 net710 vssd1 vssd1 vccd1 vccd1 net5043 sky130_fd_sc_hd__dlygate4sd3_1
X_18009_ _02238_ _02239_ _02244_ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
Xhold4527 _00784_ vssd1 vssd1 vccd1 vccd1 net5054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4538 net719 vssd1 vssd1 vccd1 vccd1 net5065 sky130_fd_sc_hd__dlygate4sd3_1
X_21020_ clknet_leaf_55_i_clk net4295 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4549 rbzero.spi_registers.texadd1\[8\] vssd1 vssd1 vccd1 vccd1 net5076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3804 net4250 vssd1 vssd1 vccd1 vccd1 net4331 sky130_fd_sc_hd__buf_1
XFILLER_0_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3815 net7905 vssd1 vssd1 vccd1 vccd1 net4342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3826 net7939 vssd1 vssd1 vccd1 vccd1 net4353 sky130_fd_sc_hd__buf_1
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3837 _01187_ vssd1 vssd1 vccd1 vccd1 net4364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3848 _03697_ vssd1 vssd1 vccd1 vccd1 net4375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3859 net2068 vssd1 vssd1 vccd1 vccd1 net4386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21922_ net364 net2597 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21853_ net295 net2684 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20804_ net971 net5726 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21784_ clknet_leaf_0_i_clk net1769 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19790__68 clknet_1_1__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
XFILLER_0_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20735_ _03909_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7120 rbzero.pov.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 net7647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7142 net3807 vssd1 vssd1 vccd1 vccd1 net7669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7153 gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 net7680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7164 rbzero.pov.ready_buffer\[73\] vssd1 vssd1 vccd1 vccd1 net7691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6430 _04383_ vssd1 vssd1 vccd1 vccd1 net6957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7175 _02742_ vssd1 vssd1 vccd1 vccd1 net7702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6441 rbzero.tex_b0\[5\] vssd1 vssd1 vccd1 vccd1 net6968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7186 _09754_ vssd1 vssd1 vccd1 vccd1 net7713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6452 net2339 vssd1 vssd1 vccd1 vccd1 net6979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7197 rbzero.color_sky\[5\] vssd1 vssd1 vccd1 vccd1 net7724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6463 rbzero.tex_g1\[31\] vssd1 vssd1 vccd1 vccd1 net6990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6474 net2970 vssd1 vssd1 vccd1 vccd1 net7001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6485 rbzero.tex_g0\[7\] vssd1 vssd1 vccd1 vccd1 net7012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5740 net1411 vssd1 vssd1 vccd1 vccd1 net6267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5751 _04144_ vssd1 vssd1 vccd1 vccd1 net6278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6496 net2315 vssd1 vssd1 vccd1 vccd1 net7023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5762 net1293 vssd1 vssd1 vccd1 vccd1 net6289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5773 rbzero.spi_registers.new_texadd\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 net6300
+ sky130_fd_sc_hd__dlygate4sd3_1
X_12020_ _05204_ _05205_ _05208_ _04955_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5784 net1323 vssd1 vssd1 vccd1 vccd1 net6311 sky130_fd_sc_hd__dlygate4sd3_1
X_21218_ clknet_leaf_120_i_clk net2942 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5795 _03455_ vssd1 vssd1 vccd1 vccd1 net6322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21149_ clknet_leaf_104_i_clk net4860 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _07098_ _07141_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__xnor2_1
X_15710_ _08749_ _08764_ _08804_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__nand3_1
X_12922_ net3893 _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nor2_1
X_16690_ net8141 _09743_ _09744_ net4280 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _08271_ _08200_ _08252_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__or3b_1
X_12853_ net5605 _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _04836_ vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__mux2_1
X_18360_ _02526_ _02539_ _02540_ _02545_ _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a32o_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _08666_ _08245_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__nand2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12784_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _10321_ _10329_ vssd1 vssd1 vccd1 vccd1 _10330_ sky130_fd_sc_hd__nand2_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _07690_ _07689_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__xor2_1
X_11735_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _04924_ vssd1 vssd1 vccd1 vccd1 _04925_
+ sky130_fd_sc_hd__mux2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ net6307 net3838 _02493_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _10261_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454_ _07583_ _07600_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11666_ _04854_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13405_ _06575_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__clkbuf_4
X_10617_ net2445 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__clkbuf_1
X_17173_ _08309_ _09165_ vssd1 vssd1 vccd1 vccd1 _10193_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14385_ _07512_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11597_ _04783_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16124_ _09204_ _09206_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13336_ _06468_ _06473_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ net2642 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _09139_ _09148_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _06319_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__xnor2_4
X_10479_ net2497 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__clkbuf_1
X_15006_ _08102_ _06159_ _08103_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__a21oi_1
X_12218_ _04921_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__or2_1
X_13198_ _06302_ _06304_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__and2b_1
XFILLER_0_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12149_ _04911_ _05334_ _05336_ _04919_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1709 _04270_ vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_16957_ _09973_ _09977_ _09978_ vssd1 vssd1 vccd1 vccd1 _09979_ sky130_fd_sc_hd__nand3_2
X_15908_ _08211_ _08294_ _08306_ _08207_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_155_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19676_ net1692 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16888_ _09617_ _09909_ vssd1 vssd1 vccd1 vccd1 _09910_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18627_ _02781_ _02784_ _04489_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__a21oi_1
X_15839_ _08893_ _08894_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_17_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18558_ net7671 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _01746_ _01747_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18489_ _02626_ net3614 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__nand2_1
XANTENNA_13 _07903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 net8467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_57 _04921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20437__186 clknet_1_0__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__inv_2
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_68 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5003 rbzero.wall_tracer.mapY\[7\] vssd1 vssd1 vccd1 vccd1 net5530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5014 _03134_ vssd1 vssd1 vccd1 vccd1 net5541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5025 net1530 vssd1 vssd1 vccd1 vccd1 net5552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22121_ clknet_leaf_54_i_clk net5378 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
Xhold5036 _03338_ vssd1 vssd1 vccd1 vccd1 net5563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5047 rbzero.tex_b1\[60\] vssd1 vssd1 vccd1 vccd1 net5574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4302 _00610_ vssd1 vssd1 vccd1 vccd1 net4829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5058 net3874 vssd1 vssd1 vccd1 vccd1 net5585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4313 net3456 vssd1 vssd1 vccd1 vccd1 net4840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5069 net1822 vssd1 vssd1 vccd1 vccd1 net5596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4324 rbzero.wall_tracer.rayAddendX\[-6\] vssd1 vssd1 vccd1 vccd1 net4851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4335 net3627 vssd1 vssd1 vccd1 vccd1 net4862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4346 net3944 vssd1 vssd1 vccd1 vccd1 net4873 sky130_fd_sc_hd__dlygate4sd3_1
X_22052_ net494 net2338 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold3601 _05680_ vssd1 vssd1 vccd1 vccd1 net4128 sky130_fd_sc_hd__clkbuf_4
Xhold3612 _04669_ vssd1 vssd1 vccd1 vccd1 net4139 sky130_fd_sc_hd__clkbuf_2
Xhold4357 _00596_ vssd1 vssd1 vccd1 vccd1 net4884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3623 _08095_ vssd1 vssd1 vccd1 vccd1 net4150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4368 net8402 vssd1 vssd1 vccd1 vccd1 net4895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3634 _05042_ vssd1 vssd1 vccd1 vccd1 net4161 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold4379 net3767 vssd1 vssd1 vccd1 vccd1 net4906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2900 net7938 vssd1 vssd1 vccd1 vccd1 net3427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3645 _05175_ vssd1 vssd1 vccd1 vccd1 net4172 sky130_fd_sc_hd__dlygate4sd3_1
X_21003_ clknet_leaf_85_i_clk _00490_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2911 _01201_ vssd1 vssd1 vccd1 vccd1 net3438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3656 _08111_ vssd1 vssd1 vccd1 vccd1 net4183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2922 _00617_ vssd1 vssd1 vccd1 vccd1 net3449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3667 net8298 vssd1 vssd1 vccd1 vccd1 net4194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3678 net7890 vssd1 vssd1 vccd1 vccd1 net4205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2933 net7870 vssd1 vssd1 vccd1 vccd1 net3460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3689 net8301 vssd1 vssd1 vccd1 vccd1 net4216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2944 _01196_ vssd1 vssd1 vccd1 vccd1 net3471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2955 net7580 vssd1 vssd1 vccd1 vccd1 net3482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2966 rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 net3493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2977 net7626 vssd1 vssd1 vccd1 vccd1 net3504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2988 net4786 vssd1 vssd1 vccd1 vccd1 net3515 sky130_fd_sc_hd__dlygate4sd3_1
X_20602__334 clknet_1_1__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__inv_2
X_21905_ net347 net2577 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21836_ net278 net999 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21767_ clknet_leaf_15_i_clk net1342 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11520_ _04670_ net4324 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand2_1
X_20718_ net5380 _03877_ _03874_ _03898_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21698_ clknet_leaf_116_i_clk net5753 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _04566_ _04555_ rbzero.spi_registers.texadd3\[1\] vssd1 vssd1 vccd1 vccd1
+ _04643_ sky130_fd_sc_hd__or3b_1
XFILLER_0_110_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20649_ clknet_1_0__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__buf_1
XFILLER_0_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14170_ _07339_ _07340_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ rbzero.spi_registers.texadd2\[22\] _04567_ _04548_ rbzero.spi_registers.texadd1\[22\]
+ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6260 rbzero.tex_b0\[45\] vssd1 vssd1 vccd1 vccd1 net6787 sky130_fd_sc_hd__dlygate4sd3_1
X_13121_ _06284_ _06288_ _06291_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__and3_1
Xhold6271 net2050 vssd1 vssd1 vccd1 vccd1 net6798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6282 _04225_ vssd1 vssd1 vccd1 vccd1 net6809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6293 net2227 vssd1 vssd1 vccd1 vccd1 net6820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5570 _04426_ vssd1 vssd1 vccd1 vccd1 net6097 sky130_fd_sc_hd__dlygate4sd3_1
X_13052_ _06210_ _06227_ _06219_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__o21ai_1
Xhold5581 _04294_ vssd1 vssd1 vccd1 vccd1 net6108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5592 _04338_ vssd1 vssd1 vccd1 vccd1 net6119 sky130_fd_sc_hd__dlygate4sd3_1
X_12003_ net4177 _05191_ _04460_ _04601_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__or4b_1
XFILLER_0_178_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4880 rbzero.wall_tracer.mapY\[10\] vssd1 vssd1 vccd1 vccd1 net5407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17860_ _02033_ _02013_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__or2b_1
Xhold4891 net1005 vssd1 vssd1 vccd1 vccd1 net5418 sky130_fd_sc_hd__dlygate4sd3_1
X_16811_ _09838_ net4547 net4649 vssd1 vssd1 vccd1 vccd1 _09839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17791_ _02021_ _02029_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19530_ net3087 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
X_16742_ _09775_ _09776_ _09773_ vssd1 vssd1 vccd1 vccd1 _09778_ sky130_fd_sc_hd__o21ai_1
X_13954_ _06857_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12905_ net3959 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__inv_2
X_20577__311 clknet_1_0__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__inv_2
X_19461_ net3486 net3906 _02947_ _02969_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__and4bb_1
X_16673_ _09739_ vssd1 vssd1 vccd1 vccd1 _09742_ sky130_fd_sc_hd__buf_4
X_13885_ _07016_ _07055_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18412_ _02593_ _02594_ rbzero.wall_tracer.rayAddendX\[1\] _09736_ vssd1 vssd1 vccd1
+ vccd1 _02595_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15624_ _08716_ _08717_ _08718_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__nand3_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _06007_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__or2_1
XFILLER_0_201_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ net5272 _03268_ _03298_ _03299_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__o211a_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ _08625_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__xor2_1
X_18343_ net3509 net5961 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__nand2_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ net39 _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__nand2_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _07489_ _07194_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11718_ net5356 net7730 _04845_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux2_1
X_18274_ net6291 net1426 _02477_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
X_15486_ _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ _05850_ net30 net31 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a21o_1
X_17225_ _10243_ _10244_ vssd1 vssd1 vccd1 vccd1 _10245_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14437_ _07556_ _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ net1209 _04828_ _04832_ net1136 vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a22o_1
Xinput11 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__03863_ clknet_0__03863_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03863_
+ sky130_fd_sc_hd__clkbuf_16
Xinput22 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_2
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput33 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_2
XFILLER_0_142_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17156_ _10173_ _10174_ vssd1 vssd1 vccd1 vccd1 _10176_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_6
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput55 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_8
X_14368_ _06924_ _07304_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__nor2_1
Xhold806 _00986_ vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _09199_ _09200_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__nor2_1
Xhold817 net6192 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13319_ net82 _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nor2_1
Xhold828 net6371 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ _09979_ _09981_ _10107_ vssd1 vssd1 vccd1 vccd1 _10108_ sky130_fd_sc_hd__a21oi_1
Xhold839 _03340_ vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14299_ _07464_ _07467_ _07468_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16038_ _09023_ _09016_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__or2b_1
XFILLER_0_110_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2207 rbzero.tex_b1\[47\] vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2218 _04424_ vssd1 vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 _04136_ vssd1 vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1506 _04153_ vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 _04132_ vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
X_17989_ _02130_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__or3b_1
Xhold1528 net6791 vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 net7474 vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
X_19728_ net5496 _03489_ _03495_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__o21a_1
XFILLER_0_205_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20443__190 clknet_1_1__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__inv_2
X_19659_ net6321 net3631 _03429_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21621_ clknet_leaf_128_i_clk net2922 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21552_ net186 net2919 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21483_ clknet_leaf_44_i_clk net1546 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20673__18 clknet_1_1__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XFILLER_0_105_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4110 _01232_ vssd1 vssd1 vccd1 vccd1 net4637 sky130_fd_sc_hd__dlygate4sd3_1
X_22104_ net166 net2299 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold4121 _09767_ vssd1 vssd1 vccd1 vccd1 net4648 sky130_fd_sc_hd__buf_4
Xhold4132 net3861 vssd1 vssd1 vccd1 vccd1 net4659 sky130_fd_sc_hd__clkbuf_2
X_20296_ net6283 net3863 _03814_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4154 net3379 vssd1 vssd1 vccd1 vccd1 net4681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3420 _02652_ vssd1 vssd1 vccd1 vccd1 net3947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4165 _00426_ vssd1 vssd1 vccd1 vccd1 net4692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3431 _00474_ vssd1 vssd1 vccd1 vccd1 net3958 sky130_fd_sc_hd__dlygate4sd3_1
X_22035_ net477 net2249 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4176 net7805 vssd1 vssd1 vccd1 vccd1 net4703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4187 _02513_ vssd1 vssd1 vccd1 vccd1 net4714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3442 net6000 vssd1 vssd1 vccd1 vccd1 net3969 sky130_fd_sc_hd__buf_1
Xhold4198 _02581_ vssd1 vssd1 vccd1 vccd1 net4725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3453 _03396_ vssd1 vssd1 vccd1 vccd1 net3980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3464 _04678_ vssd1 vssd1 vccd1 vccd1 net3991 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2730 _03553_ vssd1 vssd1 vccd1 vccd1 net3257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3475 rbzero.debug_overlay.facingY\[10\] vssd1 vssd1 vccd1 vccd1 net4002 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2741 _00712_ vssd1 vssd1 vccd1 vccd1 net3268 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3486 _08110_ vssd1 vssd1 vccd1 vccd1 net4013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2752 net5867 vssd1 vssd1 vccd1 vccd1 net3279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3497 net5982 vssd1 vssd1 vccd1 vccd1 net4024 sky130_fd_sc_hd__buf_4
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2763 _03020_ vssd1 vssd1 vccd1 vccd1 net3290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2774 rbzero.pov.spi_buffer\[30\] vssd1 vssd1 vccd1 vccd1 net3301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2785 net3223 vssd1 vssd1 vccd1 vccd1 net3312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2796 net5770 vssd1 vssd1 vccd1 vccd1 net3323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ net6936 net6591 _04287_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13670_ _06795_ _06839_ _06818_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__a31oi_2
X_10882_ net2053 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _05796_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__and3_1
Xwire90 _09787_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21819_ net261 net2825 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15340_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _08435_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_54_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ net4102 net4024 net10 vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ net5981 net3445 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__xnor2_1
X_15271_ net4496 _08133_ _08362_ _08365_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__a22o_4
X_12483_ _05203_ _05643_ _05644_ net41 vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17010_ _09603_ _10030_ vssd1 vssd1 vccd1 vccd1 _10031_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14222_ _07388_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _04528_ _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ _07143_ _07146_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11365_ rbzero.spi_registers.texadd3\[16\] rbzero.spi_registers.texadd1\[16\] rbzero.spi_registers.texadd0\[16\]
+ rbzero.spi_registers.texadd2\[16\] _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04557_
+ sky130_fd_sc_hd__mux4_2
Xhold6090 net1487 vssd1 vssd1 vccd1 vccd1 net6617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14084_ _07204_ _07249_ _07253_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__and3_1
X_18961_ net5710 net4327 net2874 vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
X_11296_ net8051 _04483_ _04488_ _04490_ _04486_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _02148_ _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__and2_1
X_13035_ _06204_ _06206_ _06208_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__or4_1
X_18892_ net1753 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
X_17843_ _10327_ _08799_ _01693_ _09976_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__or4_1
XFILLER_0_195_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17774_ _01902_ _01912_ _01910_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14986_ net4622 _08032_ _08067_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__mux2_1
X_19513_ _04102_ net3084 _03344_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16725_ net4049 net3884 _09103_ vssd1 vssd1 vccd1 vccd1 _09763_ sky130_fd_sc_hd__o21a_1
X_13937_ _06771_ _06829_ _06830_ _06833_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19444_ net4956 _03323_ _03332_ _03316_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__a211o_1
X_13868_ _06703_ _06832_ _07038_ _07036_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16656_ _04479_ _09734_ vssd1 vssd1 vccd1 vccd1 _09735_ sky130_fd_sc_hd__and2_2
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ _08658_ _08689_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12819_ _05992_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__nor2_1
X_19375_ net5101 _03283_ _03290_ _03288_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__o211a_1
X_16587_ _09676_ _09546_ _08474_ vssd1 vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__a21oi_1
X_13799_ net80 net79 vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__or2_1
XFILLER_0_201_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18326_ _02511_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15538_ _08372_ _08373_ net8033 net4877 _08383_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__o32ai_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7708 rbzero.debug_overlay.playerY\[2\] vssd1 vssd1 vccd1 vccd1 net8235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7719 _02938_ vssd1 vssd1 vccd1 vccd1 net8246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15469_ _08521_ _08563_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18257_ net3897 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17208_ _10101_ _10106_ _10105_ vssd1 vssd1 vccd1 vccd1 _10228_ sky130_fd_sc_hd__a21bo_1
X_20631__360 clknet_1_1__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__inv_2
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03846_ clknet_0__03846_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03846_
+ sky130_fd_sc_hd__clkbuf_16
X_18188_ _02407_ _02408_ _02401_ _02409_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 net6196 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17139_ _10157_ _10158_ vssd1 vssd1 vccd1 vccd1 _10159_ sky130_fd_sc_hd__nor2_1
Xhold614 _01379_ vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold625 _03560_ vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold636 net5467 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 net6212 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 net6218 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ net7083 _03707_ net4447 _03679_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 _00659_ vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20081_ _08288_ _03610_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__nor2_1
Xhold2004 _04111_ vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 net3051 vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2026 _01448_ vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 net6855 vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2048 net7290 vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1303 net7521 vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 _01552_ vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2059 _00687_ vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 net5564 vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1336 _02997_ vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1347 _01354_ vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1358 net6743 vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 _01514_ vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ clknet_leaf_58_i_clk _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_205_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21604_ clknet_leaf_131_i_clk net1318 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21535_ net169 net1838 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21466_ clknet_leaf_42_i_clk net2005 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21397_ clknet_leaf_39_i_clk net5511 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11150_ net6995 net2387 _04390_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ _04193_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20279_ net5966 net4099 _03811_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__o21a_1
Xhold3250 net3665 vssd1 vssd1 vccd1 vccd1 net3777 sky130_fd_sc_hd__clkbuf_2
X_22018_ net460 net2757 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold3261 net8416 vssd1 vssd1 vccd1 vccd1 net3788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3272 _09869_ vssd1 vssd1 vccd1 vccd1 net3799 sky130_fd_sc_hd__buf_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3283 net7989 vssd1 vssd1 vccd1 vccd1 net3810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3294 net7872 vssd1 vssd1 vccd1 vccd1 net3821 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2560 _03382_ vssd1 vssd1 vccd1 vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2571 net5744 vssd1 vssd1 vccd1 vccd1 net3098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14840_ net7794 _07937_ _07997_ net4704 vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__a211o_2
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2582 _01372_ vssd1 vssd1 vccd1 vccd1 net3109 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2593 rbzero.pov.spi_buffer\[54\] vssd1 vssd1 vccd1 vccd1 net3120 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03866_ clknet_0__03866_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03866_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1870 _03681_ vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1881 rbzero.tex_g1\[32\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ _07934_ _07936_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__and2_2
X_11983_ _05130_ _05171_ _04659_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a21bo_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1892 _01459_ vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_16510_ _09116_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13722_ _06891_ _06892_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__nor2_1
X_10934_ _04264_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__clkbuf_4
X_17490_ _01731_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16441_ _09530_ _09531_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _06751_ _06750_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__and2b_1
X_10865_ net2827 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ net52 _05744_ _05763_ net53 vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__a22o_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _09369_ _09340_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__or2b_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19160_ net1429 _03146_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__or2_1
X_13584_ _06618_ _06634_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__xnor2_4
X_10796_ net2971 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _08376_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__buf_2
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _02342_ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__clkbuf_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12535_ net55 _05700_ _05701_ net52 vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091_ net4092 net4138 _04657_ net4127 vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ _08340_ _08347_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__nor2_1
X_18042_ _02274_ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__xnor2_1
X_12466_ _04102_ _05642_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a21o_2
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14205_ _07358_ _07357_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11417_ _04496_ _04591_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__or3b_1
XFILLER_0_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15185_ _08279_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__clkbuf_4
X_12397_ _04991_ _05556_ _05564_ _04849_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a311o_1
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14136_ _07306_ _07303_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__nor2_2
X_11348_ _04517_ _04537_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a21o_1
X_19993_ net4168 _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__nor2_1
X_18944_ net3260 net7093 _03036_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
X_14067_ _07199_ _07236_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__nand2_1
X_11279_ net3975 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__buf_1
XFILLER_0_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13018_ net3875 vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__inv_2
X_18875_ net3145 net7508 _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ _02062_ _02063_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _01981_ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__xnor2_1
X_14969_ _08082_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__clkbuf_1
X_16708_ _04567_ net7665 _09747_ vssd1 vssd1 vccd1 vccd1 _09748_ sky130_fd_sc_hd__mux2_1
X_17688_ _01815_ _01819_ _01926_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ _03320_ net3652 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__and2_1
X_16639_ net7679 net3956 _09725_ vssd1 vssd1 vccd1 vccd1 _09726_ sky130_fd_sc_hd__and3b_1
XFILLER_0_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19358_ net5312 _03269_ _03280_ _03275_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18309_ net6426 net1447 _02493_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20555__291 clknet_1_0__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__inv_2
XFILLER_0_45_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19289_ net1422 _03238_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__or2_1
Xhold7538 net8420 vssd1 vssd1 vccd1 vccd1 net8065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6804 rbzero.tex_b0\[16\] vssd1 vssd1 vccd1 vccd1 net7331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7549 _02586_ vssd1 vssd1 vccd1 vccd1 net8076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6815 net2930 vssd1 vssd1 vccd1 vccd1 net7342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21320_ clknet_leaf_13_i_clk net5266 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6826 net2596 vssd1 vssd1 vccd1 vccd1 net7353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6837 rbzero.tex_r1\[53\] vssd1 vssd1 vccd1 vccd1 net7364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6848 net2895 vssd1 vssd1 vccd1 vccd1 net7375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6859 rbzero.tex_b0\[18\] vssd1 vssd1 vccd1 vccd1 net7386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21251_ clknet_leaf_0_i_clk net3558 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold400 net5219 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 net6102 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 net4300 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold433 net8125 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
X_20202_ _04459_ net3495 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__or2_1
Xhold444 net8221 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_1
X_21182_ clknet_leaf_128_i_clk net3184 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold455 net5271 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 net5287 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 net5415 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 net8228 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
X_20133_ _03689_ net7660 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__or2_1
Xhold499 net3361 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
X_20064_ _03661_ net4617 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__or2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _00914_ vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 net6575 vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 net6618 vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1133 net6698 vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 net6577 vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 net7309 vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1166 _00996_ vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 _03067_ vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 net6640 vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 _00907_ vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20966_ clknet_leaf_70_i_clk _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20897_ clknet_leaf_84_i_clk net5781 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_166_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10650_ net6737 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10581_ net5550 net1529 _04097_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _04911_ _05503_ _05505_ _04919_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21518_ clknet_leaf_7_i_clk net1498 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _04968_ vssd1 vssd1 vccd1 vccd1 _05438_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21449_ clknet_leaf_39_i_clk net1624 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ net6832 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12182_ _05213_ _04949_ _05369_ _05025_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11133_ net2361 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__clkbuf_1
X_16990_ _10011_ net4669 net4649 vssd1 vssd1 vccd1 vccd1 _10012_ sky130_fd_sc_hd__mux2_1
X_11064_ net2633 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
X_15941_ net8041 _06121_ _08491_ _09035_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__or4_4
Xhold3091 rbzero.debug_overlay.vplaneY\[-5\] vssd1 vssd1 vccd1 vccd1 net3618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18660_ _02814_ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__nand2_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _08957_ _08963_ _08965_ _08966_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__o2bb2a_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2390 net7386 vssd1 vssd1 vccd1 vccd1 net2917 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17611_ _01849_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__nor2_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _07982_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
X_19796__74 clknet_1_0__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ net4635 net4879 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03849_ clknet_0__03849_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03849_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _10062_ _09040_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11966_ net4713 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__clkbuf_4
X_14754_ net7850 _07846_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__nor2_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10917_ net2605 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
X_13705_ _06874_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__xnor2_1
X_17473_ _10367_ _10369_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__nor2_1
X_14685_ _07818_ _07853_ _07855_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__a21oi_1
X_11897_ _05066_ net3517 _05075_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19212_ net5220 _03182_ _03194_ _03189_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__o211a_1
X_16424_ _09513_ _09514_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__nor2_1
X_13636_ _06805_ _06806_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__nor2_1
X_10848_ net2595 net6223 _04238_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19143_ net5613 _03147_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__or2_1
X_16355_ _09218_ _09317_ _09315_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__a21oi_4
X_13567_ _06683_ _06737_ net79 vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__a21oi_1
X_10779_ net2429 net6114 _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15306_ _08161_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__buf_2
X_12518_ net11 _05691_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__and2b_1
X_16286_ _08226_ _08535_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19074_ net44 net6611 _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13498_ _06478_ _06467_ _06571_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18025_ _02191_ _02215_ _02217_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15237_ _08331_ _08327_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__xnor2_1
X_12449_ reg_hsync _05631_ _05054_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__mux2_2
XFILLER_0_23_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4709 net936 vssd1 vssd1 vccd1 vccd1 net5236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ _08261_ _08262_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14119_ _07288_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19976_ net1809 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
X_15099_ _08156_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__buf_4
XFILLER_0_201_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18927_ net3273 net7595 _03025_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18858_ net3351 net4825 _02993_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17809_ _01962_ _01963_ _02046_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18789_ net8243 _02921_ _02919_ net8242 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20820_ net850 net5609 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20751_ _03919_ _03920_ _03921_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_187_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8014 rbzero.debug_overlay.playerY\[-8\] vssd1 vssd1 vccd1 vccd1 net8541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7313 rbzero.wall_tracer.trackDistY\[-11\] vssd1 vssd1 vccd1 vccd1 net7840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7324 rbzero.wall_tracer.stepDistY\[-5\] vssd1 vssd1 vccd1 vccd1 net7851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7335 net4191 vssd1 vssd1 vccd1 vccd1 net7862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6601 rbzero.tex_r0\[21\] vssd1 vssd1 vccd1 vccd1 net7128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7346 net3821 vssd1 vssd1 vccd1 vccd1 net7873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7357 rbzero.traced_texVinit\[2\] vssd1 vssd1 vccd1 vccd1 net7884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6612 net2377 vssd1 vssd1 vccd1 vccd1 net7139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7368 net1086 vssd1 vssd1 vccd1 vccd1 net7895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6623 _04151_ vssd1 vssd1 vccd1 vccd1 net7150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6634 net2011 vssd1 vssd1 vccd1 vccd1 net7161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5900 _02503_ vssd1 vssd1 vccd1 vccd1 net6427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7379 net4342 vssd1 vssd1 vccd1 vccd1 net7906 sky130_fd_sc_hd__dlygate4sd3_1
X_21303_ clknet_leaf_48_i_clk net5258 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6645 _04223_ vssd1 vssd1 vccd1 vccd1 net7172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6656 rbzero.tex_r0\[50\] vssd1 vssd1 vccd1 vccd1 net7183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5911 net1245 vssd1 vssd1 vccd1 vccd1 net6438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6667 net2491 vssd1 vssd1 vccd1 vccd1 net7194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5922 rbzero.spi_registers.new_texadd\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net6449
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5933 net1197 vssd1 vssd1 vccd1 vccd1 net6460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6678 _04402_ vssd1 vssd1 vccd1 vccd1 net7205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6689 net2685 vssd1 vssd1 vccd1 vccd1 net7216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5944 rbzero.spi_registers.new_texadd\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net6471
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 net7913 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5955 net1289 vssd1 vssd1 vccd1 vccd1 net6482 sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ clknet_leaf_15_i_clk net3901 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold241 _01493_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold252 net7092 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5966 rbzero.spi_registers.new_other\[2\] vssd1 vssd1 vccd1 vccd1 net6493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5977 net1694 vssd1 vssd1 vccd1 vccd1 net6504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 net4888 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5988 rbzero.spi_registers.new_texadd\[0\]\[19\] vssd1 vssd1 vccd1 vccd1 net6515
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5999 net1409 vssd1 vssd1 vccd1 vccd1 net6526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 net5267 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
X_21165_ clknet_leaf_132_i_clk net1972 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold285 net5168 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold296 net8023 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
X_20116_ net3469 _03699_ net5760 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a21oi_1
X_21096_ clknet_leaf_11_i_clk net1861 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20047_ net7605 _03631_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nor2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _04818_ _05009_ _04821_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__o21a_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ net440 net2730 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _04825_ _04920_ _04929_ _04940_ _04844_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__o311a_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20949_ clknet_leaf_64_i_clk _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ net5544 net2122 _04160_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14470_ _07634_ _07635_ _07639_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__nand3_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20571__306 clknet_1_1__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__inv_2
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ net3406 net3641 net3857 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _06498_ _06571_ _06591_ _06492_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__a211o_1
X_10633_ net7441 net6669 _04127_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16140_ _09231_ _09232_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _06522_ _06447_ _06450_ _06453_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__or4_1
X_10564_ net2370 net6144 _04086_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux2_1
X_12303_ _04911_ _05486_ _05488_ _04928_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16071_ _09031_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__buf_2
XFILLER_0_162_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13283_ _06445_ _06447_ _06450_ _06453_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__or4_2
X_10495_ net2657 net7161 _04053_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__mux2_1
Xhold7891 _08249_ vssd1 vssd1 vccd1 vccd1 net8418 sky130_fd_sc_hd__dlygate4sd3_1
X_15022_ _08116_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__buf_4
X_12234_ rbzero.tex_g1\[39\] rbzero.tex_g1\[38\] _04837_ vssd1 vssd1 vccd1 vccd1 _05421_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19830_ net6415 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
X_12165_ _04915_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__or2_1
X_11116_ net6054 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
X_16973_ _09991_ _09993_ vssd1 vssd1 vccd1 vccd1 _09995_ sky130_fd_sc_hd__and2_1
X_12096_ net4080 _05032_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18712_ _02856_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _02864_
+ sky130_fd_sc_hd__xor2_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net2334 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
X_15924_ _08392_ _08391_ _08244_ _08386_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__a2bb2o_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_102_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19692_ net6472 net3738 _03468_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_4
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ net4560 rbzero.wall_tracer.rayAddendY\[-1\] vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__nand2_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _08947_ _08949_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _07964_ _07931_ _07967_ net7823 net3638 vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__a221o_4
X_18574_ _09769_ net5917 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nor2_1
X_15786_ _08880_ _08329_ _08691_ _08391_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__o22a_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ net4667 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__inv_2
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _10190_ _09116_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14737_ _07860_ _07804_ _07884_ net7811 vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__a211o_1
XFILLER_0_197_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11949_ rbzero.debug_overlay.facingX\[-9\] _05106_ net4161 gpout0.vpos\[5\] vssd1
+ vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a211o_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17456_ _10105_ _01692_ _01696_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14668_ net7807 _07837_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__and3_4
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _09465_ _09497_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__xnor2_4
X_13619_ _06787_ _06776_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__or2b_1
X_17387_ _08864_ _10289_ vssd1 vssd1 vccd1 vccd1 _10405_ sky130_fd_sc_hd__nor2_1
X_14599_ _07762_ _07765_ _07737_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__a21oi_1
X_19126_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__clkbuf_2
X_16338_ _09401_ _09429_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19057_ net3479 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__clkbuf_1
Xhold5207 _03057_ vssd1 vssd1 vccd1 vccd1 net5734 sky130_fd_sc_hd__dlygate4sd3_1
X_16269_ _09251_ _09256_ _09359_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5218 net3098 vssd1 vssd1 vccd1 vccd1 net5745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5229 _00756_ vssd1 vssd1 vccd1 vccd1 net5756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ net89 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__clkbuf_8
Xhold4506 net666 vssd1 vssd1 vccd1 vccd1 net5033 sky130_fd_sc_hd__buf_1
XFILLER_0_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4517 rbzero.pov.ready_buffer\[10\] vssd1 vssd1 vccd1 vccd1 net5044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4528 net714 vssd1 vssd1 vccd1 vccd1 net5055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4539 _00799_ vssd1 vssd1 vccd1 vccd1 net5066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3805 _08065_ vssd1 vssd1 vccd1 vccd1 net4332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3816 net7907 vssd1 vssd1 vccd1 vccd1 net4343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3827 net8166 vssd1 vssd1 vccd1 vccd1 net4354 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3838 net3318 vssd1 vssd1 vccd1 vccd1 net4365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3849 _01194_ vssd1 vssd1 vccd1 vccd1 net4376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19959_ net5812 net3009 _03583_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21921_ net363 net2464 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21852_ net294 net1300 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19775__55 clknet_1_0__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XFILLER_0_210_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20803_ net971 net5726 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__nor2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21783_ clknet_leaf_0_i_clk net1578 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20734_ _03910_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7110 _02722_ vssd1 vssd1 vccd1 vccd1 net7637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7121 net3921 vssd1 vssd1 vccd1 vccd1 net7648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7132 _03716_ vssd1 vssd1 vccd1 vccd1 net7659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7143 _02726_ vssd1 vssd1 vccd1 vccd1 net7670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7154 net4110 vssd1 vssd1 vccd1 vccd1 net7681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6420 rbzero.tex_b1\[23\] vssd1 vssd1 vccd1 vccd1 net6947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7165 _03657_ vssd1 vssd1 vccd1 vccd1 net7692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6431 net2150 vssd1 vssd1 vccd1 vccd1 net6958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7176 _02743_ vssd1 vssd1 vccd1 vccd1 net7703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6442 net1943 vssd1 vssd1 vccd1 vccd1 net6969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7187 _02735_ vssd1 vssd1 vccd1 vccd1 net7714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6453 _04157_ vssd1 vssd1 vccd1 vccd1 net6980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7198 net3651 vssd1 vssd1 vccd1 vccd1 net7725 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20414__165 clknet_1_0__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__inv_2
Xhold6464 net2566 vssd1 vssd1 vccd1 vccd1 net6991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6475 rbzero.pov.ready_buffer\[5\] vssd1 vssd1 vccd1 vccd1 net7002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5730 net1200 vssd1 vssd1 vccd1 vccd1 net6257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6486 net2354 vssd1 vssd1 vccd1 vccd1 net7013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5741 _04387_ vssd1 vssd1 vccd1 vccd1 net6268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6497 rbzero.tex_b0\[39\] vssd1 vssd1 vccd1 vccd1 net7024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5752 net1207 vssd1 vssd1 vccd1 vccd1 net6279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5763 rbzero.spi_registers.new_texadd\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net6290
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5774 net1328 vssd1 vssd1 vccd1 vccd1 net6301 sky130_fd_sc_hd__dlygate4sd3_1
X_21217_ clknet_leaf_120_i_clk net3040 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5785 rbzero.spi_registers.new_texadd\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net6312
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5796 net1267 vssd1 vssd1 vccd1 vccd1 net6323 sky130_fd_sc_hd__dlygate4sd3_1
X_21148_ clknet_leaf_103_i_clk net3743 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_21079_ clknet_leaf_71_i_clk _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13970_ _07137_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _06039_ net3848 net4044 net3807 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15640_ _08729_ _08731_ _08734_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__nand3_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12852_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__clkbuf_4
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _04979_ vssd1 vssd1 vccd1 vccd1 _04993_
+ sky130_fd_sc_hd__mux2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _05957_ _05958_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _08199_ _08195_ net8425 _08192_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__o2bb2a_4
X_20495__237 clknet_1_1__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__inv_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17310_ _10326_ _10328_ vssd1 vssd1 vccd1 vccd1 _10329_ sky130_fd_sc_hd__xor2_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_139_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _07656_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__and2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _02476_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17241_ _10259_ net4657 _10260_ vssd1 vssd1 vccd1 vccd1 _10261_ sky130_fd_sc_hd__mux2_1
X_20679__24 clknet_1_0__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
X_14453_ _07622_ _07623_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__nor2b_1
X_11665_ net3406 net1361 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10616_ net7200 net7184 _04116_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13404_ net73 _06544_ _06546_ _06556_ _06574_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a221oi_4
X_17172_ _10189_ _10191_ vssd1 vssd1 vccd1 vccd1 _10192_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14384_ _07531_ _07553_ _07554_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a21oi_1
X_11596_ net2474 _04784_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_148_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ _06472_ _06441_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__nor2_1
X_16123_ _08115_ _09214_ _09215_ net4613 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_150_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10547_ net6872 net7055 _04075_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16054_ _09146_ _09147_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__nor2_1
X_13266_ _06404_ _06354_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nand2_2
X_10478_ net6140 net6952 _04042_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20389__142 clknet_1_1__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__inv_2
X_12217_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _04933_ vssd1 vssd1 vccd1 vccd1 _05404_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15005_ net4865 vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__buf_6
X_13197_ _06268_ _06269_ _06300_ _06301_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__a31o_2
XFILLER_0_208_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ _04938_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or2_1
X_19744_ clknet_1_0__leaf__03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__buf_1
X_12079_ _05266_ _05267_ _05206_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__mux2_1
X_16956_ _09674_ _09677_ _09675_ vssd1 vssd1 vccd1 vccd1 _09978_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15907_ _08211_ _08207_ _08294_ _08305_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__or4_1
X_19675_ net6599 net3863 _03457_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16887_ _08204_ _09354_ vssd1 vssd1 vccd1 vccd1 _09909_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18626_ _02781_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15838_ _08859_ _08895_ _08932_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__and3_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18557_ _02725_ net7669 _06242_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
X_15769_ _08129_ _08223_ _08224_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__a21o_4
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17508_ _10395_ _01748_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__nor2_1
X_18488_ net5892 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17439_ _10340_ _10342_ _10339_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_145_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 _08295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_36 net3469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_47 _03202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 _04942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20450_ clknet_1_0__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_69 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19109_ net5526 _03126_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__05847_ _05847_ vssd1 vssd1 vccd1 vccd1 clknet_0__05847_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5004 net1611 vssd1 vssd1 vccd1 vccd1 net5531 sky130_fd_sc_hd__buf_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5015 _00762_ vssd1 vssd1 vccd1 vccd1 net5542 sky130_fd_sc_hd__dlygate4sd3_1
X_22120_ clknet_leaf_55_i_clk net5342 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
Xhold5026 rbzero.wall_tracer.mapX\[6\] vssd1 vssd1 vccd1 vccd1 net5553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5037 _00899_ vssd1 vssd1 vccd1 vccd1 net5564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5048 _04323_ vssd1 vssd1 vccd1 vccd1 net5575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4303 net3530 vssd1 vssd1 vccd1 vccd1 net4830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4314 rbzero.spi_registers.got_new_texadd\[2\] vssd1 vssd1 vccd1 vccd1 net4841
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5059 rbzero.tex_b1\[14\] vssd1 vssd1 vccd1 vccd1 net5586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4325 net781 vssd1 vssd1 vccd1 vccd1 net4852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22051_ net493 net2326 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold4336 _04475_ vssd1 vssd1 vccd1 vccd1 net4863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4347 rbzero.wall_tracer.trackDistY\[-9\] vssd1 vssd1 vccd1 vccd1 net4874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3602 _03802_ vssd1 vssd1 vccd1 vccd1 net4129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4358 net918 vssd1 vssd1 vccd1 vccd1 net4885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3613 _05174_ vssd1 vssd1 vccd1 vccd1 net4140 sky130_fd_sc_hd__buf_1
Xhold4369 rbzero.wall_tracer.trackDistY\[4\] vssd1 vssd1 vccd1 vccd1 net4896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3624 _00459_ vssd1 vssd1 vccd1 vccd1 net4151 sky130_fd_sc_hd__dlygate4sd3_1
X_21002_ clknet_leaf_85_i_clk _00489_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3635 _05046_ vssd1 vssd1 vccd1 vccd1 net4162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3646 _05628_ vssd1 vssd1 vccd1 vccd1 net4173 sky130_fd_sc_hd__buf_2
Xhold2901 net4899 vssd1 vssd1 vccd1 vccd1 net3428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2912 rbzero.pov.ready_buffer\[44\] vssd1 vssd1 vccd1 vccd1 net3439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3657 _00465_ vssd1 vssd1 vccd1 vccd1 net4184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3668 net8115 vssd1 vssd1 vccd1 vccd1 net4195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2923 net7852 vssd1 vssd1 vccd1 vccd1 net3450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3679 net7892 vssd1 vssd1 vccd1 vccd1 net4206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2934 net7770 vssd1 vssd1 vccd1 vccd1 net3461 sky130_fd_sc_hd__buf_2
Xhold2945 net7941 vssd1 vssd1 vccd1 vccd1 net3472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2956 _00742_ vssd1 vssd1 vccd1 vccd1 net3483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2967 _02552_ vssd1 vssd1 vccd1 vccd1 net3494 sky130_fd_sc_hd__clkbuf_4
Xhold2978 _03734_ vssd1 vssd1 vccd1 vccd1 net3505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2989 net5204 vssd1 vssd1 vccd1 vccd1 net3516 sky130_fd_sc_hd__buf_1
XFILLER_0_173_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21904_ net346 net2016 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21835_ net277 net2002 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21766_ clknet_leaf_83_i_clk net3997 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20717_ _03894_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__xnor2_1
X_21697_ clknet_leaf_115_i_clk net5861 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ rbzero.spi_registers.texadd2\[1\] _04566_ _04567_ _04020_ vssd1 vssd1 vccd1
+ vccd1 _04642_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11381_ rbzero.spi_registers.texadd3\[22\] _04567_ _04554_ vssd1 vssd1 vccd1 vccd1
+ _04573_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6250 _04300_ vssd1 vssd1 vccd1 vccd1 net6777 sky130_fd_sc_hd__dlygate4sd3_1
X_13120_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6261 net1982 vssd1 vssd1 vccd1 vccd1 net6788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6272 rbzero.spi_registers.new_mapd\[1\] vssd1 vssd1 vccd1 vccd1 net6799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6283 net1962 vssd1 vssd1 vccd1 vccd1 net6810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6294 rbzero.tex_r0\[39\] vssd1 vssd1 vccd1 vccd1 net6821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5560 rbzero.tex_r1\[20\] vssd1 vssd1 vccd1 vccd1 net6087 sky130_fd_sc_hd__dlygate4sd3_1
X_13051_ _06203_ _06206_ _06208_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__a21oi_1
Xhold5571 net905 vssd1 vssd1 vccd1 vccd1 net6098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5582 net925 vssd1 vssd1 vccd1 vccd1 net6109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5593 net998 vssd1 vssd1 vccd1 vccd1 net6120 sky130_fd_sc_hd__dlygate4sd3_1
X_12002_ net4127 _04468_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nand2_1
Xhold4870 _00861_ vssd1 vssd1 vccd1 vccd1 net5397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4881 net894 vssd1 vssd1 vccd1 vccd1 net5408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4892 rbzero.mapdyw\[0\] vssd1 vssd1 vccd1 vccd1 net5419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16810_ _06058_ _09836_ _09837_ vssd1 vssd1 vccd1 vccd1 _09838_ sky130_fd_sc_hd__o21ai_1
X_17790_ _02026_ _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16741_ _09773_ _09775_ _09776_ vssd1 vssd1 vccd1 vccd1 _09777_ sky130_fd_sc_hd__or3_1
X_13953_ _07122_ _07123_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19460_ net5452 _03334_ _03342_ _03339_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _06076_ _06077_ _06078_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__a211o_1
X_16672_ _09736_ vssd1 vssd1 vccd1 vccd1 _09741_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _07014_ _07015_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__and2_1
X_18411_ _02591_ _02592_ _04481_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a21o_1
X_15623_ _08221_ _08279_ _08318_ _08241_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__o22ai_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\] _06009_
+ _06010_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__or4_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _03205_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19754__36 clknet_1_0__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_0_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ net3509 net5961 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _08646_ _08647_ _08648_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__a21oi_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ net38 _05931_ _05934_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__a211o_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _07072_ _07233_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11717_ _04843_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nor2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ net4074 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15485_ _08389_ net8414 _08392_ _08161_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12697_ _05873_ _05874_ net31 vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17224_ _10241_ _10242_ vssd1 vssd1 vccd1 vccd1 _10244_ sky130_fd_sc_hd__nand2_1
X_11648_ _04837_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14436_ _07512_ _07555_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__03862_ clknet_0__03862_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03862_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
Xinput34 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_2
XFILLER_0_108_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17155_ _10173_ _10174_ vssd1 vssd1 vccd1 vccd1 _10175_ sky130_fd_sc_hd__nor2_1
Xinput45 i_reg_outs_enb vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_6
XFILLER_0_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11579_ _04765_ _04766_ _04768_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__nand3_1
X_14367_ _06924_ _07413_ net569 vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold807 net3737 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16106_ _09055_ _09072_ _09054_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__a21oi_1
Xhold818 _00592_ vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ _06465_ _06477_ _06484_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__or4_2
X_17086_ _10101_ _10106_ vssd1 vssd1 vccd1 vccd1 _10107_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14298_ _07464_ _07467_ _07468_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__a21o_1
Xhold829 _03830_ vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _09017_ _09022_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ _06264_ _06419_ _06307_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2208 net2622 vssd1 vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2219 _01053_ vssd1 vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1507 _01490_ vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1518 _01509_ vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ _02130_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__o21ba_1
Xhold1529 _03114_ vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
X_19727_ net5496 _03489_ net2310 vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a21boi_1
X_16939_ _09959_ _09960_ vssd1 vssd1 vccd1 vccd1 _09961_ sky130_fd_sc_hd__xnor2_1
X_19658_ net6432 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18609_ _05164_ net4423 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19589_ net1542 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21620_ clknet_leaf_128_i_clk net3188 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21551_ net185 net1954 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21482_ clknet_leaf_43_i_clk net1249 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4100 net8172 vssd1 vssd1 vccd1 vccd1 net4627 sky130_fd_sc_hd__dlygate4sd3_1
X_22103_ net165 net1978 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
Xhold4111 net684 vssd1 vssd1 vccd1 vccd1 net4638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4122 _09822_ vssd1 vssd1 vccd1 vccd1 net4649 sky130_fd_sc_hd__buf_4
XFILLER_0_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4133 net4265 vssd1 vssd1 vccd1 vccd1 net4660 sky130_fd_sc_hd__buf_1
X_20295_ net6452 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
Xhold4144 net8188 vssd1 vssd1 vccd1 vccd1 net4671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3410 _02982_ vssd1 vssd1 vccd1 vccd1 net3937 sky130_fd_sc_hd__dlygate4sd3_1
X_22034_ net476 net2961 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
Xhold3421 net4822 vssd1 vssd1 vccd1 vccd1 net3948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4166 net3425 vssd1 vssd1 vccd1 vccd1 net4693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4177 _07868_ vssd1 vssd1 vccd1 vccd1 net4704 sky130_fd_sc_hd__clkbuf_2
Xhold3432 net7686 vssd1 vssd1 vccd1 vccd1 net3959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4188 _04005_ vssd1 vssd1 vccd1 vccd1 net4715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3443 _03117_ vssd1 vssd1 vccd1 vccd1 net3970 sky130_fd_sc_hd__buf_1
Xhold3454 _00942_ vssd1 vssd1 vccd1 vccd1 net3981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4199 _02584_ vssd1 vssd1 vccd1 vccd1 net4726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2720 _04285_ vssd1 vssd1 vccd1 vccd1 net3247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3465 _03640_ vssd1 vssd1 vccd1 vccd1 net3992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2731 _01118_ vssd1 vssd1 vccd1 vccd1 net3258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3476 _03748_ vssd1 vssd1 vccd1 vccd1 net4003 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2742 net7535 vssd1 vssd1 vccd1 vccd1 net3269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3487 _00464_ vssd1 vssd1 vccd1 vccd1 net4014 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2753 _03068_ vssd1 vssd1 vccd1 vccd1 net3280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3498 _03786_ vssd1 vssd1 vccd1 vccd1 net4025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20526__266 clknet_1_1__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__inv_2
XFILLER_0_138_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2764 _00671_ vssd1 vssd1 vccd1 vccd1 net3291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2775 net3207 vssd1 vssd1 vccd1 vccd1 net3302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2786 _03579_ vssd1 vssd1 vccd1 vccd1 net3313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2797 _03050_ vssd1 vssd1 vccd1 vccd1 net3324 sky130_fd_sc_hd__dlygate4sd3_1
X_10950_ net6713 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10881_ net6756 net6092 _04253_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire80 _06655_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_6
X_12620_ net25 net24 vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__nor2_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21818_ net260 net1990 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ net4128 _05043_ _05730_ net3996 _05691_ net12 vssd1 vssd1 vccd1 vccd1 _05732_
+ sky130_fd_sc_hd__mux4_1
X_21749_ clknet_leaf_131_i_clk net4689 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11502_ net8207 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12482_ net4066 _05646_ _05642_ net71 _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a221o_1
X_15270_ _08124_ _08364_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14221_ _06696_ _07391_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nor2_1
X_11433_ _04525_ _04527_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14152_ _06699_ _07198_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11364_ rbzero.spi_registers.texadd3\[15\] rbzero.spi_registers.texadd1\[15\] rbzero.spi_registers.texadd0\[15\]
+ rbzero.spi_registers.texadd2\[15\] _04554_ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_
+ sky130_fd_sc_hd__mux4_2
Xhold6080 net1755 vssd1 vssd1 vccd1 vccd1 net6607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13103_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nor2_1
Xhold6091 rbzero.spi_registers.new_texadd\[0\]\[21\] vssd1 vssd1 vccd1 vccd1 net6618
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14083_ _07204_ _07249_ _07253_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a21oi_1
X_18960_ net1789 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5390 _02738_ vssd1 vssd1 vccd1 vccd1 net5917 sky130_fd_sc_hd__dlygate4sd3_1
X_17911_ _02145_ _02147_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__nand2_1
X_13034_ _06207_ net4526 _06209_ net4589 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a2bb2o_1
X_18891_ net1752 net7155 _03003_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17842_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__xnor2_1
X_17773_ _02010_ _02011_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _08090_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19512_ _03352_ net3218 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__nor2_1
X_16724_ _09753_ _09760_ _09761_ vssd1 vssd1 vccd1 vccd1 _09762_ sky130_fd_sc_hd__a21bo_1
X_13936_ _07105_ _07106_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__xor2_1
XFILLER_0_159_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19443_ net1561 net3519 _03141_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__and3_1
X_16655_ net3452 net3628 _09733_ vssd1 vssd1 vccd1 vccd1 _09734_ sky130_fd_sc_hd__or3_4
X_13867_ _07036_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15606_ _08694_ _08700_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__xnor2_4
X_12818_ _05978_ _05976_ _05977_ _05993_ _05991_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__o2111a_1
X_19374_ net6372 _03284_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__or2_1
X_16586_ net3587 _09413_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__nand2_1
X_13798_ _06962_ _06963_ _06967_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18325_ _02512_ net4714 _02511_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15537_ net3626 _08162_ _08167_ _08433_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__o211a_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _05904_ _05921_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7709 rbzero.debug_overlay.playerX\[0\] vssd1 vssd1 vccd1 vccd1 net8236 sky130_fd_sc_hd__dlygate4sd3_1
X_18256_ _02469_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__clkbuf_1
X_15468_ _08540_ _08562_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ _10224_ _10225_ _10106_ vssd1 vssd1 vccd1 vccd1 _10227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _07413_ _07233_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03845_ clknet_0__03845_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03845_
+ sky130_fd_sc_hd__clkbuf_16
X_18187_ _02403_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__inv_2
X_15399_ _08137_ net8042 vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__nand2_4
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _10155_ _10156_ vssd1 vssd1 vccd1 vccd1 _10158_ sky130_fd_sc_hd__and2_1
Xhold604 net6198 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 net6186 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _01125_ vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold637 net5469 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _01419_ vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 net6220 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ _10088_ _10089_ vssd1 vssd1 vccd1 vccd1 _10090_ sky130_fd_sc_hd__xor2_1
XFILLER_0_204_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20080_ net3433 _03660_ net4328 _03628_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__o211a_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _01528_ vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 _03576_ vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2027 net7195 vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2038 _01377_ vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1304 _03157_ vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2049 _04261_ vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 net7102 vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1326 net6734 vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1337 _00650_ vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 net6706 vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 _03570_ vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20982_ clknet_leaf_58_i_clk _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21603_ clknet_leaf_134_i_clk net3047 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21534_ clknet_leaf_130_i_clk net4946 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7__f_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21465_ clknet_leaf_17_i_clk net2600 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20416_ clknet_1_1__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__buf_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21396_ clknet_leaf_39_i_clk net5520 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11080_ net6950 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
X_20278_ _03689_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3240 net4905 vssd1 vssd1 vccd1 vccd1 net3767 sky130_fd_sc_hd__dlygate4sd3_1
X_22017_ net459 net1855 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3251 rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 net3778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3262 net7965 vssd1 vssd1 vccd1 vccd1 net3789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3273 _09870_ vssd1 vssd1 vccd1 vccd1 net3800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3284 net3295 vssd1 vssd1 vccd1 vccd1 net3811 sky130_fd_sc_hd__clkbuf_2
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3295 net3804 vssd1 vssd1 vccd1 vccd1 net3822 sky130_fd_sc_hd__clkbuf_2
Xhold2550 net2807 vssd1 vssd1 vccd1 vccd1 net3077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2561 _00932_ vssd1 vssd1 vccd1 vccd1 net3088 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 _03059_ vssd1 vssd1 vccd1 vccd1 net3099 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2583 rbzero.pov.spi_buffer\[10\] vssd1 vssd1 vccd1 vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03865_ clknet_0__03865_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03865_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2594 net1558 vssd1 vssd1 vccd1 vccd1 net3121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1860 net7203 vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1871 net4285 vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _07914_ _07935_ _07913_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__mux2_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1882 net6992 vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_11982_ _05143_ _05170_ _05121_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__o21ai_1
Xhold1893 net7130 vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13721_ _06783_ _06886_ _06890_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__a21oi_1
X_10933_ net7435 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _09524_ _09529_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10864_ net7431 net7145 _04171_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__mux2_1
X_13652_ _06791_ _06822_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__xor2_1
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ net19 _05760_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nor2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _09338_ _09444_ _09443_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__a21o_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ net7373 net7001 _04205_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__mux2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _06753_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18110_ _02341_ net3787 _02320_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
X_15322_ _08200_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__clkbuf_4
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _05711_ _05712_ _05697_ _05714_ net12 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__o221a_1
X_19090_ _09733_ net4096 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18041_ _02275_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__xor2_1
X_15253_ _08340_ _08347_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12465_ net6122 _05643_ _05644_ clknet_1_1__leaf__05645_ _05646_ vssd1 vssd1 vccd1
+ vccd1 _05647_ sky130_fd_sc_hd__a221o_2
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14204_ _07283_ _07320_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__xor2_2
X_11416_ _04553_ _04556_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__or2_1
X_12396_ _04967_ _05568_ _05572_ _04818_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o311a_1
X_15184_ _08277_ _08278_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14135_ _06771_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__clkbuf_4
X_11347_ _04515_ _04538_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19992_ _03484_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18943_ net7463 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
X_14066_ _07199_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__or2_1
X_11278_ net5922 vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13017_ net3820 _06191_ _06192_ net4655 vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_158_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18874_ _02992_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__clkbuf_4
X_20509__250 clknet_1_1__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__inv_2
X_17825_ _01997_ _02060_ _02061_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _01993_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14968_ net4483 _07991_ _08079_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16707_ _04489_ _09734_ vssd1 vssd1 vccd1 vccd1 _09747_ sky130_fd_sc_hd__or2_4
X_13919_ _07030_ _07070_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__nand2_1
X_17687_ _01815_ _01819_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14899_ net4277 _08037_ _08043_ vssd1 vssd1 vccd1 vccd1 _08044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19426_ net2060 net3651 _03310_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16638_ _08092_ vssd1 vssd1 vccd1 vccd1 _09725_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19357_ net6378 _03271_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__or2_1
X_16569_ _08880_ _09170_ _09403_ _08417_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18308_ net6530 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__clkbuf_1
Xhold7506 net8436 vssd1 vssd1 vccd1 vccd1 net8033 sky130_fd_sc_hd__clkbuf_2
Xhold7517 _08313_ vssd1 vssd1 vccd1 vccd1 net8044 sky130_fd_sc_hd__dlygate4sd3_1
X_19288_ net8118 _03236_ net598 _03230_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7528 _08274_ vssd1 vssd1 vccd1 vccd1 net8055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7539 rbzero.traced_texa\[9\] vssd1 vssd1 vccd1 vccd1 net8066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6805 net2345 vssd1 vssd1 vccd1 vccd1 net7332 sky130_fd_sc_hd__dlygate4sd3_1
X_18239_ _09788_ _02454_ _02155_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a21o_1
Xhold6816 rbzero.tex_b1\[43\] vssd1 vssd1 vccd1 vccd1 net7343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6827 rbzero.tex_g0\[55\] vssd1 vssd1 vccd1 vccd1 net7354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6838 net2780 vssd1 vssd1 vccd1 vccd1 net7365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6849 rbzero.tex_b0\[48\] vssd1 vssd1 vccd1 vccd1 net7376 sky130_fd_sc_hd__dlygate4sd3_1
X_21250_ clknet_leaf_7_i_clk net3594 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold401 net5221 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 net6104 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 net7885 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20201_ net3494 net1875 _03709_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__mux2_1
Xhold434 net4278 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 net8070 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03859_ _03859_ vssd1 vssd1 vccd1 vccd1 clknet_0__03859_ sky130_fd_sc_hd__clkbuf_16
X_21181_ clknet_leaf_128_i_clk net3058 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold456 net5273 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold467 net5289 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
X_20132_ rbzero.debug_overlay.facingX\[-5\] net3435 _03710_ vssd1 vssd1 vccd1 vccd1
+ _03716_ sky130_fd_sc_hd__mux2_1
Xhold478 net5417 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 net8004 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20063_ net4616 _08145_ _03614_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__mux2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 net6565 vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 _00960_ vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 net6620 vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 net6700 vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 _03370_ vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 net6694 vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 net6503 vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 _00714_ vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _04306_ vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ clknet_leaf_71_i_clk _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20896_ _03312_ net1099 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ net6930 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21517_ clknet_leaf_5_i_clk net1336 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ _04921_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21448_ clknet_leaf_19_i_clk net3625 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_other
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ net6830 net2527 _04423_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _05258_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__buf_4
X_21379_ clknet_leaf_9_i_clk net5011 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ net6946 net2648 _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
Xhold990 net6825 vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ net6866 net2632 _04353_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__mux2_1
X_15940_ net3453 _09033_ _09034_ _08442_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__a31o_1
Xhold3070 _03093_ vssd1 vssd1 vccd1 vccd1 net3597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3081 net7652 vssd1 vssd1 vccd1 vccd1 net3608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3092 _02762_ vssd1 vssd1 vccd1 vccd1 net3619 sky130_fd_sc_hd__clkbuf_4
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ _08942_ _08959_ _08961_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__a21bo_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2380 net2810 vssd1 vssd1 vccd1 vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
X_17610_ _01732_ _01735_ _01733_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2391 _04439_ vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ net4496 _07981_ _07976_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__mux2_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ net4528 net4848 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__nor2_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03848_ clknet_0__03848_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03848_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 net7070 vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
X_17541_ _01690_ _01681_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or2b_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _07843_ _07820_ _07842_ _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ rbzero.debug_overlay.vplaneX\[0\] _05093_ _05095_ rbzero.debug_overlay.vplaneX\[-3\]
+ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _06683_ _06737_ _06634_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21oi_1
X_17472_ _10392_ _01713_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__xnor2_1
X_10916_ net7423 net6854 _04276_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14684_ net8442 _07854_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ net4108 _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19211_ net6516 _03183_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or2_1
X_16423_ _09383_ _09384_ _09381_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _06801_ _06804_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10847_ net2400 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19142_ net5432 _03145_ _03154_ _03149_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__o211a_1
X_16354_ _09338_ _09445_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_184_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13566_ _06736_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10778_ _04193_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ _08359_ _08399_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__xnor2_2
X_19073_ _04458_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__buf_4
X_12517_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__inv_2
X_16285_ _09374_ _09375_ _09376_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13497_ _06606_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18024_ _02174_ _02177_ _02175_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15236_ _08280_ _08294_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12448_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ net3457 _08236_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__nand2_1
X_12379_ _05306_ _05559_ _05563_ _05263_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a211o_1
XFILLER_0_205_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _06923_ _07259_ _06693_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19975_ net7312 net1866 _09725_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__mux2_1
X_15098_ net4268 _08118_ _06119_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14049_ _07209_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__xnor2_1
X_18926_ net6438 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18857_ net3330 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17808_ _01962_ _01963_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a21oi_1
X_18788_ _02933_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nand2_1
X_17739_ _01975_ _01976_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__and2_1
XFILLER_0_203_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20750_ net822 net4980 vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19409_ net5509 _03302_ _03309_ _03299_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8015 _09092_ vssd1 vssd1 vccd1 vccd1 net8542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7303 rbzero.wall_tracer.stepDistX\[2\] vssd1 vssd1 vccd1 vccd1 net7830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7314 net3748 vssd1 vssd1 vccd1 vccd1 net7841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7325 net4378 vssd1 vssd1 vccd1 vccd1 net7852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7336 net647 vssd1 vssd1 vccd1 vccd1 net7863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6602 net2032 vssd1 vssd1 vccd1 vccd1 net7129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7347 rbzero.wall_tracer.stepDistX\[4\] vssd1 vssd1 vccd1 vccd1 net7874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6613 rbzero.tex_r0\[55\] vssd1 vssd1 vccd1 vccd1 net7140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7358 net4201 vssd1 vssd1 vccd1 vccd1 net7885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7369 rbzero.traced_texVinit\[4\] vssd1 vssd1 vccd1 vccd1 net7896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6624 net2295 vssd1 vssd1 vccd1 vccd1 net7151 sky130_fd_sc_hd__dlygate4sd3_1
X_21302_ clknet_leaf_48_i_clk net5366 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6635 _04055_ vssd1 vssd1 vccd1 vccd1 net7162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6646 net2403 vssd1 vssd1 vccd1 vccd1 net7173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5901 net1448 vssd1 vssd1 vccd1 vccd1 net6428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6657 net2676 vssd1 vssd1 vccd1 vccd1 net7184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5912 rbzero.spi_registers.new_texadd\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net6439
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5923 net1465 vssd1 vssd1 vccd1 vccd1 net6450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6668 rbzero.tex_b1\[42\] vssd1 vssd1 vccd1 vccd1 net7195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6679 net2388 vssd1 vssd1 vccd1 vccd1 net7206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5934 _04408_ vssd1 vssd1 vccd1 vccd1 net6461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 net4688 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
X_21233_ clknet_leaf_123_i_clk net1615 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5945 net986 vssd1 vssd1 vccd1 vccd1 net6472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5956 rbzero.spi_registers.new_texadd\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net6483
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 net5259 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 net5112 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5967 net1061 vssd1 vssd1 vccd1 vccd1 net6494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5978 rbzero.tex_g0\[18\] vssd1 vssd1 vccd1 vccd1 net6505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 net4515 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 net7187 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ clknet_leaf_131_i_clk net1575 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5989 net1570 vssd1 vssd1 vccd1 vccd1 net6516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 net5269 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 net5170 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 net5211 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20115_ net5759 _03615_ _03659_ _03703_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__o211a_1
X_21095_ clknet_leaf_11_i_clk net1437 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20046_ _03483_ _03650_ _03608_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a21o_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ net439 net2189 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _04932_ _04935_ _04939_ _04928_ net84 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a221o_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ clknet_leaf_66_i_clk _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ net5690 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__clkbuf_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _04462_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20879_ _02752_ _02758_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__or2b_1
XFILLER_0_181_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13420_ net561 net560 _06496_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a21oi_1
X_10632_ net6174 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10563_ net1116 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _04915_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__or2_1
X_16070_ _08401_ _08402_ _09025_ _09031_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__or4_1
Xhold7870 _08201_ vssd1 vssd1 vccd1 vccd1 net8397 sky130_fd_sc_hd__dlygate4sd3_1
X_10494_ net2500 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _06451_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__xnor2_2
X_15021_ net3628 _06117_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__or2b_1
X_12233_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _04838_ vssd1 vssd1 vccd1 vccd1 _05420_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12164_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _05239_ vssd1 vssd1 vccd1 vccd1 _05352_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11115_ net2149 net6052 _04375_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__mux2_1
X_16972_ _09991_ _09993_ vssd1 vssd1 vccd1 vccd1 _09994_ sky130_fd_sc_hd__nor2_1
X_12095_ _04849_ _05224_ _05244_ _05265_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__o32a_1
XFILLER_0_21_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11046_ net7346 net7401 _04342_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
X_15923_ _08221_ _08241_ _08418_ _08392_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__or4_1
X_18711_ net8113 _02537_ _02855_ net4799 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__o211ai_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19691_ net1463 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__clkbuf_1
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18642_ net3678 rbzero.wall_tracer.rayAddendY\[-2\] _02791_ vssd1 vssd1 vccd1 vccd1
+ _02799_ sky130_fd_sc_hd__o21a_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _08948_ _08329_ _08691_ _08916_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__o22a_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _07914_ _07935_ _07965_ _07966_ net531 net7785 vssd1 vssd1 vccd1 vccd1 _07967_
+ sky130_fd_sc_hd__mux4_2
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ net5916 _02737_ _09788_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
X_15785_ _08221_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__buf_2
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12997_ _06164_ net3787 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nor2_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17524_ _01763_ _01764_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__nand2_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _07904_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11948_ rbzero.debug_overlay.facingX\[-6\] _05102_ _05090_ rbzero.debug_overlay.facingX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _10105_ _01692_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a21oi_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ net564 _07834_ _07836_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__nand3_1
X_11879_ net4106 net4058 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16406_ _09467_ _09496_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13618_ _06747_ _06748_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17386_ _10402_ _10403_ vssd1 vssd1 vccd1 vccd1 _10404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _07767_ _07766_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19125_ net886 _03140_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__and2_1
X_16337_ _09426_ _09428_ vssd1 vssd1 vccd1 vccd1 _09429_ sky130_fd_sc_hd__xnor2_1
X_13549_ net567 _06634_ net79 net80 vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a211o_2
XFILLER_0_82_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19056_ net7585 net7579 net3397 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
X_16268_ _09251_ _09256_ _09359_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__05794_ _05794_ vssd1 vssd1 vccd1 vccd1 clknet_0__05794_ sky130_fd_sc_hd__clkbuf_16
Xhold5208 net2941 vssd1 vssd1 vccd1 vccd1 net5735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5219 _03612_ vssd1 vssd1 vccd1 vccd1 net5746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18007_ _02242_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15219_ _08114_ net8044 vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__nand2_1
Xhold4507 _01647_ vssd1 vssd1 vccd1 vccd1 net5034 sky130_fd_sc_hd__dlygate4sd3_1
X_16199_ net3841 _06122_ _09181_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__a21boi_4
Xhold4518 net610 vssd1 vssd1 vccd1 vccd1 net5045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4529 rbzero.spi_registers.texadd1\[20\] vssd1 vssd1 vccd1 vccd1 net5056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3806 _00434_ vssd1 vssd1 vccd1 vccd1 net4333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3817 net8215 vssd1 vssd1 vccd1 vccd1 net4344 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3828 _00767_ vssd1 vssd1 vccd1 vccd1 net4355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_i_clk clknet_4_0__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold3839 net8167 vssd1 vssd1 vccd1 vccd1 net4366 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20366__121 clknet_1_1__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__inv_2
X_19958_ net2191 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
X_18909_ net2486 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
X_19889_ net3074 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
X_21920_ net362 net3106 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
X_21851_ net293 net2136 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20802_ _03964_ _03965_ _03966_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21782_ clknet_leaf_6_i_clk net1687 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20733_ net1106 net5340 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7100 net3504 vssd1 vssd1 vccd1 vccd1 net7627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7122 _03499_ vssd1 vssd1 vccd1 vccd1 net7649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7133 net3436 vssd1 vssd1 vccd1 vccd1 net7660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7144 net3808 vssd1 vssd1 vccd1 vccd1 net7671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6410 rbzero.spi_registers.new_leak\[0\] vssd1 vssd1 vccd1 vccd1 net6937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7155 _01247_ vssd1 vssd1 vccd1 vccd1 net7682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6421 net2274 vssd1 vssd1 vccd1 vccd1 net6948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7166 rbzero.spi_registers.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 net7693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6432 rbzero.spi_registers.new_vshift\[5\] vssd1 vssd1 vccd1 vccd1 net6959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7177 rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1 net7704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6443 _04453_ vssd1 vssd1 vccd1 vccd1 net6970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7188 gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 net7715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6454 net2340 vssd1 vssd1 vccd1 vccd1 net6981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7199 _05548_ vssd1 vssd1 vccd1 vccd1 net7726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6465 _04212_ vssd1 vssd1 vccd1 vccd1 net6992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5720 net1182 vssd1 vssd1 vccd1 vccd1 net6247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5731 rbzero.tex_r1\[35\] vssd1 vssd1 vccd1 vccd1 net6258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6476 net1970 vssd1 vssd1 vccd1 vccd1 net7003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5742 net1412 vssd1 vssd1 vccd1 vccd1 net6269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6487 rbzero.tex_g1\[47\] vssd1 vssd1 vccd1 vccd1 net7014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6498 net1929 vssd1 vssd1 vccd1 vccd1 net7025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5753 rbzero.spi_registers.new_texadd\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 net6280
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21216_ clknet_leaf_121_i_clk net3225 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5764 net1281 vssd1 vssd1 vccd1 vccd1 net6291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5775 _03448_ vssd1 vssd1 vccd1 vccd1 net6302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5786 net1310 vssd1 vssd1 vccd1 vccd1 net6313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5797 rbzero.spi_registers.new_texadd\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net6324
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21147_ clknet_leaf_104_i_clk net4810 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_21078_ clknet_leaf_76_i_clk _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20029_ net3443 _03609_ net5869 _03316_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a211o_1
X_12920_ net2587 _06061_ net4642 net4366 _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ _05985_ net7775 vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nand2_4
XFILLER_0_186_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ _04967_ _04975_ _04990_ _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a211o_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _08634_ _08660_ _08664_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__or2_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _07689_ _07690_ _07691_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nor3b_2
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _04836_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__buf_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ net4648 vssd1 vssd1 vccd1 vccd1 _10260_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _06699_ _07457_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ net3405 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13403_ _06563_ _06569_ _06570_ _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__a211o_1
X_10615_ net2960 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__clkbuf_1
X_17171_ _10190_ _08616_ vssd1 vssd1 vccd1 vccd1 _10191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14383_ _07532_ _07552_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11595_ net1023 net4312 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16122_ net4612 _08115_ _08038_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__o21ai_1
X_13334_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__clkbuf_4
X_10546_ net6717 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _09144_ _09145_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13265_ net559 vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__buf_2
X_10477_ net2689 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _06115_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__inv_2
X_12216_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _04951_ vssd1 vssd1 vccd1 vccd1 _05403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ _06355_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12147_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _04978_ vssd1 vssd1 vccd1 vccd1 _05335_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19743_ clknet_1_0__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__buf_1
X_12078_ rbzero.tex_r1\[49\] rbzero.tex_r1\[48\] _04979_ vssd1 vssd1 vccd1 vccd1 _05267_
+ sky130_fd_sc_hd__mux2_1
X_16955_ _08905_ _09976_ _09972_ vssd1 vssd1 vccd1 vccd1 _09977_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ net6118 net2735 _04331_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux2_1
X_15906_ _08999_ _09000_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__and2_1
X_16886_ _08864_ _09354_ _09618_ _09617_ _09506_ vssd1 vssd1 vccd1 vccd1 _09908_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19674_ net1417 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15837_ _08925_ _08928_ _08929_ _08931_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__o211a_1
X_18625_ _02782_ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__or2b_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15768_ _08280_ _08458_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__nor2_1
X_18556_ net3552 _09818_ _02723_ _02724_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17507_ _09915_ _09345_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__or2_1
X_14719_ _07841_ _07888_ _07843_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__a21o_1
X_18487_ rbzero.wall_tracer.rayAddendX\[6\] _02663_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02665_ sky130_fd_sc_hd__mux2_1
X_15699_ _08739_ _08766_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__nand2_1
X_17438_ _10429_ _01679_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__xnor2_1
XANTENNA_15 _09094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_37 net3592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_48 _04021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17369_ _10385_ _10386_ vssd1 vssd1 vccd1 vccd1 _10387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_59 _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19108_ net2185 _03125_ net5571 _03128_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5005 _00387_ vssd1 vssd1 vccd1 vccd1 net5532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5016 net2039 vssd1 vssd1 vccd1 vccd1 net5543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19039_ net3746 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5027 net2006 vssd1 vssd1 vccd1 vccd1 net5554 sky130_fd_sc_hd__buf_1
Xhold5038 net1852 vssd1 vssd1 vccd1 vccd1 net5565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5049 net2286 vssd1 vssd1 vccd1 vccd1 net5576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4304 rbzero.spi_registers.spi_cmd\[1\] vssd1 vssd1 vccd1 vccd1 net4831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4315 net1043 vssd1 vssd1 vccd1 vccd1 net4842 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22050_ net492 net1385 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold4326 _01650_ vssd1 vssd1 vccd1 vccd1 net4853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4337 _06055_ vssd1 vssd1 vccd1 vccd1 net4864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3603 _01248_ vssd1 vssd1 vccd1 vccd1 net4130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4348 net3931 vssd1 vssd1 vccd1 vccd1 net4875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4359 rbzero.wall_tracer.rayAddendX\[-7\] vssd1 vssd1 vccd1 vccd1 net4886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3614 _05462_ vssd1 vssd1 vccd1 vccd1 net4141 sky130_fd_sc_hd__clkbuf_4
X_21001_ clknet_leaf_85_i_clk _00488_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3625 net5754 vssd1 vssd1 vccd1 vccd1 net4152 sky130_fd_sc_hd__buf_1
Xhold3636 _05047_ vssd1 vssd1 vccd1 vccd1 net4163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3647 _08098_ vssd1 vssd1 vccd1 vccd1 net4174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2902 net4731 vssd1 vssd1 vccd1 vccd1 net3429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2913 net2758 vssd1 vssd1 vccd1 vccd1 net3440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3658 rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 net4185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3669 _00850_ vssd1 vssd1 vccd1 vccd1 net4196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2924 net3974 vssd1 vssd1 vccd1 vccd1 net3451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2935 net4493 vssd1 vssd1 vccd1 vccd1 net3462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2946 net7634 vssd1 vssd1 vccd1 vccd1 net3473 sky130_fd_sc_hd__clkbuf_4
Xhold2957 net7831 vssd1 vssd1 vccd1 vccd1 net3484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2968 _03760_ vssd1 vssd1 vccd1 vccd1 net3495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2979 _01210_ vssd1 vssd1 vccd1 vccd1 net3506 sky130_fd_sc_hd__dlygate4sd3_1
X_21903_ net345 net1966 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21834_ net276 net1354 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20420__170 clknet_1_1__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__inv_2
X_21765_ clknet_leaf_83_i_clk net4100 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20716_ _03895_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__and2b_1
XFILLER_0_191_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21696_ clknet_leaf_115_i_clk net4620 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ _04503_ _04564_ _04565_ _04571_ _04496_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__o311a_1
XFILLER_0_34_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6240 rbzero.tex_b0\[17\] vssd1 vssd1 vccd1 vccd1 net6767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6251 net1921 vssd1 vssd1 vccd1 vccd1 net6778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6262 _04409_ vssd1 vssd1 vccd1 vccd1 net6789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6273 net1997 vssd1 vssd1 vccd1 vccd1 net6800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6284 rbzero.tex_g1\[41\] vssd1 vssd1 vccd1 vccd1 net6811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6295 net2101 vssd1 vssd1 vccd1 vccd1 net6822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5550 _03480_ vssd1 vssd1 vccd1 vccd1 net6077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5561 net933 vssd1 vssd1 vccd1 vccd1 net6088 sky130_fd_sc_hd__dlygate4sd3_1
X_13050_ _06185_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_116_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold5572 gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5583 gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12001_ net4091 _04682_ net4095 _04022_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__or4_1
Xhold5594 gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4860 rbzero.spi_registers.texadd1\[10\] vssd1 vssd1 vccd1 vccd1 net5387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4871 net996 vssd1 vssd1 vccd1 vccd1 net5398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4882 _00390_ vssd1 vssd1 vccd1 vccd1 net5409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4893 net1013 vssd1 vssd1 vccd1 vccd1 net5420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ net4049 net3884 net5666 net5554 _09102_ vssd1 vssd1 vccd1 vccd1 _09776_ sky130_fd_sc_hd__o41a_1
X_13952_ _06719_ _06698_ _07121_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ net2968 net1161 net832 net1611 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__or4_1
X_16671_ net4361 _09737_ _09740_ _07981_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20503__245 clknet_1_1__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__inv_2
XFILLER_0_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13883_ _07051_ _07053_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and2_1
X_15622_ _08266_ _08328_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__nor2_1
X_18410_ _02591_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12834_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__xor2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19390_ net6180 _03270_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _02519_ _02520_ _02521_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__o21a_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _08627_ _08645_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__nor2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ net38 _05937_ _05939_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and4b_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _07413_ _07198_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__nor2_1
X_11716_ net7569 _04905_ _04821_ net5509 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ net6337 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__clkbuf_1
X_15484_ _08161_ _08168_ net8414 _08384_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12696_ _04020_ _04495_ net7678 _04500_ net28 _05850_ vssd1 vssd1 vccd1 vccd1 _05874_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17223_ _10241_ _10242_ vssd1 vssd1 vccd1 vccd1 _10243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ _07560_ _07605_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__nor2_1
X_11647_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__03861_ clknet_0__03861_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03861_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_4
X_17154_ _10039_ _10048_ _10046_ vssd1 vssd1 vccd1 vccd1 _10174_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
Xinput35 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14366_ _07488_ _07494_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__xnor2_4
X_11578_ net1284 _04766_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand3_1
Xinput46 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_6
X_16105_ _09129_ _09198_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold808 _03473_ vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
X_13317_ _06485_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__or2_1
X_10529_ net2982 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__clkbuf_1
X_17085_ _10102_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _10106_ sky130_fd_sc_hd__o21a_2
Xhold819 net6439 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
X_14297_ _07402_ _07405_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__xnor2_1
X_16036_ _09001_ _09010_ _09008_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__a21o_1
X_20584__317 clknet_1_0__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__inv_2
XFILLER_0_161_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13248_ net8068 _06266_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _06347_ _06349_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _06350_
+ sky130_fd_sc_hd__mux2_4
Xhold2209 _04337_ vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1508 net6923 vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_80_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17987_ _02109_ _02110_ _02107_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1519 net3792 vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
X_19726_ net3705 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__clkbuf_1
X_16938_ _09272_ _09165_ vssd1 vssd1 vccd1 vccd1 _09960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19657_ net6430 net3583 _03429_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux2_1
X_16869_ _09630_ _09889_ _09890_ vssd1 vssd1 vccd1 vccd1 _09891_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_95_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18608_ net8129 _02508_ _09739_ net4531 _02768_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a221o_1
X_20478__222 clknet_1_1__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__inv_2
XFILLER_0_181_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19588_ net6597 net3596 net1779 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__mux2_1
X_18539_ net3893 _06041_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21550_ net184 net2347 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21481_ clknet_leaf_43_i_clk net1213 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4101 net3408 vssd1 vssd1 vccd1 vccd1 net4628 sky130_fd_sc_hd__dlygate4sd3_1
X_22102_ net164 net2853 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
Xhold4112 net8346 vssd1 vssd1 vccd1 vccd1 net4639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4123 net7969 vssd1 vssd1 vccd1 vccd1 net4650 sky130_fd_sc_hd__dlygate4sd3_1
X_20294_ net6450 net2204 _03814_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4134 _08063_ vssd1 vssd1 vccd1 vccd1 net4661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4145 _00415_ vssd1 vssd1 vccd1 vccd1 net4672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3400 rbzero.debug_overlay.facingY\[0\] vssd1 vssd1 vccd1 vccd1 net3927 sky130_fd_sc_hd__dlygate4sd3_1
X_22033_ net475 net2446 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
Xhold4156 _08048_ vssd1 vssd1 vccd1 vccd1 net4683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3411 _00643_ vssd1 vssd1 vccd1 vccd1 net3938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3422 rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 net3949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4167 net4299 vssd1 vssd1 vccd1 vccd1 net4694 sky130_fd_sc_hd__clkbuf_2
Xhold4178 net4225 vssd1 vssd1 vccd1 vccd1 net4705 sky130_fd_sc_hd__buf_4
Xhold3433 _06081_ vssd1 vssd1 vccd1 vccd1 net3960 sky130_fd_sc_hd__clkbuf_2
Xhold4189 net8106 vssd1 vssd1 vccd1 vccd1 net4716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3444 net7682 vssd1 vssd1 vccd1 vccd1 net3971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2710 net3191 vssd1 vssd1 vccd1 vccd1 net3237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3455 net5504 vssd1 vssd1 vccd1 vccd1 net3982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2721 _01371_ vssd1 vssd1 vccd1 vccd1 net3248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3466 net5909 vssd1 vssd1 vccd1 vccd1 net3993 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_48_i_clk clknet_4_8__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2732 rbzero.pov.spi_buffer\[42\] vssd1 vssd1 vccd1 vccd1 net3259 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3477 _03749_ vssd1 vssd1 vccd1 vccd1 net4004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3488 net4037 vssd1 vssd1 vccd1 vccd1 net4015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 _03062_ vssd1 vssd1 vccd1 vccd1 net3270 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2754 _00715_ vssd1 vssd1 vccd1 vccd1 net3281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3499 _01245_ vssd1 vssd1 vccd1 vccd1 net4026 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2765 net3341 vssd1 vssd1 vccd1 vccd1 net3292 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2776 _03551_ vssd1 vssd1 vccd1 vccd1 net3303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2787 _01142_ vssd1 vssd1 vccd1 vccd1 net3314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2798 _00698_ vssd1 vssd1 vccd1 vccd1 net3325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10880_ net2692 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21817_ net259 net2241 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ net6044 vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__buf_1
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21748_ clknet_leaf_132_i_clk net3578 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11501_ _04671_ _04673_ _04676_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and4_1
X_12481_ net50 _05643_ _05644_ net49 _05649_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21679_ clknet_leaf_124_i_clk net3307 vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14220_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ _04525_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ _07283_ _07320_ _07321_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_85_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ _04505_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6070 net1203 vssd1 vssd1 vccd1 vccd1 net6597 sky130_fd_sc_hd__dlygate4sd3_1
X_13102_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] _06271_
+ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a31oi_2
Xhold6081 _04094_ vssd1 vssd1 vccd1 vccd1 net6608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14082_ _07250_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__nand2_1
Xhold6092 net1649 vssd1 vssd1 vccd1 vccd1 net6619 sky130_fd_sc_hd__dlygate4sd3_1
X_11294_ _04478_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__buf_4
Xhold5380 net5791 vssd1 vssd1 vccd1 vccd1 net5907 sky130_fd_sc_hd__dlygate4sd3_1
X_17910_ _02145_ _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13033_ net3751 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__inv_2
Xhold5391 _02739_ vssd1 vssd1 vccd1 vccd1 net5918 sky130_fd_sc_hd__dlygate4sd3_1
X_18890_ net7047 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4690 _00836_ vssd1 vssd1 vccd1 vccd1 net5217 sky130_fd_sc_hd__dlygate4sd3_1
X_17841_ net8008 _09181_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17772_ _02008_ _02009_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__and2_1
X_14984_ net4388 _08030_ _08067_ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19511_ net5978 _03139_ _03364_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13935_ _06576_ _06832_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16723_ net3999 _09102_ vssd1 vssd1 vccd1 vccd1 _09761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19442_ net3646 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__clkbuf_1
X_16654_ net4122 vssd1 vssd1 vccd1 vccd1 _09733_ sky130_fd_sc_hd__inv_2
X_13866_ _06706_ _06796_ _07035_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__o21ai_1
X_15605_ _08697_ _08699_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__xnor2_4
X_12817_ _05978_ net3761 net4416 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__nand3b_1
X_16585_ net8035 _08494_ _09673_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__or3b_1
X_19373_ net5001 _03283_ _03289_ _03288_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13797_ _06962_ _06963_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__nand3_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15536_ _08372_ _08373_ net4877 _08630_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__or4_1
X_18324_ net4713 net693 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ net35 _05905_ _05922_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a31o_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18255_ _02468_ net4498 net4782 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_4
X_15467_ _08541_ _08561_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ net31 vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17206_ _10106_ _10224_ _10225_ vssd1 vssd1 vccd1 vccd1 _10226_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418_ _07539_ _07540_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03844_ clknet_0__03844_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03844_
+ sky130_fd_sc_hd__clkbuf_16
X_18186_ net3766 net4481 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__or2_1
X_15398_ _06121_ net4877 _08366_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17137_ _10155_ _10156_ vssd1 vssd1 vccd1 vccd1 _10157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14349_ _07514_ _07517_ _07518_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nand3_1
Xhold605 _01353_ vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 net6188 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 net4611 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold638 net6238 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17068_ _08509_ _09170_ vssd1 vssd1 vccd1 vccd1 _10089_ sky130_fd_sc_hd__or2_1
Xhold649 net6463 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16019_ _09111_ _09112_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 net7380 vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 _01139_ vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2028 net7197 vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 net6990 vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 net4394 vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 _04110_ vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1327 net6736 vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1338 rbzero.pov.mosi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1349 net6708 vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19709_ net6134 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
X_20981_ clknet_leaf_57_i_clk _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21602_ clknet_leaf_134_i_clk net2508 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21533_ clknet_leaf_130_i_clk net3826 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21464_ clknet_leaf_17_i_clk net2646 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20532__271 clknet_1_1__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__inv_2
XFILLER_0_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21395_ clknet_leaf_39_i_clk net5503 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20277_ net5966 net4099 vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3230 net3409 vssd1 vssd1 vccd1 vccd1 net3757 sky130_fd_sc_hd__clkbuf_2
Xhold3241 net3012 vssd1 vssd1 vccd1 vccd1 net3768 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22016_ net458 net2096 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3252 net5953 vssd1 vssd1 vccd1 vccd1 net3779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3263 net3205 vssd1 vssd1 vccd1 vccd1 net3790 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3274 net7958 vssd1 vssd1 vccd1 vccd1 net3801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2540 net2393 vssd1 vssd1 vccd1 vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3296 net7654 vssd1 vssd1 vccd1 vccd1 net3823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2551 _03535_ vssd1 vssd1 vccd1 vccd1 net3078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2562 net7432 vssd1 vssd1 vccd1 vccd1 net3089 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 _00706_ vssd1 vssd1 vccd1 vccd1 net3100 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03864_ clknet_0__03864_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03864_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2584 net3101 vssd1 vssd1 vccd1 vccd1 net3111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1850 net7138 vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2595 _03578_ vssd1 vssd1 vccd1 vccd1 net3122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1861 net7205 vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1872 net7048 vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
X_11981_ _05150_ _05169_ _04670_ net4161 vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__o2bb2a_1
Xhold1883 _01437_ vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1894 net7132 vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ _06783_ _06886_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__and3_1
X_10932_ net7433 net3263 _04276_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ _06807_ _06821_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10863_ net6589 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__buf_1
XFILLER_0_151_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12602_ net18 _05775_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__o21ai_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _09446_ _09447_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _06701_ _06705_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__xor2_1
X_10794_ net2567 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _08412_ _08415_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__nand2_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ net54 _05713_ net50 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a21oi_1
X_20615__346 clknet_1_1__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__inv_2
XFILLER_0_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _02201_ _02211_ _02209_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _08342_ _08345_ _08346_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_48_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12464_ net5 _05633_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ _07345_ _07373_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11415_ _04496_ _04552_ _04604_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__o31a_1
X_15183_ net4485 _08136_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__nor2_1
X_12395_ _05574_ _05576_ _05579_ _05465_ _05263_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14134_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__buf_2
X_11346_ rbzero.texu_hot\[5\] _04514_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or2_1
X_19991_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18942_ net3166 net7461 _03036_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
X_14065_ _07234_ _07235_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11277_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ net3835 vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18873_ net3020 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ _01997_ _02060_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20360__116 clknet_1_0__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__inv_2
X_17755_ _01991_ _01992_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__and2_1
X_14967_ _08081_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16706_ net8079 _09745_ _09746_ net8034 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a22o_1
X_13918_ _07032_ _07085_ _07087_ _07088_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__or4_4
X_17686_ _01818_ _01925_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14898_ _04481_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__clkbuf_4
X_19425_ _08092_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13849_ _07006_ _07018_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__o21bai_1
X_16637_ net3955 net3858 vssd1 vssd1 vccd1 vccd1 _09724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19356_ net5396 _03269_ _03279_ _03275_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__o211a_1
X_16568_ _09403_ _08244_ _08666_ _09288_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__and4b_1
XFILLER_0_18_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ net6528 net3866 _02493_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
X_15519_ _08613_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__clkbuf_4
X_16499_ _09460_ _09587_ _09588_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__o21ai_4
Xhold7507 net7816 vssd1 vssd1 vccd1 vccd1 net8034 sky130_fd_sc_hd__clkbuf_4
X_19287_ net597 _03238_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__or2_1
Xhold7518 _08314_ vssd1 vssd1 vccd1 vccd1 net8045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7529 rbzero.wall_tracer.stepDistY\[-3\] vssd1 vssd1 vccd1 vccd1 net8056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6806 rbzero.pov.ready_buffer\[40\] vssd1 vssd1 vccd1 vccd1 net7333 sky130_fd_sc_hd__dlygate4sd3_1
X_18238_ _02452_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6817 net2937 vssd1 vssd1 vccd1 vccd1 net7344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6828 net2923 vssd1 vssd1 vccd1 vccd1 net7355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6839 rbzero.pov.spi_buffer\[51\] vssd1 vssd1 vccd1 vccd1 net7366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18169_ _02392_ net3790 _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
Xhold402 net5363 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _01071_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20200_ net7155 _03743_ net4699 _03732_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__03858_ _03858_ vssd1 vssd1 vccd1 vccd1 clknet_0__03858_ sky130_fd_sc_hd__clkbuf_16
X_21180_ clknet_leaf_101_i_clk net1948 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold424 net5391 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold435 net5323 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold446 net5279 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 net8180 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 net5395 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
X_20131_ net3362 _03707_ net4463 _03679_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold479 net5427 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20062_ net5929 _03660_ net3441 _03628_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__o211a_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 net6567 vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 net5525 vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _00987_ vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 _01301_ vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _00922_ vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20562__297 clknet_1_0__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__inv_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1157 _00653_ vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1168 _03461_ vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1179 net1751 vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ clknet_leaf_73_i_clk _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ net4936 net6111 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21516_ clknet_leaf_6_i_clk net1464 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21447_ clknet_leaf_25_i_clk net1766 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ net6098 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _04821_ _05350_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or3_2
X_21378_ clknet_leaf_9_i_clk net5023 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11131_ _04264_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__clkbuf_4
X_20329_ net6180 net3583 _03813_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold980 _00593_ vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 net6827 vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net5591 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
Xhold3060 net8343 vssd1 vssd1 vccd1 vccd1 net3587 sky130_fd_sc_hd__buf_1
Xhold3071 _00734_ vssd1 vssd1 vccd1 vccd1 net3598 sky130_fd_sc_hd__dlygate4sd3_1
X_15870_ _08943_ _08964_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__xnor2_1
Xhold3082 _03721_ vssd1 vssd1 vccd1 vccd1 net3609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3093 _03771_ vssd1 vssd1 vccd1 vccd1 net3620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2370 _01024_ vssd1 vssd1 vccd1 vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2381 _04176_ vssd1 vssd1 vccd1 vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
X_14821_ net7824 _07979_ _07980_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__a21o_2
XFILLER_0_203_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2392 _01039_ vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03847_ clknet_0__03847_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03847_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1680 _00950_ vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1691 net7072 vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
X_17540_ _01670_ _01672_ _01674_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__o21ai_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _07841_ _07852_ _07857_ net7850 vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__a211oi_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ net3661 _05108_ _05152_ net4160 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ net80 _06734_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__or2_1
X_10915_ net6237 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
X_17471_ _01711_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__nor2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14683_ _07784_ _07786_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ net4057 _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19210_ net5165 _03182_ _03193_ _03189_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__o211a_1
X_16422_ _09511_ _09512_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__xnor2_1
X_13634_ _06801_ _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__and2_1
X_10846_ net6223 net7049 _04238_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20539__277 clknet_1_1__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__inv_2
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ _09443_ _09444_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__and2b_1
X_19141_ net1637 _03147_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__or2_1
X_13565_ _06681_ _06727_ _06663_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__or3b_4
XFILLER_0_82_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ net2177 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ _08397_ _08398_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19072_ net3852 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__clkbuf_1
X_12516_ net11 _05691_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__nand2_1
X_16284_ _09373_ _09250_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13496_ _06620_ _06627_ _06557_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15235_ _08322_ _08329_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__nor2_1
X_18023_ _02220_ _02221_ _02228_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__o21a_1
X_12447_ _05630_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15166_ net3457 _08236_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__or2_1
X_12378_ _05517_ _05560_ _05562_ _05465_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__o211a_1
X_14117_ _07254_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__inv_2
X_11329_ rbzero.texu_hot\[2\] _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19974_ net1867 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
X_15097_ net7776 _08190_ _08191_ _08124_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__o211a_1
X_14048_ _07210_ _07218_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__xor2_1
X_18925_ net6436 net3407 _03025_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18856_ net3329 net4591 _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17807_ _01855_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__xnor2_1
X_18787_ _02866_ net4838 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__nand2_1
X_15999_ _08983_ _08985_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__xor2_4
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17738_ _01975_ _01976_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__nor2_1
X_17669_ _01794_ _09403_ _01793_ _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__o31a_1
X_19408_ net2146 _03303_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7304 net4400 vssd1 vssd1 vccd1 vccd1 net7831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7315 _06551_ vssd1 vssd1 vccd1 vccd1 net7842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7326 net3450 vssd1 vssd1 vccd1 vccd1 net7853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6603 rbzero.tex_g0\[59\] vssd1 vssd1 vccd1 vccd1 net7130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7348 net4521 vssd1 vssd1 vccd1 vccd1 net7875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6614 net2384 vssd1 vssd1 vccd1 vccd1 net7141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7359 net950 vssd1 vssd1 vccd1 vccd1 net7886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6625 rbzero.tex_g1\[26\] vssd1 vssd1 vccd1 vccd1 net7152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21301_ clknet_leaf_43_i_clk net5187 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6636 net2012 vssd1 vssd1 vccd1 vccd1 net7163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6647 rbzero.pov.spi_buffer\[65\] vssd1 vssd1 vccd1 vccd1 net7174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5902 net8276 vssd1 vssd1 vccd1 vccd1 net6429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6658 rbzero.tex_g0\[54\] vssd1 vssd1 vccd1 vccd1 net7185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5913 net1346 vssd1 vssd1 vccd1 vccd1 net6440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6669 net2554 vssd1 vssd1 vccd1 vccd1 net7196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5924 _03820_ vssd1 vssd1 vccd1 vccd1 net6451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5935 net1198 vssd1 vssd1 vccd1 vccd1 net6462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold210 _01106_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
X_21232_ clknet_leaf_123_i_clk net3347 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold221 net5020 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5946 rbzero.spi_registers.new_texadd\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net6473
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 net5261 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5957 net1462 vssd1 vssd1 vccd1 vccd1 net6484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 net5114 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5968 rbzero.spi_registers.new_texadd\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net6495
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5979 net1269 vssd1 vssd1 vccd1 vccd1 net6506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 net4851 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ clknet_leaf_134_i_clk net1864 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold265 net4605 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 net6091 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold287 net5303 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
X_20114_ net3469 _03698_ _03615_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__o21ai_1
Xhold298 net5213 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21094_ clknet_leaf_12_i_clk net1516 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20045_ net3682 _03646_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__or2_1
X_20644__372 clknet_1_1__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__inv_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20343__100 clknet_1_0__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__inv_2
XFILLER_0_147_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21996_ net438 net1091 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20947_ clknet_leaf_77_i_clk net4334 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ net5688 net5544 _04160_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__mux2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04857_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
X_20878_ _09739_ _02756_ net4600 _02508_ net8100 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ net6172 net2993 _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13350_ _06471_ _06520_ _06466_ _06469_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__o211a_1
X_10562_ net6144 net6195 _04086_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _05239_ vssd1 vssd1 vccd1 vccd1 _05487_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13281_ _06385_ _06352_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__or2_2
X_10493_ net7161 net7165 _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7882 _08151_ vssd1 vssd1 vccd1 vccd1 net8409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7893 _08435_ vssd1 vssd1 vccd1 vccd1 net8420 sky130_fd_sc_hd__dlygate4sd3_1
X_15020_ _08114_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__buf_4
X_12232_ _04949_ _05416_ _05418_ _05213_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12163_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _05237_ vssd1 vssd1 vccd1 vccd1 _05351_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ net2537 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
X_16971_ _09653_ _09695_ _09992_ vssd1 vssd1 vccd1 vccd1 _09993_ sky130_fd_sc_hd__a21oi_2
X_12094_ _04991_ _05273_ _05282_ _04821_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18710_ _09747_ net4798 _02862_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__or3_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ net7041 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
X_15922_ _08415_ _08419_ _08412_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__a21bo_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ net6484 net3562 _03468_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ net5805 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__clkbuf_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _08401_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__clkbuf_4
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14804_ _07818_ _07804_ _07875_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__a21o_1
XFILLER_0_207_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18572_ _09756_ _09759_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__xnor2_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _08869_ _08870_ _08871_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__o21ai_2
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ net3932 vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _10163_ _09060_ _01762_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__o21ai_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ net4399 _07903_ _07872_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ net3719 _05103_ _05093_ rbzero.debug_overlay.facingX\[0\] vssd1 vssd1 vccd1
+ vccd1 _05136_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17454_ _10106_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14666_ _07832_ _07834_ _07836_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__a21o_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ net5205 net5911 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16405_ _09477_ _09495_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__xor2_2
X_13617_ _06776_ _06787_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__xnor2_1
X_10829_ net3249 net6211 _04227_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17385_ _10400_ _10401_ vssd1 vssd1 vccd1 vccd1 _10403_ sky130_fd_sc_hd__and2_1
X_14597_ _07737_ _07762_ _07765_ _07766_ _07767_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ net6816 net3375 _03139_ net4451 _08093_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__o311a_1
X_16336_ _09291_ _09302_ _09427_ vssd1 vssd1 vccd1 vccd1 _09428_ sky130_fd_sc_hd__a21bo_1
X_13548_ _06662_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16267_ _09357_ _09358_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__xnor2_1
X_19055_ net3867 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13479_ _06648_ _06649_ _06538_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5209 rbzero.pov.ready_buffer\[56\] vssd1 vssd1 vccd1 vccd1 net5736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15218_ _06010_ _06349_ _04510_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__mux2_1
X_18006_ _02055_ _02058_ _02056_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a21bo_1
X_16198_ _09286_ _09290_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4508 net667 vssd1 vssd1 vccd1 vccd1 net5035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4519 _01240_ vssd1 vssd1 vccd1 vccd1 net5046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _08220_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3807 net1793 vssd1 vssd1 vccd1 vccd1 net4334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3818 _01186_ vssd1 vssd1 vccd1 vccd1 net4345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3829 net1291 vssd1 vssd1 vccd1 vccd1 net4356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19957_ net7175 net5812 _03583_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18908_ net6649 net6954 _03014_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
X_19888_ net3256 net6436 _03550_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18839_ _02968_ _02978_ _02980_ net5864 net3935 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a32o_1
XFILLER_0_207_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21850_ net292 net2287 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20801_ _03878_ _03967_ net8229 _03883_ net5522 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21781_ clknet_leaf_9_i_clk net1357 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_20732_ net1106 net5340 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7101 rbzero.spi_registers.spi_buffer\[18\] vssd1 vssd1 vccd1 vccd1 net7628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7112 _03729_ vssd1 vssd1 vccd1 vccd1 net7639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7123 _03501_ vssd1 vssd1 vccd1 vccd1 net7650 sky130_fd_sc_hd__dlygate4sd3_1
X_20594_ clknet_1_1__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6400 rbzero.tex_r1\[3\] vssd1 vssd1 vccd1 vccd1 net6927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7145 rbzero.pov.spi_counter\[3\] vssd1 vssd1 vccd1 vccd1 net7672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6411 net2447 vssd1 vssd1 vccd1 vccd1 net6938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7156 net3971 vssd1 vssd1 vccd1 vccd1 net7683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6422 _04363_ vssd1 vssd1 vccd1 vccd1 net6949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7167 rbzero.spi_registers.spi_counter\[3\] vssd1 vssd1 vccd1 vccd1 net7694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6433 net2223 vssd1 vssd1 vccd1 vccd1 net6960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7178 net3682 vssd1 vssd1 vccd1 vccd1 net7705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6444 net1944 vssd1 vssd1 vccd1 vccd1 net6971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5710 net1140 vssd1 vssd1 vccd1 vccd1 net6237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7189 net4091 vssd1 vssd1 vccd1 vccd1 net7716 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold6455 rbzero.tex_r0\[59\] vssd1 vssd1 vccd1 vccd1 net6982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5721 rbzero.tex_b1\[52\] vssd1 vssd1 vccd1 vccd1 net6248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6466 net2409 vssd1 vssd1 vccd1 vccd1 net6993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6477 rbzero.tex_g1\[10\] vssd1 vssd1 vccd1 vccd1 net7004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5732 net1235 vssd1 vssd1 vccd1 vccd1 net6259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5743 rbzero.tex_b1\[12\] vssd1 vssd1 vccd1 vccd1 net6270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6488 net2288 vssd1 vssd1 vccd1 vccd1 net7015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6499 _04416_ vssd1 vssd1 vccd1 vccd1 net7026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5754 net1278 vssd1 vssd1 vccd1 vccd1 net6281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5765 rbzero.tex_g1\[0\] vssd1 vssd1 vccd1 vccd1 net6292 sky130_fd_sc_hd__dlygate4sd3_1
X_21215_ clknet_leaf_120_i_clk net2831 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5776 net1329 vssd1 vssd1 vccd1 vccd1 net6303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5787 rbzero.spi_registers.new_texadd\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 net6314
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5798 net1349 vssd1 vssd1 vccd1 vccd1 net6325 sky130_fd_sc_hd__dlygate4sd3_1
X_21146_ clknet_leaf_103_i_clk net3465 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_21077_ clknet_leaf_71_i_clk _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20028_ net5868 _03631_ _03606_ _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12850_ _05989_ _05995_ _06021_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or4b_1
XFILLER_0_198_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04844_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__clkbuf_8
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nand2_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21979_ net421 net2228 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _07624_ _07649_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__xor2_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__buf_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _07617_ _07620_ _07621_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _04847_ _04848_ _04849_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or4_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13402_ _06493_ _06572_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__nor2_1
X_10614_ net7403 net7200 _04116_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__mux2_1
X_17170_ _08374_ vssd1 vssd1 vccd1 vccd1 _10190_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14382_ _07532_ _07552_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__xor2_4
X_11594_ net1023 net4312 vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _09212_ _09213_ net7779 vssd1 vssd1 vccd1 vccd1 _09215_ sky130_fd_sc_hd__o21ai_1
X_13333_ _06407_ _06467_ _06478_ _06433_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and4b_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ net2641 net6715 _04075_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _09144_ _09145_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13264_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__buf_6
Xhold7690 net5779 vssd1 vssd1 vccd1 vccd1 net8217 sky130_fd_sc_hd__clkbuf_4
X_10476_ net6952 net7123 _04042_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_1
X_15003_ net740 _08100_ net3985 vssd1 vssd1 vccd1 vccd1 _08101_ sky130_fd_sc_hd__mux2_1
X_12215_ _04943_ _05399_ _05401_ _04928_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__o211a_1
X_13195_ _06356_ _06357_ _06361_ net8217 _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19811_ clknet_1_1__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__buf_1
XFILLER_0_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _05220_ vssd1 vssd1 vccd1 vccd1 _05334_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19742_ net4944 net7656 _03505_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__a21oi_1
X_12077_ rbzero.tex_r1\[51\] rbzero.tex_r1\[50\] _04979_ vssd1 vssd1 vccd1 vccd1 _05266_
+ sky130_fd_sc_hd__mux2_1
X_16954_ _09974_ _09975_ vssd1 vssd1 vccd1 vccd1 _09976_ sky130_fd_sc_hd__and2_2
XFILLER_0_194_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11028_ net5671 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
X_15905_ _08543_ _08535_ _08998_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__o21ai_1
X_19673_ net6419 net2205 _03457_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16885_ _09905_ _09906_ vssd1 vssd1 vccd1 vccd1 _09907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_159_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ net4686 rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02783_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15836_ _08888_ _08930_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__and2_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18555_ _06057_ _06050_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__nor2_1
X_15767_ _08838_ _08840_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__xor2_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ net4306 net4044 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__xnor2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17506_ _09915_ _09225_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14718_ _07818_ _07863_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__nand2_1
X_18486_ _02536_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__buf_4
X_20396__148 clknet_1_1__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__inv_2
X_15698_ _08787_ _08792_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17437_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ net7811 _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_16 _09735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net4173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _10262_ _10264_ vssd1 vssd1 vccd1 vccd1 _10386_ sky130_fd_sc_hd__nor2_1
XANTENNA_49 _04021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19107_ net5570 _03126_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__or2_1
X_16319_ net4624 _06123_ _09410_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17299_ _10187_ _10317_ vssd1 vssd1 vccd1 vccd1 _10318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5006 net1612 vssd1 vssd1 vccd1 vccd1 net5533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5017 rbzero.tex_r0\[10\] vssd1 vssd1 vccd1 vccd1 net5544 sky130_fd_sc_hd__dlygate4sd3_1
X_19038_ net3838 net3745 net3398 vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5028 _00523_ vssd1 vssd1 vccd1 vccd1 net5555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5039 rbzero.tex_b0\[1\] vssd1 vssd1 vccd1 vccd1 net5566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4305 net3083 vssd1 vssd1 vccd1 vccd1 net4832 sky130_fd_sc_hd__buf_1
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4316 _03425_ vssd1 vssd1 vccd1 vccd1 net4843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4327 net782 vssd1 vssd1 vccd1 vccd1 net4854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4338 _06056_ vssd1 vssd1 vccd1 vccd1 net4865 sky130_fd_sc_hd__clkbuf_2
Xhold3604 gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 net4131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3615 _08096_ vssd1 vssd1 vccd1 vccd1 net4142 sky130_fd_sc_hd__dlygate4sd3_1
X_21000_ clknet_leaf_83_i_clk _00487_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3626 _04717_ vssd1 vssd1 vccd1 vccd1 net4153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3637 _05546_ vssd1 vssd1 vccd1 vccd1 net4164 sky130_fd_sc_hd__clkbuf_4
Xhold2903 net8374 vssd1 vssd1 vccd1 vccd1 net3430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3648 _00462_ vssd1 vssd1 vccd1 vccd1 net4175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2914 _03664_ vssd1 vssd1 vccd1 vccd1 net3441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3659 net3336 vssd1 vssd1 vccd1 vccd1 net4186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2925 _04654_ vssd1 vssd1 vccd1 vccd1 net3452 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1__f__03509_ clknet_0__03509_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03509_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2936 rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 net3715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2947 net4376 vssd1 vssd1 vccd1 vccd1 net3474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2958 net7693 vssd1 vssd1 vccd1 vccd1 net3485 sky130_fd_sc_hd__clkbuf_2
Xhold2969 _03761_ vssd1 vssd1 vccd1 vccd1 net3496 sky130_fd_sc_hd__dlygate4sd3_1
X_21902_ net344 net2902 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21833_ net275 net2939 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21764_ clknet_leaf_83_i_clk net4093 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20455__201 clknet_1_0__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__inv_2
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20715_ net960 net5380 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21695_ clknet_leaf_110_i_clk net3442 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6230 rbzero.tex_r1\[54\] vssd1 vssd1 vccd1 vccd1 net6757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6241 net1952 vssd1 vssd1 vccd1 vccd1 net6768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6252 rbzero.tex_b0\[15\] vssd1 vssd1 vccd1 vccd1 net6779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6263 net1983 vssd1 vssd1 vccd1 vccd1 net6790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6274 rbzero.tex_b0\[21\] vssd1 vssd1 vccd1 vccd1 net6801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6285 net1935 vssd1 vssd1 vccd1 vccd1 net6812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5540 rbzero.spi_registers.new_texadd\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net6067
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6296 _04133_ vssd1 vssd1 vccd1 vccd1 net6823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5551 net2415 vssd1 vssd1 vccd1 vccd1 net6078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5562 _04080_ vssd1 vssd1 vccd1 vccd1 net6089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5573 net1095 vssd1 vssd1 vccd1 vccd1 net6100 sky130_fd_sc_hd__dlygate4sd3_1
X_12000_ _05182_ _05187_ _05188_ _04702_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__or4b_2
Xhold5584 net1098 vssd1 vssd1 vccd1 vccd1 net6111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4850 _01608_ vssd1 vssd1 vccd1 vccd1 net5377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5595 net1092 vssd1 vssd1 vccd1 vccd1 net6122 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4861 net1011 vssd1 vssd1 vccd1 vccd1 net5388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4872 rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 net5399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4883 net895 vssd1 vssd1 vccd1 vccd1 net5410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4894 _00781_ vssd1 vssd1 vccd1 vccd1 net5421 sky130_fd_sc_hd__dlygate4sd3_1
X_21129_ clknet_leaf_32_i_clk net3809 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13951_ _06719_ _06698_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__or3_1
XFILLER_0_199_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12902_ net2277 net2058 net1006 net894 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__or4_1
X_13882_ _07049_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nor2_1
X_16670_ net4615 _09737_ _09740_ _07975_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15621_ _08220_ _08240_ _08279_ _08317_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ _06008_ _05953_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__xnor2_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _05155_ net3565 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _08350_ _08337_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__xnor2_4
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _05905_ _05940_ net37 vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_185_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11715_ _04844_ _04845_ _04853_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o31a_1
X_14503_ _07638_ _07637_ _07636_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15483_ _08570_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__xnor2_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18271_ net6335 net1493 _02477_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ net4133 net4089 _05851_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__mux2_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _10058_ _10118_ _10117_ vssd1 vssd1 vccd1 vccd1 _10242_ sky130_fd_sc_hd__a21oi_1
X_11646_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__buf_4
X_14434_ _07580_ _07603_ _07604_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_1_1__f__03860_ clknet_0__03860_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03860_
+ sky130_fd_sc_hd__clkbuf_16
Xinput14 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
X_17153_ _10162_ _10172_ vssd1 vssd1 vccd1 vccd1 _10173_ sky130_fd_sc_hd__xnor2_1
X_14365_ _07521_ _07527_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__xor2_4
Xinput25 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_4
Xinput36 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
X_11577_ net1101 net4230 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput47 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_4
X_16104_ _09195_ _09197_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13316_ _06424_ _06426_ _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__and3b_1
X_17084_ _08905_ net4877 _10104_ _09970_ vssd1 vssd1 vccd1 vccd1 _10105_ sky130_fd_sc_hd__or4_4
X_10528_ net7087 net7439 _04064_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14296_ _07464_ _07465_ _07466_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__nand3_1
Xhold809 _01004_ vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16035_ _09067_ _09128_ vssd1 vssd1 vccd1 vccd1 _09129_ sky130_fd_sc_hd__xnor2_1
X_13247_ _06387_ _06409_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__nor2_1
X_10459_ net2348 net6581 _04031_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13178_ _06339_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12129_ _04921_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__or2_1
X_17986_ _02132_ _02097_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__and2b_1
XFILLER_0_202_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1509 net6925 vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
X_19725_ _03489_ net3704 _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__and3b_1
X_16937_ _09957_ _09958_ vssd1 vssd1 vccd1 vccd1 _09959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19656_ net6621 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__clkbuf_1
X_16868_ _09611_ _09613_ _09609_ vssd1 vssd1 vccd1 vccd1 _09890_ sky130_fd_sc_hd__a21oi_1
X_18607_ _02767_ _08038_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__nor2_1
X_15819_ _08896_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__or2_1
X_19587_ net1393 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
X_16799_ _09826_ _09824_ net4631 _06057_ vssd1 vssd1 vccd1 vccd1 _09828_ sky130_fd_sc_hd__a31o_1
X_19745__27 clknet_1_1__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
XFILLER_0_88_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18538_ net3894 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18469_ _02617_ net4698 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21480_ clknet_leaf_16_i_clk net1379 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22101_ net163 net2121 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4102 net8350 vssd1 vssd1 vccd1 vccd1 net4629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4113 net744 vssd1 vssd1 vccd1 vccd1 net4640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4124 net3836 vssd1 vssd1 vccd1 vccd1 net4651 sky130_fd_sc_hd__clkbuf_2
X_20293_ net1460 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4135 _00433_ vssd1 vssd1 vccd1 vccd1 net4662 sky130_fd_sc_hd__dlygate4sd3_1
X_22032_ net474 net2678 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
Xhold4146 net3560 vssd1 vssd1 vccd1 vccd1 net4673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3401 _03746_ vssd1 vssd1 vccd1 vccd1 net3928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4157 _00420_ vssd1 vssd1 vccd1 vccd1 net4684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3412 rbzero.spi_registers.spi_cmd\[2\] vssd1 vssd1 vccd1 vccd1 net3939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3423 net2872 vssd1 vssd1 vccd1 vccd1 net3950 sky130_fd_sc_hd__clkbuf_2
Xhold4168 _08055_ vssd1 vssd1 vccd1 vccd1 net4695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3434 _02731_ vssd1 vssd1 vccd1 vccd1 net3961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4179 _08061_ vssd1 vssd1 vccd1 vccd1 net4706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2700 net1788 vssd1 vssd1 vccd1 vccd1 net3227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3445 _04472_ vssd1 vssd1 vccd1 vccd1 net3972 sky130_fd_sc_hd__clkbuf_1
Xhold2711 _03594_ vssd1 vssd1 vccd1 vccd1 net3238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3456 _04737_ vssd1 vssd1 vccd1 vccd1 net3983 sky130_fd_sc_hd__buf_1
Xhold2722 net7513 vssd1 vssd1 vccd1 vccd1 net3249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3467 _01177_ vssd1 vssd1 vccd1 vccd1 net3994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2733 net2330 vssd1 vssd1 vccd1 vccd1 net3260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3478 _01218_ vssd1 vssd1 vccd1 vccd1 net4005 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3489 net4039 vssd1 vssd1 vccd1 vccd1 net4016 sky130_fd_sc_hd__clkbuf_4
Xhold2744 _00709_ vssd1 vssd1 vccd1 vccd1 net3271 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2755 rbzero.pov.spi_buffer\[57\] vssd1 vssd1 vccd1 vccd1 net3282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2766 _03026_ vssd1 vssd1 vccd1 vccd1 net3293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2777 _01116_ vssd1 vssd1 vccd1 vccd1 net3304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2788 net5858 vssd1 vssd1 vccd1 vccd1 net3315 sky130_fd_sc_hd__clkbuf_2
Xhold2799 net7689 vssd1 vssd1 vccd1 vccd1 net3326 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21816_ net258 net1019 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21747_ clknet_leaf_98_i_clk net3622 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11500_ _04677_ _04681_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__and4b_1
XFILLER_0_109_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ net6 _05654_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21678_ clknet_leaf_124_i_clk net3222 vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11431_ rbzero.texu_hot\[0\] _04524_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14150_ _07312_ _07319_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ _04504_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__buf_4
Xhold6060 net1587 vssd1 vssd1 vccd1 vccd1 net6587 sky130_fd_sc_hd__dlygate4sd3_1
X_13101_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__and2_1
Xhold6071 rbzero.spi_registers.new_texadd\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net6598
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6082 net1756 vssd1 vssd1 vccd1 vccd1 net6609 sky130_fd_sc_hd__dlygate4sd3_1
X_14081_ _06577_ _06839_ _07251_ net5902 vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6093 _03453_ vssd1 vssd1 vccd1 vccd1 net6620 sky130_fd_sc_hd__dlygate4sd3_1
X_11293_ _04486_ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5370 rbzero.pov.ready_buffer\[71\] vssd1 vssd1 vccd1 vccd1 net5897 sky130_fd_sc_hd__dlygate4sd3_1
X_13032_ _06207_ net4526 _06201_ net3790 vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__a22o_1
Xhold5381 _03639_ vssd1 vssd1 vccd1 vccd1 net5908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5392 _00620_ vssd1 vssd1 vccd1 vccd1 net5919 sky130_fd_sc_hd__dlygate4sd3_1
X_17840_ _02076_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4680 _03790_ vssd1 vssd1 vccd1 vccd1 net5207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4691 net859 vssd1 vssd1 vccd1 vccd1 net5218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3990 net7935 vssd1 vssd1 vccd1 vccd1 net4517 sky130_fd_sc_hd__dlygate4sd3_1
X_17771_ _02008_ _02009_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__nor2_1
X_14983_ _08089_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
X_19510_ net2147 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
X_16722_ _09756_ _09759_ _09757_ vssd1 vssd1 vccd1 vccd1 _09760_ sky130_fd_sc_hd__a21o_1
X_13934_ _07104_ _06796_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19441_ _03320_ net3645 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__and2_1
X_16653_ net4089 net5949 _09732_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o21a_1
X_13865_ _06706_ _07035_ _06813_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15604_ _08339_ _08698_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__xnor2_4
X_19372_ net6470 _03284_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__or2_1
X_12816_ _05948_ _05976_ _05977_ _05991_ _05978_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a311oi_4
X_16584_ _08573_ _09673_ net4891 vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__a21o_1
X_13796_ _06964_ _06965_ _06966_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ net3565 net5033 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ net8041 _08124_ _08381_ _08382_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__or4_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ net35 net36 _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__and3_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18254_ net3591 _02467_ _02313_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__o21ai_1
X_15466_ _08550_ _08560_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12678_ _05851_ net4156 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17205_ _10222_ _10223_ _10221_ vssd1 vssd1 vccd1 vccd1 _10225_ sky130_fd_sc_hd__a21o_1
X_11629_ _04809_ _04808_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__and2b_1
X_14417_ _07566_ _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03843_ clknet_0__03843_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03843_
+ sky130_fd_sc_hd__clkbuf_16
X_18185_ net3766 net4481 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nand2_2
X_15397_ net8041 _06120_ _08491_ _08408_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__or4b_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17136_ _08542_ _09612_ _10032_ _10031_ vssd1 vssd1 vccd1 vccd1 _10156_ sky130_fd_sc_hd__o31a_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14348_ _07514_ _07517_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__a21o_1
Xhold606 net6857 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 _01523_ vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 net4260 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ _10086_ _10087_ vssd1 vssd1 vccd1 vccd1 _10088_ sky130_fd_sc_hd__nand2_1
Xhold639 net6240 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ _07334_ _07382_ _07380_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16018_ _08543_ _08614_ _09063_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__o21ai_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _04203_ vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2018 net7337 vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _01319_ vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 net6650 vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 _01529_ vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1328 _01504_ vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__xnor2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1339 net1808 vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
X_19708_ net6132 net3583 _03456_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_100_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20980_ clknet_leaf_58_i_clk _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_19639_ net6388 net3562 _03441_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21601_ clknet_leaf_130_i_clk net3232 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_115_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21532_ clknet_leaf_130_i_clk net3924 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20336__94 clknet_1_0__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__inv_2
XFILLER_0_209_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21463_ clknet_leaf_42_i_clk net2207 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21394_ clknet_leaf_39_i_clk net5486 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20567__302 clknet_1_1__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__inv_2
XFILLER_0_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20276_ net4092 _03806_ _03809_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3220 _00732_ vssd1 vssd1 vccd1 vccd1 net3747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22015_ net457 net1835 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
Xhold3242 rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 net3769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3253 _00611_ vssd1 vssd1 vccd1 vccd1 net3780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3264 net7960 vssd1 vssd1 vccd1 vccd1 net3791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2530 _03017_ vssd1 vssd1 vccd1 vccd1 net3057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3275 net7967 vssd1 vssd1 vccd1 vccd1 net3802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2541 _04033_ vssd1 vssd1 vccd1 vccd1 net3068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3286 net5873 vssd1 vssd1 vccd1 vccd1 net3813 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3297 _03503_ vssd1 vssd1 vccd1 vccd1 net3824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2552 _01102_ vssd1 vssd1 vccd1 vccd1 net3079 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2563 net7434 vssd1 vssd1 vccd1 vccd1 net3090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03863_ clknet_0__03863_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03863_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2574 net3110 vssd1 vssd1 vccd1 vccd1 net3101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1840 net7406 vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2585 _03005_ vssd1 vssd1 vccd1 vccd1 net3112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1851 _01449_ vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2596 _01141_ vssd1 vssd1 vccd1 vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ _04670_ _04658_ _05159_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a22o_1
Xhold1862 _01073_ vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1873 _04241_ vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 net7366 vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1895 _01400_ vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_10931_ net3247 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ net6587 net2826 _04171_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__mux2_1
X_13650_ _06810_ _06820_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12601_ _05760_ _05778_ _05779_ _05780_ net21 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_184_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13581_ _06712_ _06750_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ net7001 net6991 _04205_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ _08401_ _08411_ _08180_ _08414_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12532_ net14 net15 vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nor2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ _08306_ _08328_ _08343_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__or3_1
X_12463_ clknet_4_8__leaf_i_clk vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__buf_1
X_14202_ _07344_ _07343_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__and2b_1
X_11414_ _04584_ _04543_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15182_ _08117_ _08275_ _08276_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__a21oi_4
X_12394_ _05577_ _05578_ _05276_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14133_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11345_ _04519_ _04534_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a21o_1
X_19990_ net40 _03605_ _03122_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18941_ net2585 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
X_14064_ _06696_ _07194_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11276_ _04471_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_8
XFILLER_0_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ net4723 vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__inv_2
X_18872_ net3019 net7490 _02993_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _01979_ _01980_ _01977_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17754_ _01991_ _01992_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14966_ net4373 _07981_ _08079_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16705_ net8067 _09745_ _09746_ net7837 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a22o_1
X_13917_ _07067_ _07069_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__nor2_1
X_17685_ _01918_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14897_ net4569 _08034_ _08036_ net3787 net4744 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_i_clk clknet_4_10__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19424_ net5049 _03310_ _03319_ _03316_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__a211o_1
X_16636_ net3859 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__clkbuf_1
X_13848_ _06974_ _07007_ _07017_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19355_ net6283 _03271_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16567_ _08391_ _09165_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__or2_1
X_13779_ _06902_ _06904_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ net6605 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__clkbuf_1
X_15518_ _06121_ _08612_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19286_ net5129 _03236_ _03239_ _03230_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__o211a_1
X_16498_ _09461_ _09575_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7508 _06092_ vssd1 vssd1 vccd1 vccd1 net8035 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_47_i_clk clknet_4_8__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18237_ _02442_ _02445_ _02443_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__o21ai_1
X_15449_ _08338_ _08542_ _08543_ _08142_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_170_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6807 net816 vssd1 vssd1 vccd1 vccd1 net7334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6818 rbzero.tex_b1\[38\] vssd1 vssd1 vccd1 vccd1 net7345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6829 _04256_ vssd1 vssd1 vccd1 vccd1 net7356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18168_ net4782 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold403 net5365 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold414 net7882 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ _10136_ _10137_ _10013_ _10138_ vssd1 vssd1 vccd1 vccd1 _10139_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03857_ _03857_ vssd1 vssd1 vccd1 vccd1 clknet_0__03857_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold425 net5393 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _02328_ _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__xnor2_1
Xhold436 net5325 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold447 net5281 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 net8031 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20130_ net4462 _03711_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__or2_1
Xhold469 net5397 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20061_ net3440 _03485_ _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__a211o_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _00975_ vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _03375_ vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 net6642 vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1136 net7954 vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 rbzero.row_render.size\[8\] vssd1 vssd1 vccd1 vccd1 net3686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 net6569 vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _00993_ vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ clknet_leaf_77_i_clk _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ net4936 net63 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21515_ clknet_leaf_8_i_clk net1455 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21446_ clknet_leaf_19_i_clk net2955 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21377_ clknet_leaf_12_i_clk net5290 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ net2083 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20328_ net6082 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold970 net6423 vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 net6404 vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net2632 net5589 _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
Xhold992 _01507_ vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
X_20259_ net4111 _09733_ _03797_ _03794_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__a22o_1
Xhold3050 _03774_ vssd1 vssd1 vccd1 vccd1 net3577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3061 _02458_ vssd1 vssd1 vccd1 vccd1 net3588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3072 net7827 vssd1 vssd1 vccd1 vccd1 net3599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3083 _01203_ vssd1 vssd1 vccd1 vccd1 net3610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3094 _03772_ vssd1 vssd1 vccd1 vccd1 net3621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2360 net7356 vssd1 vssd1 vccd1 vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2371 net8192 vssd1 vssd1 vccd1 vccd1 net2898 sky130_fd_sc_hd__buf_2
X_14820_ net8354 _07910_ _07915_ net7793 net3638 vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_192_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2382 _01469_ vssd1 vssd1 vccd1 vccd1 net2909 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2393 net3055 vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03846_ clknet_0__03846_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03846_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20621__351 clknet_1_1__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__inv_2
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1670 net4696 vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1681 net7156 vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751_ _07918_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__clkbuf_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1692 _01366_ vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11963_ net3565 _05106_ _05114_ net3509 vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a22o_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06705_ _06808_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__nor2_2
X_17470_ _01709_ _01710_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__and2_1
X_10914_ net6235 net2604 _04276_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _07510_ _07787_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__xnor2_1
X_11894_ net3919 _05071_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _09262_ _08392_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__nor2_1
X_10845_ net2024 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13633_ _06802_ _06775_ _06803_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19140_ net5505 _03145_ net1134 _03149_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16352_ _09440_ _09442_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10776_ net6114 net7105 _04194_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__mux2_1
X_13564_ _06719_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15303_ _08377_ _08388_ _08396_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__nand3_1
XFILLER_0_165_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19071_ net5895 net3940 _03104_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
X_12515_ net15 _05695_ net11 net12 vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__and4b_1
X_16283_ _09135_ _09249_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__nand2_1
X_13495_ _06547_ _06664_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ _02256_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__xnor2_1
X_15234_ _08328_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__clkbuf_4
X_12446_ reg_vsync _04477_ _05054_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__mux2_4
XFILLER_0_180_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12377_ _04922_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15165_ net4293 _08259_ _08124_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14116_ _06577_ _07251_ net542 _07104_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__a211o_1
X_11328_ rbzero.spi_registers.texadd3\[8\] rbzero.spi_registers.texadd1\[8\] rbzero.spi_registers.texadd0\[8\]
+ rbzero.spi_registers.texadd2\[8\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux4_2
X_19973_ net54 net1866 _03109_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__mux2_1
X_15096_ net3372 _06033_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18924_ net3081 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
X_11259_ net5566 net1836 _04104_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__mux2_1
X_14047_ _07216_ _07217_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18855_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__clkbuf_4
X_17806_ _02043_ _02044_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18786_ _02866_ net4838 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15998_ _09091_ net8542 vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__and2_1
X_19787__66 clknet_1_1__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
XFILLER_0_206_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17737_ _10190_ _09225_ _01748_ _01863_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__o31a_1
XFILLER_0_171_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ net4485 _07917_ _08068_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17668_ _01791_ _01792_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__nand2_1
X_19407_ net5518 _03302_ _03308_ _03299_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16619_ _09707_ _09708_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__or2_1
X_17599_ _01737_ _01738_ _01838_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19338_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7305 net4718 vssd1 vssd1 vccd1 vccd1 net7832 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7316 _07840_ vssd1 vssd1 vccd1 vccd1 net7843 sky130_fd_sc_hd__buf_2
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7327 rbzero.traced_texVinit\[8\] vssd1 vssd1 vccd1 vccd1 net7854 sky130_fd_sc_hd__dlygate4sd3_1
X_19269_ net6562 _03217_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6604 net2420 vssd1 vssd1 vccd1 vccd1 net7131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7349 rbzero.wall_tracer.stepDistY\[-10\] vssd1 vssd1 vccd1 vccd1 net7876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21300_ clknet_leaf_44_i_clk net5083 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6615 rbzero.pov.ready_buffer\[26\] vssd1 vssd1 vccd1 vccd1 net7142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6626 net2515 vssd1 vssd1 vccd1 vccd1 net7153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6637 rbzero.tex_r1\[44\] vssd1 vssd1 vccd1 vccd1 net7164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6648 net2190 vssd1 vssd1 vccd1 vccd1 net7175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5903 net1432 vssd1 vssd1 vccd1 vccd1 net6430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5914 rbzero.tex_b1\[44\] vssd1 vssd1 vccd1 vccd1 net6441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6659 net2691 vssd1 vssd1 vccd1 vccd1 net7186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21231_ clknet_leaf_125_i_clk net3017 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold200 net5008 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5925 net1466 vssd1 vssd1 vccd1 vccd1 net6452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold211 net5140 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5936 rbzero.spi_registers.new_mapd\[11\] vssd1 vssd1 vccd1 vccd1 net6463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold222 net5022 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5947 net1307 vssd1 vssd1 vccd1 vccd1 net6474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5958 rbzero.spi_registers.new_other\[3\] vssd1 vssd1 vccd1 vccd1 net6485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 net5116 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 net5144 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ clknet_leaf_130_i_clk net2766 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold255 net4853 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5969 net1576 vssd1 vssd1 vccd1 vccd1 net6496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 net5160 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 net6093 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20113_ _03352_ net6063 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__nor2_1
Xhold288 net5305 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 net5060 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
X_21093_ clknet_leaf_12_i_clk net1510 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20044_ net3431 _03609_ net5899 _03316_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a211o_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ net437 net3358 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ clknet_leaf_69_i_clk net4663 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _02753_ net4599 net4424 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a21bo_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ _04104_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10561_ net2272 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _04913_ vssd1 vssd1 vccd1 vccd1 _05486_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13280_ net8217 _06329_ _06332_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o21ai_2
Xhold7850 _06016_ vssd1 vssd1 vccd1 vccd1 net8377 sky130_fd_sc_hd__dlygate4sd3_1
X_10492_ _04030_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__clkbuf_4
Xhold7872 _08431_ vssd1 vssd1 vccd1 vccd1 net8399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ _04847_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__or2_1
Xhold7883 _08152_ vssd1 vssd1 vccd1 vccd1 net8410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21429_ clknet_leaf_36_i_clk net1563 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12162_ _04942_ _05337_ _05341_ _05349_ _04817_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__o311a_1
XFILLER_0_124_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11113_ net6052 net6890 _04375_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux2_1
X_16970_ _09692_ _09694_ vssd1 vssd1 vccd1 vccd1 _09992_ sky130_fd_sc_hd__nor2_1
X_12093_ _05275_ _05278_ _05281_ _05213_ _04825_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ net2333 net7039 _04342_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15921_ _08393_ _08395_ _08390_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__a21bo_1
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18640_ rbzero.wall_tracer.rayAddendY\[-2\] _02797_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _08691_ _08329_ net8423 net7836 vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__and4bb_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 _01349_ vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _07881_ _07884_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ net4035 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _08876_ _08877_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__nor2_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ net4500 _06169_ net4508 _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__o22a_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17522_ _10163_ _09060_ _01762_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__or3_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14734_ _07869_ _07902_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__or2b_2
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11946_ _05116_ _05131_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__or3b_4
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17453_ _09537_ _01694_ _10350_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14665_ _07825_ _07835_ _07439_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__and3b_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _05060_ _05063_ net3919 net4057 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16404_ _09493_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__nor2_1
X_13616_ _06777_ _06785_ _06786_ _06779_ _06784_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__o32a_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ net2030 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__clkbuf_1
X_17384_ _10400_ _10401_ vssd1 vssd1 vccd1 vccd1 _10402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14596_ _07710_ _07718_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ net3374 _03141_ net4450 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a21o_1
X_16335_ _09301_ _09299_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__or2b_1
X_13547_ _06713_ _06717_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__xnor2_1
X_10759_ net6205 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__clkbuf_1
X_19054_ net7629 net7585 net3398 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
X_16266_ _08543_ _09116_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__nor2_1
X_13478_ _06491_ _06584_ _06585_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18005_ _02240_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15217_ net5902 _06502_ _07902_ _08113_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__a31o_1
X_12429_ _05608_ _05610_ _05613_ _05233_ _04967_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16197_ _09287_ _09289_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4509 rbzero.spi_registers.texadd1\[21\] vssd1 vssd1 vccd1 vccd1 net5036 sky130_fd_sc_hd__dlygate4sd3_1
X_15148_ _08204_ _08205_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3808 net8153 vssd1 vssd1 vccd1 vccd1 net4335 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3819 net3416 vssd1 vssd1 vccd1 vccd1 net4346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20628__357 clknet_1_0__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__inv_2
X_19956_ net2928 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
X_15079_ net4277 _08117_ _08148_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__a21o_1
XFILLER_0_208_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18907_ net3290 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
X_19887_ net3257 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18838_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18769_ net3761 _09736_ _02917_ _04490_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20800_ _03965_ _03966_ _03964_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21780_ clknet_leaf_3_i_clk net1504 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20731_ _03904_ _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7102 net3866 vssd1 vssd1 vccd1 vccd1 net7629 sky130_fd_sc_hd__dlygate4sd3_1
X_20373__127 clknet_1_0__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__inv_2
Xhold7113 net3687 vssd1 vssd1 vccd1 vccd1 net7640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7135 _03718_ vssd1 vssd1 vccd1 vccd1 net7662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6401 net1958 vssd1 vssd1 vccd1 vccd1 net6928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7146 net3707 vssd1 vssd1 vccd1 vccd1 net7673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6412 rbzero.tex_r1\[61\] vssd1 vssd1 vccd1 vccd1 net6939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7157 rbzero.pov.spi_counter\[1\] vssd1 vssd1 vccd1 vccd1 net7684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6423 net2275 vssd1 vssd1 vccd1 vccd1 net6950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7168 _02966_ vssd1 vssd1 vccd1 vccd1 net7695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6434 _03394_ vssd1 vssd1 vccd1 vccd1 net6961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7179 _02745_ vssd1 vssd1 vccd1 vccd1 net7706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6445 rbzero.tex_b0\[59\] vssd1 vssd1 vccd1 vccd1 net6972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5700 net1188 vssd1 vssd1 vccd1 vccd1 net6227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6456 net2530 vssd1 vssd1 vccd1 vccd1 net6983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5711 net6579 vssd1 vssd1 vccd1 vccd1 net6238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6467 rbzero.tex_b0\[53\] vssd1 vssd1 vccd1 vccd1 net6994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5722 net1158 vssd1 vssd1 vccd1 vccd1 net6249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5733 _04063_ vssd1 vssd1 vccd1 vccd1 net6260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6478 net2738 vssd1 vssd1 vccd1 vccd1 net7005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6489 rbzero.tex_r0\[34\] vssd1 vssd1 vccd1 vccd1 net7016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5744 net1225 vssd1 vssd1 vccd1 vccd1 net6271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21214_ clknet_leaf_120_i_clk net1560 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5755 rbzero.spi_registers.new_texadd\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net6282
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5766 net1596 vssd1 vssd1 vccd1 vccd1 net6293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5777 rbzero.spi_registers.new_texadd\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 net6304
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5788 net1468 vssd1 vssd1 vccd1 vccd1 net6315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5799 rbzero.pov.spi_buffer\[71\] vssd1 vssd1 vccd1 vccd1 net6326 sky130_fd_sc_hd__dlygate4sd3_1
X_21145_ clknet_leaf_104_i_clk net4801 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_21076_ clknet_leaf_76_i_clk _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20027_ net3443 _08295_ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _04983_ _04989_ _04825_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__o21a_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _05952_
+ _05955_ _05950_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a221oi_4
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ net420 net2051 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _04832_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__buf_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20929_ clknet_leaf_60_i_clk net4746 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _07616_ _07615_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__and2b_1
X_11662_ net87 net88 net85 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13401_ _06467_ _06432_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__mux2_1
X_10613_ net7011 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11593_ _04779_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14381_ _07534_ _07550_ _07551_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_92_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ net7779 _09212_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__or3_1
X_10544_ net6090 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__clkbuf_1
X_13332_ _06495_ net554 vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__nand2_4
XFILLER_0_84_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16051_ _08229_ _08323_ _09004_ _09002_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7680 net3433 vssd1 vssd1 vccd1 vccd1 net8207 sky130_fd_sc_hd__dlymetal6s2s_1
X_10475_ net2781 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13263_ _06389_ _06407_ _06413_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__or4bb_4
Xhold7691 _00000_ vssd1 vssd1 vccd1 vccd1 net8218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _06145_ _08099_ net1013 _06102_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__a2bb2o_1
X_12214_ _04930_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__or2_1
Xhold6990 rbzero.tex_r0\[13\] vssd1 vssd1 vccd1 vccd1 net7517 sky130_fd_sc_hd__dlygate4sd3_1
X_13194_ _06362_ _06363_ _06364_ _04491_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a22o_2
X_12145_ _04818_ _05307_ _05315_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__a31o_1
X_19810_ clknet_1_0__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__buf_1
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ _04967_ _05248_ _05254_ _04818_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__o311a_1
X_19741_ net4944 net7656 _03493_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__o21ai_1
X_16953_ net4388 _06124_ vssd1 vssd1 vccd1 vccd1 _09975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ net2735 net5669 _04331_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15904_ _08529_ _08535_ _08998_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19672_ net1347 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__clkbuf_1
X_16884_ _08127_ net7818 vssd1 vssd1 vccd1 vccd1 _09906_ sky130_fd_sc_hd__and2_1
XFILLER_0_188_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18623_ net4686 rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02782_
+ sky130_fd_sc_hd__nor2_1
X_15835_ _08886_ _08887_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__nand2_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18554_ _06049_ _06034_ _06047_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__or3_1
X_15766_ _08833_ _08842_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__xnor2_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ net4315 _06062_ _06048_ net1803 _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__o221a_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _08167_ net4914 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__nand2_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ _07821_ _07861_ _07886_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__a21oi_1
X_18485_ _02654_ _02655_ _02662_ _02526_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a2bb2o_1
X_11929_ net3536 _05113_ _05114_ net3339 _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15697_ _08790_ _08791_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__nand2_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ _10430_ _10431_ _01676_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nand3_1
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14648_ _07804_ _07817_ _07818_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _10009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _10383_ _10384_ vssd1 vssd1 vccd1 vccd1 _10385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_39 net4490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ _07739_ _07749_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19106_ net4347 _03125_ net890 _03128_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__o211a_1
X_16318_ _09409_ _09174_ _06122_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__a21o_2
X_17298_ _08338_ _10316_ vssd1 vssd1 vccd1 vccd1 _10317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19037_ net3839 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__clkbuf_1
Xhold5007 rbzero.spi_registers.new_other\[4\] vssd1 vssd1 vccd1 vccd1 net5534 sky130_fd_sc_hd__dlygate4sd3_1
X_16249_ _09270_ _09246_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5018 _04165_ vssd1 vssd1 vccd1 vccd1 net5545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5029 net2007 vssd1 vssd1 vccd1 vccd1 net5556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4306 _02472_ vssd1 vssd1 vccd1 vccd1 net4833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4317 net1044 vssd1 vssd1 vccd1 vccd1 net4844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3605 net4120 vssd1 vssd1 vccd1 vccd1 net4132 sky130_fd_sc_hd__buf_4
Xhold3616 _00460_ vssd1 vssd1 vccd1 vccd1 net4143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3627 _04726_ vssd1 vssd1 vccd1 vccd1 net4154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3638 _08097_ vssd1 vssd1 vccd1 vccd1 net4165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2904 net7700 vssd1 vssd1 vccd1 vccd1 net3431 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3649 gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 net4176 sky130_fd_sc_hd__buf_2
Xclkbuf_1_1__f__03508_ clknet_0__03508_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03508_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2915 net5930 vssd1 vssd1 vccd1 vccd1 net3442 sky130_fd_sc_hd__dlygate4sd3_1
X_19939_ net3284 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
Xhold2926 _08378_ vssd1 vssd1 vccd1 vccd1 net3453 sky130_fd_sc_hd__buf_2
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2937 net5776 vssd1 vssd1 vccd1 vccd1 net3464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2948 net7916 vssd1 vssd1 vccd1 vccd1 net3475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2959 _02967_ vssd1 vssd1 vccd1 vccd1 net3486 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_103_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21901_ net343 net3204 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21832_ net274 net2556 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21763_ clknet_leaf_83_i_clk net4072 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20714_ net960 net5380 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nor2_1
X_21694_ clknet_leaf_24_i_clk net4022 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6220 _04395_ vssd1 vssd1 vccd1 vccd1 net6747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6231 net2131 vssd1 vssd1 vccd1 vccd1 net6758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6242 _04440_ vssd1 vssd1 vccd1 vccd1 net6769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6253 net1721 vssd1 vssd1 vccd1 vccd1 net6780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6264 rbzero.spi_registers.sclk_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6275 net1824 vssd1 vssd1 vccd1 vccd1 net6802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5530 gpout5.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6286 _04202_ vssd1 vssd1 vccd1 vccd1 net6813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5541 net2075 vssd1 vssd1 vccd1 vccd1 net6068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5552 rbzero.spi_registers.new_texadd\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net6079
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6297 net2102 vssd1 vssd1 vccd1 vccd1 net6824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5563 net934 vssd1 vssd1 vccd1 vccd1 net6090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5574 _04016_ vssd1 vssd1 vccd1 vccd1 net6101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4840 rbzero.spi_registers.texadd1\[22\] vssd1 vssd1 vccd1 vccd1 net5367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5585 _04019_ vssd1 vssd1 vccd1 vccd1 net6112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4851 net885 vssd1 vssd1 vccd1 vccd1 net5378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5596 _04003_ vssd1 vssd1 vccd1 vccd1 net6123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4862 _00817_ vssd1 vssd1 vccd1 vccd1 net5389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4873 net872 vssd1 vssd1 vccd1 vccd1 net5400 sky130_fd_sc_hd__buf_1
XFILLER_0_79_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4884 rbzero.spi_registers.texadd1\[19\] vssd1 vssd1 vccd1 vccd1 net5411 sky130_fd_sc_hd__dlygate4sd3_1
X_21128_ clknet_leaf_33_i_clk net4046 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_1
Xhold4895 net1014 vssd1 vssd1 vccd1 vccd1 net5422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21059_ clknet_leaf_68_i_clk _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13950_ _06813_ _06695_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__or2_1
X_12901_ net3431 net3998 vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ _07042_ _07048_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _08682_ _08713_ _08714_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__nand3_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12832_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _08627_ _08645_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__xor2_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12763_ net51 _05902_ _05915_ net40 vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a22o_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _07638_ _07636_ _07637_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__nand3_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18270_ net6476 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__buf_1
X_11714_ _04885_ _04903_ net654 net3388 _04861_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a2111o_2
X_15482_ _08571_ _08576_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__nand2_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _04648_ _04461_ _04468_ _04023_ _05851_ _05850_ vssd1 vssd1 vccd1 vccd1 _05872_
+ sky130_fd_sc_hd__mux4_1
X_17221_ _10182_ _10240_ vssd1 vssd1 vccd1 vccd1 _10241_ sky130_fd_sc_hd__xnor2_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _07581_ _07602_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__nor2_1
X_11645_ net4450 _04813_ _04834_ _04794_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_86_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17152_ _10170_ _10171_ vssd1 vssd1 vccd1 vccd1 _10172_ sky130_fd_sc_hd__nor2_1
Xinput15 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_2
X_14364_ _07485_ _07496_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11576_ net1101 net4230 vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__nand2_1
Xinput26 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
Xinput37 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16103_ _09015_ _09050_ _09196_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
XFILLER_0_107_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13315_ _06430_ _06432_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__nand2_1
X_10527_ net5549 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__clkbuf_1
X_17083_ _08573_ _09673_ vssd1 vssd1 vccd1 vccd1 _10104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ _06832_ _07233_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ _09126_ _09127_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__nor2_1
X_10458_ net2027 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__clkbuf_1
X_13246_ net8217 _06416_ _06415_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13177_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
X_12128_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _04950_ vssd1 vssd1 vccd1 vccd1 _05316_
+ sky130_fd_sc_hd__mux2_1
X_17985_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__xor2_1
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16936_ _08880_ _09292_ _08246_ _09288_ vssd1 vssd1 vccd1 vccd1 _09958_ sky130_fd_sc_hd__a2bb2o_1
X_12059_ _04949_ _05245_ _05247_ _05233_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__o211a_1
X_19724_ net7273 _03492_ net2310 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a21boi_2
X_16867_ _09632_ _09597_ vssd1 vssd1 vccd1 vccd1 _09889_ sky130_fd_sc_hd__or2b_1
X_19655_ net6619 net3481 _03429_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__mux2_1
X_15818_ _08902_ _08911_ _08912_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__a21oi_1
X_18606_ net4423 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__inv_2
X_19586_ net6464 net3745 net1779 vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__mux2_1
X_20404__156 clknet_1_0__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__inv_2
X_16798_ _09824_ net4631 _09826_ vssd1 vssd1 vccd1 vccd1 _09827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18537_ _02709_ net5974 _06242_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
X_15749_ _08833_ _08842_ _08843_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ _02614_ _02632_ _02607_ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17419_ _10435_ _10436_ vssd1 vssd1 vccd1 vccd1 _10437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18399_ net4724 rbzero.wall_tracer.rayAddendX\[1\] vssd1 vssd1 vccd1 vccd1 _02582_
+ sky130_fd_sc_hd__or2_1
X_20361_ clknet_1_1__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__buf_1
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22100_ net162 net2133 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4103 net3889 vssd1 vssd1 vccd1 vccd1 net4630 sky130_fd_sc_hd__clkbuf_2
X_20292_ net6510 net4038 _03814_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4114 net5936 vssd1 vssd1 vccd1 vccd1 net4641 sky130_fd_sc_hd__buf_1
Xhold4125 net8404 vssd1 vssd1 vccd1 vccd1 net4652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22031_ net473 net1440 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4136 net3477 vssd1 vssd1 vccd1 vccd1 net4663 sky130_fd_sc_hd__dlygate4sd3_1
X_20485__228 clknet_1_1__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__inv_2
XFILLER_0_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4147 net4290 vssd1 vssd1 vccd1 vccd1 net4674 sky130_fd_sc_hd__buf_4
Xhold3402 _03747_ vssd1 vssd1 vccd1 vccd1 net3929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3413 net3851 vssd1 vssd1 vccd1 vccd1 net3940 sky130_fd_sc_hd__clkbuf_2
Xhold4158 net3013 vssd1 vssd1 vccd1 vccd1 net4685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3424 _03781_ vssd1 vssd1 vccd1 vccd1 net3951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4169 _00425_ vssd1 vssd1 vccd1 vccd1 net4696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3435 net7688 vssd1 vssd1 vccd1 vccd1 net3962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2701 _03573_ vssd1 vssd1 vccd1 vccd1 net3228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3446 net8053 vssd1 vssd1 vccd1 vccd1 net3973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 _01156_ vssd1 vssd1 vccd1 vccd1 net3239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3457 _06103_ vssd1 vssd1 vccd1 vccd1 net3984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2723 _04233_ vssd1 vssd1 vccd1 vccd1 net3250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3468 net6043 vssd1 vssd1 vccd1 vccd1 net3995 sky130_fd_sc_hd__buf_1
Xhold2734 _03565_ vssd1 vssd1 vccd1 vccd1 net3261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3479 net4047 vssd1 vssd1 vccd1 vccd1 net4006 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2745 rbzero.pov.spi_buffer\[34\] vssd1 vssd1 vccd1 vccd1 net3272 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2756 net2860 vssd1 vssd1 vccd1 vccd1 net3283 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2767 _00676_ vssd1 vssd1 vccd1 vccd1 net3294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2778 net7271 vssd1 vssd1 vccd1 vccd1 net3305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2789 net5860 vssd1 vssd1 vccd1 vccd1 net3316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21815_ net257 net1799 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
X_20379__133 clknet_1_1__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__inv_2
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire83 net1608 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21746_ clknet_leaf_134_i_clk net3541 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21677_ clknet_leaf_124_i_clk net2891 vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _04496_ _04617_ _04619_ _04621_ _04494_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ rbzero.spi_registers.texadd2\[14\] _04506_ _04507_ _04552_ vssd1 vssd1 vccd1
+ vccd1 _04553_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6050 rbzero.spi_registers.new_leak\[4\] vssd1 vssd1 vccd1 vccd1 net6577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6061 _04249_ vssd1 vssd1 vccd1 vccd1 net6588 sky130_fd_sc_hd__dlygate4sd3_1
X_13100_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xor2_2
XFILLER_0_81_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6072 net1691 vssd1 vssd1 vccd1 vccd1 net6599 sky130_fd_sc_hd__dlygate4sd3_1
X_14080_ _06914_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__inv_2
X_11292_ net3976 net4083 _04485_ net3871 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6083 rbzero.spi_registers.mosi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6094 net1650 vssd1 vssd1 vccd1 vccd1 net6621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5360 net3370 vssd1 vssd1 vccd1 vccd1 net5887 sky130_fd_sc_hd__buf_2
Xhold5371 net3015 vssd1 vssd1 vccd1 vccd1 net5898 sky130_fd_sc_hd__buf_1
X_13031_ net4669 vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__inv_2
Xhold5382 _03641_ vssd1 vssd1 vccd1 vccd1 net5909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5393 net3966 vssd1 vssd1 vccd1 vccd1 net5920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4670 net880 vssd1 vssd1 vccd1 vccd1 net5197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4681 _03791_ vssd1 vssd1 vccd1 vccd1 net5208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4692 rbzero.spi_registers.texadd0\[19\] vssd1 vssd1 vccd1 vccd1 net5219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17770_ _01818_ _01925_ _01815_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a21boi_1
Xclkbuf_4_12__f_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold3980 net7981 vssd1 vssd1 vccd1 vccd1 net4507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3991 net3378 vssd1 vssd1 vccd1 vccd1 net4518 sky130_fd_sc_hd__clkbuf_2
X_14982_ net4756 _08028_ _08079_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16721_ _09757_ _09758_ vssd1 vssd1 vccd1 vccd1 _09759_ sky130_fd_sc_hd__nor2_1
X_13933_ net83 vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_199_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19440_ net2232 net3644 _03323_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ net4089 net5949 _09720_ vssd1 vssd1 vccd1 vccd1 _09732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13864_ net80 _06708_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15603_ _08349_ _08348_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__and2b_1
X_12815_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__inv_2
X_19371_ net5025 _03283_ _03287_ _03288_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16583_ net3507 _09413_ _08441_ _09672_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__a22o_2
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13795_ _06768_ _06931_ _06727_ _06758_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__and4_1
X_18322_ _05155_ net693 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nand2_1
X_15534_ _08571_ _08574_ _08575_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__a21o_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ net4103 net4024 net34 vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20590__323 clknet_1_1__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__inv_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18253_ net4413 net3590 _06057_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a21o_1
X_15465_ _08558_ _08559_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12677_ _05849_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17204_ _10221_ _10222_ _10223_ vssd1 vssd1 vccd1 vccd1 _10224_ sky130_fd_sc_hd__nand3_1
X_14416_ _07564_ _07565_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__03842_ clknet_0__03842_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03842_
+ sky130_fd_sc_hd__clkbuf_16
X_11628_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__clkbuf_8
X_18184_ _02406_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15396_ _08133_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__buf_2
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17135_ _10153_ _10154_ vssd1 vssd1 vccd1 vccd1 _10155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _07472_ _07475_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ net3642 vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__inv_2
Xhold607 _03153_ vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 net2800 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17066_ _08391_ _09292_ _09411_ _08880_ vssd1 vssd1 vccd1 vccd1 _10087_ sky130_fd_sc_hd__o22ai_1
Xhold629 net5463 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14278_ _07436_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16017_ _08529_ _08614_ _09063_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13229_ _06310_ _06367_ _06381_ _06385_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a31o_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2008 _01445_ vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 _04330_ vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 net6652 vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1318 net6839 vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
X_17968_ _08612_ _09181_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__nor2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 net3018 vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_19707_ net6078 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
X_16919_ _09641_ _09642_ vssd1 vssd1 vccd1 vccd1 _09941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899_ _02000_ _02039_ _02037_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19638_ net1484 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19569_ net6397 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21600_ clknet_leaf_130_i_clk net3212 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21531_ clknet_leaf_135_i_clk net3710 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21462_ clknet_leaf_18_i_clk net2106 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21393_ clknet_leaf_39_i_clk net5462 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20275_ _03689_ net4099 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3210 rbzero.spi_registers.spi_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net3737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22014_ net456 net2407 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold3221 net7840 vssd1 vssd1 vccd1 vccd1 net3748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3232 _02891_ vssd1 vssd1 vccd1 vccd1 net3759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3243 net1878 vssd1 vssd1 vccd1 vccd1 net3770 sky130_fd_sc_hd__clkbuf_4
Xhold3254 net7664 vssd1 vssd1 vccd1 vccd1 net3781 sky130_fd_sc_hd__buf_2
Xhold2520 _01090_ vssd1 vssd1 vccd1 vccd1 net3047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3265 rbzero.spi_registers.mosi vssd1 vssd1 vccd1 vccd1 net3792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3276 net3359 vssd1 vssd1 vccd1 vccd1 net3803 sky130_fd_sc_hd__clkbuf_2
Xhold2531 _00668_ vssd1 vssd1 vccd1 vccd1 net3058 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2542 _01596_ vssd1 vssd1 vccd1 vccd1 net3069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3287 net5875 vssd1 vssd1 vccd1 vccd1 net3814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3298 net7657 vssd1 vssd1 vccd1 vccd1 net3825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2553 net7612 vssd1 vssd1 vccd1 vccd1 net3080 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 _01370_ vssd1 vssd1 vccd1 vccd1 net3091 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03862_ clknet_0__03862_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03862_
+ sky130_fd_sc_hd__clkbuf_16
Xhold1830 net7098 vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2575 _03530_ vssd1 vssd1 vccd1 vccd1 net3102 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1841 _04370_ vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2586 _00657_ vssd1 vssd1 vccd1 vccd1 net3113 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1852 net5665 vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 rbzero.pov.spi_buffer\[36\] vssd1 vssd1 vccd1 vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1863 net7223 vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1874 _01411_ vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ net7532 net7433 _04276_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1885 _03574_ vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1896 net6913 vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ net2477 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12600_ net19 net18 net20 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a21o_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ _06741_ _06749_ _06718_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__o21a_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10792_ net6993 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _05700_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__inv_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21729_ clknet_leaf_101_i_clk net4419 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15250_ _08343_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__xnor2_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12462_ _05633_ net5 vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__and2b_1
X_14201_ _07333_ _07371_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__nand2_1
X_11413_ _04542_ _04515_ _04540_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_93 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_93/HI o_rgb[0] sky130_fd_sc_hd__conb_1
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ net4539 _08123_ _06118_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04951_ vssd1 vssd1 vccd1 vccd1 _05578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14132_ _07243_ _07279_ _07299_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__a22o_4
X_20433__182 clknet_1_0__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__inv_2
X_11344_ _04517_ _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18940_ net3214 net7334 _03036_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
X_14063_ _06699_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__nor2_1
X_11275_ _04023_ _04470_ net4133 net4089 vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__or4b_1
Xhold5190 rbzero.tex_b1\[49\] vssd1 vssd1 vccd1 vccd1 net5717 sky130_fd_sc_hd__dlygate4sd3_1
X_13014_ _06166_ _06168_ _06171_ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__and4b_1
XFILLER_0_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18871_ net2469 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
X_17822_ _01999_ _01969_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17753_ _01872_ _01881_ _01879_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a21oi_1
X_14965_ _08080_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19802__79 clknet_1_1__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__inv_2
X_16704_ net991 _09745_ _09746_ net8088 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a22o_1
X_13916_ _07040_ _07066_ _07086_ _07079_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__a2bb2o_1
X_17684_ _01807_ _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14896_ rbzero.wall_tracer.visualWallDist\[-8\] _08037_ _08038_ vssd1 vssd1 vccd1
+ vccd1 _08042_ sky130_fd_sc_hd__o21a_1
X_16635_ _09721_ net3858 _09722_ vssd1 vssd1 vccd1 vccd1 _09723_ sky130_fd_sc_hd__and3_1
X_19423_ net2441 net3902 _03141_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13847_ _06974_ _07007_ _07017_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ _09535_ _09538_ _09534_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__a21bo_1
X_19354_ net5360 _03269_ _03278_ _03275_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13778_ net549 _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15517_ net8265 _08119_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__nand2_4
X_18305_ net6603 net3674 _02493_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ net38 net37 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__and2b_1
X_19285_ net1286 _03238_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__or2_1
X_16497_ _09576_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7509 rbzero.wall_tracer.stepDistY\[-6\] vssd1 vssd1 vccd1 vccd1 net8036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18236_ _02450_ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__nand2_1
X_15448_ _08529_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6808 rbzero.tex_g1\[21\] vssd1 vssd1 vccd1 vccd1 net7335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6819 net2706 vssd1 vssd1 vccd1 vccd1 net7346 sky130_fd_sc_hd__dlygate4sd3_1
X_18167_ _09809_ _02390_ _02391_ _09880_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15379_ _08473_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17118_ _10015_ vssd1 vssd1 vccd1 vccd1 _10138_ sky130_fd_sc_hd__inv_2
Xhold404 net5311 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03856_ _03856_ vssd1 vssd1 vccd1 vccd1 clknet_0__03856_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ _02329_ net3730 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__or2b_1
Xhold415 net4878 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold426 net5359 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 net6113 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 net2796 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ _10068_ _10069_ vssd1 vssd1 vccd1 vccd1 _10070_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold459 net6471 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20060_ net5929 _03610_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 net6453 vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _00925_ vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 net6644 vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1137 net4586 vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1148 net8112 vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 net6571 vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20597__329 clknet_1_0__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__inv_2
XFILLER_0_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20962_ clknet_leaf_74_i_clk _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20893_ _03312_ net2614 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21514_ clknet_leaf_8_i_clk net1351 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21445_ clknet_leaf_17_i_clk net3088 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21376_ clknet_leaf_46_i_clk net5107 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20327_ net6080 net3481 _03813_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold960 net6616 vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 _01005_ vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11060_ _04193_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__clkbuf_4
Xhold982 _02491_ vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 net6487 vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_20258_ net3970 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__inv_2
Xhold3040 _03751_ vssd1 vssd1 vccd1 vccd1 net3567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3051 _01235_ vssd1 vssd1 vccd1 vccd1 net3578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3062 _02464_ vssd1 vssd1 vccd1 vccd1 net3589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3073 net8329 vssd1 vssd1 vccd1 vccd1 net3600 sky130_fd_sc_hd__dlygate4sd3_1
X_20189_ net4733 _03744_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or2_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3084 rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 net3611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2350 net7952 vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3095 _01234_ vssd1 vssd1 vccd1 vccd1 net3622 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2361 _01397_ vssd1 vssd1 vccd1 vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2372 net5828 vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2383 net8310 vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03845_ clknet_0__03845_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03845_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 _03542_ vssd1 vssd1 vccd1 vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1660 net7094 vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1671 net5844 vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__buf_1
X_14750_ net4539 _07917_ _07872_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__mux2_1
Xhold1682 net7158 vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ net3660 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__clkbuf_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1693 net6682 vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _06866_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__and2b_1
X_10913_ _04264_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__clkbuf_4
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _07818_ _07849_ _07851_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__o21ba_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ net4107 _05081_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16420_ _09509_ _09510_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__and2_1
X_13632_ _06756_ _06760_ _06766_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__and3_1
X_10844_ net7049 net7111 _04238_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xsplit42 _07304_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
X_16351_ _09440_ _09442_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__nor2_1
X_13563_ _06663_ _06673_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10775_ net2534 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15302_ _08377_ _08388_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19070_ net3941 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__clkbuf_1
X_12514_ _05690_ _05692_ _05693_ _05694_ net14 vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a32o_1
X_16282_ _08996_ _09373_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13494_ _06547_ _06630_ _06543_ _06505_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__o211a_1
X_18021_ _02196_ _02197_ _02198_ _02199_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__o22a_1
X_15233_ net4535 _08162_ _08126_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__o21bai_4
X_12445_ _05629_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ _08258_ net3433 net7776 vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__mux2_1
X_12376_ rbzero.tex_b1\[27\] rbzero.tex_b1\[26\] _04924_ vssd1 vssd1 vccd1 vccd1 _05561_
+ sky130_fd_sc_hd__mux2_1
X_14115_ _07256_ _07264_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11327_ rbzero.texu_hot\[3\] _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19972_ net6667 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ _08188_ _08189_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__and2_1
X_18923_ net3256 net7613 _03025_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
X_14046_ _07211_ _07215_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or2_1
X_11258_ net5628 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_114_i_clk clknet_4_3__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18854_ net2873 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11189_ net2726 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17805_ _01857_ _01938_ _01937_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a21oi_1
X_18785_ net6048 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__clkbuf_1
X_15997_ net8220 net8227 net4182 vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _08071_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
X_17736_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_129_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17667_ _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14879_ net8370 _07988_ _07869_ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19406_ net1671 _03303_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ _09704_ _09706_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17598_ _01737_ _01738_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16549_ _09503_ _09638_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19337_ net1020 _03140_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7306 _06436_ vssd1 vssd1 vccd1 vccd1 net7833 sky130_fd_sc_hd__buf_2
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19268_ net5308 _03216_ _03227_ _03219_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__o211a_1
Xhold7328 net4228 vssd1 vssd1 vccd1 vccd1 net7855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7339 rbzero.wall_tracer.stepDistX\[-5\] vssd1 vssd1 vccd1 vccd1 net7866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6605 _04252_ vssd1 vssd1 vccd1 vccd1 net7132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18219_ _02427_ _02430_ _02428_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__o21a_1
Xhold6616 net1915 vssd1 vssd1 vccd1 vccd1 net7143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19199_ net5372 _03182_ _03187_ _03176_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__o211a_1
Xhold6627 rbzero.pov.ready_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net7154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6638 net2499 vssd1 vssd1 vccd1 vccd1 net7165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21230_ clknet_leaf_126_i_clk net1981 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6649 _03590_ vssd1 vssd1 vccd1 vccd1 net7176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5904 _03454_ vssd1 vssd1 vccd1 vccd1 net6431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5915 net1352 vssd1 vssd1 vccd1 vccd1 net6442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 net5010 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5926 rbzero.spi_registers.new_texadd\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net6453
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5937 net1176 vssd1 vssd1 vccd1 vccd1 net6464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 net5142 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold223 net5192 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5948 rbzero.spi_registers.spi_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net6475 sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ clknet_leaf_130_i_clk net3353 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5959 net1076 vssd1 vssd1 vccd1 vccd1 net6486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 net5118 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 net5146 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold256 net5176 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold267 net5162 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _01393_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
X_20112_ _03699_ _03700_ _03701_ net3553 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 net7333 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
X_21092_ clknet_leaf_47_i_clk net1633 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20043_ net5898 _03631_ _03647_ _03648_ _03607_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__o221a_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ net436 net1928 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ clknet_leaf_69_i_clk net4677 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _09739_ net4424 _04010_ _02508_ net8097 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ net6195 net6922 _04086_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20651__378 clknet_1_0__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__inv_2
XFILLER_0_107_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7840 net3776 vssd1 vssd1 vccd1 vccd1 net8367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7851 _08182_ vssd1 vssd1 vccd1 vccd1 net8378 sky130_fd_sc_hd__dlygate4sd3_1
X_10491_ net6977 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7873 _08432_ vssd1 vssd1 vccd1 vccd1 net8400 sky130_fd_sc_hd__buf_1
XFILLER_0_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _04837_ vssd1 vssd1 vccd1 vccd1 _05417_
+ sky130_fd_sc_hd__mux2_1
Xhold7884 _08153_ vssd1 vssd1 vccd1 vccd1 net8411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21428_ clknet_leaf_36_i_clk net2234 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7895 _08174_ vssd1 vssd1 vccd1 vccd1 net8422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12161_ _05343_ _05345_ _05348_ _04988_ _04824_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_i_clk clknet_4_11__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21359_ clknet_leaf_7_i_clk net5179 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11112_ net6892 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
X_12092_ _05279_ _05280_ _04977_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__mux2_1
Xhold790 net6414 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ net2778 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
X_15920_ _08993_ _09014_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__xnor2_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_0__f_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_46_i_clk clknet_4_8__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _08941_ _08945_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__xor2_1
X_20545__283 clknet_1_0__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__inv_2
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2180 _04347_ vssd1 vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2191 rbzero.tex_r1\[25\] vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
X_14802_ net7813 _07876_ _07879_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__and3_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15782_ _08861_ _08875_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__and2_1
X_18570_ net7714 net4034 net4648 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ net3757 vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__inv_2
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1490 net7227 vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _08472_ _08614_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__or2_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ net7839 _07898_ _07901_ net7833 vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__o211ai_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11945_ _05074_ _05094_ _05133_ net4118 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _09537_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__nor2_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ _06696_ _07360_ _07442_ net8491 vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__o211a_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19792__70 clknet_1_1__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_0_19_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11876_ _04665_ net3918 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__or2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16403_ _09491_ _09492_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ _06730_ _06728_ _06721_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__a21oi_1
X_17383_ _10151_ _10278_ _10281_ vssd1 vssd1 vccd1 vccd1 _10401_ sky130_fd_sc_hd__a21oi_1
X_10827_ net6211 net6750 _04227_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14595_ _07739_ _07748_ _07747_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16334_ _09408_ _09425_ vssd1 vssd1 vccd1 vccd1 _09426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19122_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__clkbuf_4
X_13546_ _06714_ _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10758_ net2288 net6203 _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19053_ net7617 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__clkbuf_1
X_16265_ _09352_ _09353_ _09356_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13477_ _06462_ _06571_ _06578_ _06551_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__a211o_1
XFILLER_0_168_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10689_ net7348 net7095 _04149_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15216_ _08307_ _08310_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__nand2_2
XFILLER_0_164_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18004_ net4762 net4388 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__or2_1
X_12428_ _05611_ _05612_ _04984_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ _08402_ _09165_ _09288_ net7836 vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _08206_ _08221_ _08229_ _08241_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12359_ _04656_ net4067 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__nor2_1
Xhold3809 net8154 vssd1 vssd1 vccd1 vccd1 net4336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19955_ net2927 net7175 _03583_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__mux2_1
X_15078_ net7765 net8413 vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__nand2_1
X_14029_ _07138_ _07137_ _07186_ _07188_ _07189_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__a32o_2
X_18906_ net3173 net7548 _03014_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
X_19886_ net7516 net3256 _03550_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__mux2_1
X_18837_ net3935 net1547 net3909 net5845 vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__and4_1
XFILLER_0_175_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ _02915_ _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__xnor2_1
X_17719_ _01956_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18699_ _02832_ _02838_ _02826_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20730_ net5252 _03877_ _03874_ _03908_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7103 rbzero.wall_tracer.mapX\[5\] vssd1 vssd1 vccd1 vccd1 net7630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7125 _03720_ vssd1 vssd1 vccd1 vccd1 net7652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7136 net3691 vssd1 vssd1 vccd1 vccd1 net7663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6402 _04099_ vssd1 vssd1 vccd1 vccd1 net6929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7147 _03496_ vssd1 vssd1 vccd1 vccd1 net7674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6413 net2026 vssd1 vssd1 vccd1 vccd1 net6940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7158 net3703 vssd1 vssd1 vccd1 vccd1 net7685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6424 rbzero.tex_r1\[51\] vssd1 vssd1 vccd1 vccd1 net6951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7169 rbzero.spi_registers.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 net7696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6435 rbzero.tex_r0\[9\] vssd1 vssd1 vccd1 vccd1 net6962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5701 _04183_ vssd1 vssd1 vccd1 vccd1 net6228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6446 net2279 vssd1 vssd1 vccd1 vccd1 net6973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6457 rbzero.tex_r1\[23\] vssd1 vssd1 vccd1 vccd1 net6984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5712 net1165 vssd1 vssd1 vccd1 vccd1 net6239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6468 net2167 vssd1 vssd1 vccd1 vccd1 net6995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5723 _04332_ vssd1 vssd1 vccd1 vccd1 net6250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6479 _04235_ vssd1 vssd1 vccd1 vccd1 net7006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5734 net1236 vssd1 vssd1 vccd1 vccd1 net6261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5745 _04376_ vssd1 vssd1 vccd1 vccd1 net6272 sky130_fd_sc_hd__dlygate4sd3_1
X_21213_ clknet_leaf_118_i_clk net2428 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5756 net1263 vssd1 vssd1 vccd1 vccd1 net6283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5767 _04246_ vssd1 vssd1 vccd1 vccd1 net6294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5778 net1301 vssd1 vssd1 vccd1 vccd1 net6305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5789 rbzero.spi_registers.new_texadd\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net6316
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21144_ clknet_leaf_102_i_clk net3754 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_21075_ clknet_leaf_76_i_clk _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20026_ _03615_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21977_ net419 net1996 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer60 _06734_ vssd1 vssd1 vccd1 vccd1 net3607 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _04911_ _04914_ _04918_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__o211a_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ clknet_leaf_60_i_clk net4673 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _04802_ _04814_ _04822_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nor3_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20859_ net4229 _04001_ _04002_ _10009_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a22o_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13400_ _06528_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__buf_2
XFILLER_0_193_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10612_ net7009 net2959 _04116_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14380_ _07535_ _07549_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__nor2_1
X_11592_ _04777_ _04778_ net1616 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13331_ _06434_ _06442_ _06454_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__or4_4
X_10543_ net1839 net6088 _04075_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16050_ _09142_ _09143_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7670 _03929_ vssd1 vssd1 vccd1 vccd1 net8197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ _06424_ _06426_ _06430_ _06432_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__and4b_1
X_10474_ net7123 net7365 _04042_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__mux2_1
Xhold7681 rbzero.traced_texa\[4\] vssd1 vssd1 vccd1 vccd1 net8208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7692 net8541 vssd1 vssd1 vccd1 vccd1 net8219 sky130_fd_sc_hd__dlygate4sd3_1
X_15001_ _06102_ _06158_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__or2_1
X_12213_ rbzero.tex_g1\[23\] rbzero.tex_g1\[22\] _04923_ vssd1 vssd1 vccd1 vccd1 _05400_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6980 rbzero.pov.ready_buffer\[9\] vssd1 vssd1 vccd1 vccd1 net7507 sky130_fd_sc_hd__dlygate4sd3_1
X_13193_ _06296_ _06299_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__xor2_2
Xhold6991 net3356 vssd1 vssd1 vccd1 vccd1 net7518 sky130_fd_sc_hd__dlygate4sd3_1
X_12144_ _04991_ _05323_ _05331_ _04849_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a31o_1
XFILLER_0_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19740_ net3825 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__clkbuf_1
X_12075_ _05233_ _05257_ _05262_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a211o_1
X_16952_ _09676_ _09546_ _06124_ vssd1 vssd1 vccd1 vccd1 _09974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11026_ net5720 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
X_15903_ _08995_ _08997_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19671_ net6440 net4038 _03457_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
X_16883_ _09903_ _09904_ vssd1 vssd1 vccd1 vccd1 _09905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18622_ _02771_ _02772_ _02773_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__o21a_1
X_15834_ _08889_ _08885_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__nand2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ net4045 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__clkbuf_1
X_15765_ _08831_ _08845_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__xnor2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ net1817 _06061_ _06043_ net4324 vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__o22a_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _01679_ _10429_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__or2b_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ net4019 _05115_ _05116_ net3682 _04659_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a221o_1
X_14716_ net8444 _07849_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__nor2_1
X_15696_ _08719_ _08789_ _08788_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__a21o_1
X_18484_ _02660_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__xnor2_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17435_ _10430_ _10431_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14647_ net7807 vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__buf_2
X_11859_ net4115 net4132 net4145 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _10009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ net4651 net4522 vssd1 vssd1 vccd1 vccd1 _10384_ sky130_fd_sc_hd__or2_1
X_14578_ _07747_ _07748_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19105_ net889 _03126_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__or2_1
X_16317_ net3542 _08491_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__nand2_1
X_13529_ _06607_ _06617_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17297_ _08421_ _08424_ _08426_ vssd1 vssd1 vccd1 vccd1 _10316_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ _09239_ _09240_ _09339_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19036_ net7698 net3838 net3398 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5008 net1700 vssd1 vssd1 vccd1 vccd1 net5535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5019 net2123 vssd1 vssd1 vccd1 vccd1 net5546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16179_ _08509_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__clkbuf_4
Xhold4307 _03386_ vssd1 vssd1 vccd1 vccd1 net4834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4318 _00964_ vssd1 vssd1 vccd1 vccd1 net4845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4329 _02907_ vssd1 vssd1 vccd1 vccd1 net4856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3606 _04024_ vssd1 vssd1 vccd1 vccd1 net4133 sky130_fd_sc_hd__clkbuf_4
Xhold3617 gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 net4144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3628 _04752_ vssd1 vssd1 vccd1 vccd1 net4155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3639 _00461_ vssd1 vssd1 vccd1 vccd1 net4166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2905 net5900 vssd1 vssd1 vccd1 vccd1 net3432 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03507_ clknet_0__03507_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03507_
+ sky130_fd_sc_hd__clkbuf_16
X_19938_ net3312 net3283 _03572_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__mux2_1
Xhold2916 net8236 vssd1 vssd1 vccd1 vccd1 net3443 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2927 _08421_ vssd1 vssd1 vccd1 vccd1 net3454 sky130_fd_sc_hd__clkbuf_2
Xhold2938 net5778 vssd1 vssd1 vccd1 vccd1 net3465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2949 net7998 vssd1 vssd1 vccd1 vccd1 net3476 sky130_fd_sc_hd__dlygate4sd3_1
X_19869_ net6512 net3173 _03539_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21900_ net342 net2037 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21831_ net273 net2779 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21762_ clknet_leaf_112_i_clk _01249_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20713_ _03889_ _03890_ _03891_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21693_ clknet_leaf_24_i_clk net3685 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19771__51 clknet_1_0__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_0_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6210 net1854 vssd1 vssd1 vccd1 vccd1 net6737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6221 net1762 vssd1 vssd1 vccd1 vccd1 net6748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6232 _04043_ vssd1 vssd1 vccd1 vccd1 net6759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6243 net1953 vssd1 vssd1 vccd1 vccd1 net6770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6254 _04442_ vssd1 vssd1 vccd1 vccd1 net6781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5520 _02932_ vssd1 vssd1 vccd1 vccd1 net6047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6265 net2055 vssd1 vssd1 vccd1 vccd1 net6792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6276 rbzero.tex_b0\[57\] vssd1 vssd1 vccd1 vccd1 net6803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5531 net919 vssd1 vssd1 vccd1 vccd1 net6058 sky130_fd_sc_hd__clkbuf_2
Xhold6287 net1936 vssd1 vssd1 vccd1 vccd1 net6814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5542 _03479_ vssd1 vssd1 vccd1 vccd1 net6069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6298 rbzero.tex_r0\[38\] vssd1 vssd1 vccd1 vccd1 net6825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5553 net1590 vssd1 vssd1 vccd1 vccd1 net6080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5564 rbzero.tex_g0\[52\] vssd1 vssd1 vccd1 vccd1 net6091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5575 rbzero.tex_b0\[50\] vssd1 vssd1 vccd1 vccd1 net6102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4830 _00885_ vssd1 vssd1 vccd1 vccd1 net5357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4841 net946 vssd1 vssd1 vccd1 vccd1 net5368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5586 rbzero.tex_g1\[38\] vssd1 vssd1 vccd1 vccd1 net6113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4852 rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 net5379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5597 rbzero.pov.spi_buffer\[19\] vssd1 vssd1 vccd1 vccd1 net6124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4863 net1012 vssd1 vssd1 vccd1 vccd1 net5390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4874 _01603_ vssd1 vssd1 vccd1 vccd1 net5401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4885 net989 vssd1 vssd1 vccd1 vccd1 net5412 sky130_fd_sc_hd__dlygate4sd3_1
X_21127_ clknet_leaf_33_i_clk net3850 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_1
Xhold4896 rbzero.spi_registers.texadd1\[11\] vssd1 vssd1 vccd1 vccd1 net5423 sky130_fd_sc_hd__dlygate4sd3_1
X_20462__207 clknet_1_0__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__inv_2
X_21058_ clknet_4_13__leaf_i_clk _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12900_ net3431 net3998 vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nand2_1
X_20009_ _03609_ net3544 vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or2_1
X_13880_ _07038_ _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12831_ _05952_ _05955_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__xor2_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _08642_ _08643_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__a21oi_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ net4066 _05902_ _05915_ net71 _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a221o_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _07662_ _07671_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__and2_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ net3388 _04886_ _04901_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a211o_1
X_20657__384 clknet_1_1__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__inv_2
X_15481_ _08571_ _08574_ _08575_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__nand3_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _05863_ _05867_ _05868_ _05853_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a221o_2
XFILLER_0_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17220_ _10237_ _10239_ vssd1 vssd1 vccd1 vccd1 _10240_ sky130_fd_sc_hd__xor2_2
XFILLER_0_182_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20356__112 clknet_1_1__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__inv_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _07581_ _07602_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__xor2_2
X_11644_ _04792_ _04793_ _04789_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ _10164_ _10065_ _10169_ vssd1 vssd1 vccd1 vccd1 _10171_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14363_ _07531_ _07533_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor2_2
X_11575_ _04763_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__nand2_1
Xinput16 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
Xinput27 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dlymetal6s2s_1
X_16102_ _09047_ _09049_ vssd1 vssd1 vccd1 vccd1 _09196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput38 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
XFILLER_0_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13314_ _06467_ _06433_ _06403_ _06468_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__and4_1
Xinput49 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_8
X_10526_ net2152 net5547 _04064_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_1
X_17082_ _08905_ _09970_ vssd1 vssd1 vccd1 vccd1 _10103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20675__20 clknet_1_1__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
X_14294_ _07306_ _07304_ _07280_ _07308_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16033_ _09012_ _09110_ _09125_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ _06303_ _06304_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__and2_1
X_10457_ net6581 net6940 _04031_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ rbzero.wall_tracer.visualWallDist\[-9\] _06010_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _05306_ _05310_ _05314_ _04967_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a211o_1
XFILLER_0_209_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17984_ _02094_ _02095_ _02134_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__o21a_1
X_19723_ net5496 net7685 net5280 _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__and4bb_1
X_16935_ _08880_ _08391_ _09170_ _09292_ vssd1 vssd1 vccd1 vccd1 _09957_ sky130_fd_sc_hd__or4_1
X_12058_ _04977_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__or2_1
X_11009_ net2114 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
X_19654_ net6403 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__clkbuf_1
X_16866_ _08611_ _09593_ net7818 _09887_ vssd1 vssd1 vccd1 vccd1 _09888_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18605_ net4530 _02765_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__xor2_1
X_15817_ _08904_ _08910_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__and2_1
X_19585_ net1478 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
X_16797_ _09813_ _09814_ _09815_ vssd1 vssd1 vccd1 vccd1 _09826_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18536_ net7690 _06061_ _02245_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
X_15748_ _08836_ _08841_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__or2b_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18467_ _02643_ net4820 net8085 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__o21ai_2
X_15679_ _08160_ _08225_ _08227_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17418_ _08472_ _08616_ vssd1 vssd1 vccd1 vccd1 _10436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18398_ net4724 rbzero.wall_tracer.rayAddendX\[1\] vssd1 vssd1 vccd1 vccd1 _02581_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17349_ _10237_ _10239_ vssd1 vssd1 vccd1 vccd1 _10368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19019_ net4030 net1493 _03078_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
X_20291_ net1305 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
Xhold4104 _09825_ vssd1 vssd1 vccd1 vccd1 net4631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4115 _06037_ vssd1 vssd1 vccd1 vccd1 net4642 sky130_fd_sc_hd__clkbuf_2
X_22030_ net472 net2583 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
Xhold4126 net3841 vssd1 vssd1 vccd1 vccd1 net4653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4137 net7985 vssd1 vssd1 vccd1 vccd1 net4664 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__05688_ _05688_ vssd1 vssd1 vccd1 vccd1 clknet_0__05688_ sky130_fd_sc_hd__clkbuf_16
Xhold3403 _01217_ vssd1 vssd1 vccd1 vccd1 net3930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4148 _08062_ vssd1 vssd1 vccd1 vccd1 net4675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4159 rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 net4686 sky130_fd_sc_hd__clkbuf_4
Xhold3414 _03107_ vssd1 vssd1 vccd1 vccd1 net3941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3425 _03782_ vssd1 vssd1 vccd1 vccd1 net3952 sky130_fd_sc_hd__dlygate4sd3_1
X_19808__85 clknet_1_0__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__inv_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3436 _00618_ vssd1 vssd1 vccd1 vccd1 net3963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2702 _01136_ vssd1 vssd1 vccd1 vccd1 net3229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3447 rbzero.trace_state\[2\] vssd1 vssd1 vccd1 vccd1 net3974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2713 rbzero.tex_r1\[39\] vssd1 vssd1 vccd1 vccd1 net3240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3458 _06114_ vssd1 vssd1 vccd1 vccd1 net3985 sky130_fd_sc_hd__buf_1
Xhold2724 _01418_ vssd1 vssd1 vccd1 vccd1 net3251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3469 _05731_ vssd1 vssd1 vccd1 vccd1 net3996 sky130_fd_sc_hd__clkbuf_4
Xhold2735 _01129_ vssd1 vssd1 vccd1 vccd1 net3262 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2746 net1358 vssd1 vssd1 vccd1 vccd1 net3273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2757 _03580_ vssd1 vssd1 vccd1 vccd1 net3284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2768 net7990 vssd1 vssd1 vccd1 vccd1 net3295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2779 _03604_ vssd1 vssd1 vccd1 vccd1 net3306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21814_ net256 net1662 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire84 _04851_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21745_ clknet_leaf_131_i_clk net4638 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21676_ clknet_leaf_124_i_clk net3050 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20627_ clknet_1_0__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__buf_1
XFILLER_0_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _04509_ _04547_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6040 _03440_ vssd1 vssd1 vccd1 vccd1 net6567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6051 net1671 vssd1 vssd1 vccd1 vccd1 net6578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6062 net1588 vssd1 vssd1 vccd1 vccd1 net6589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6073 rbzero.spi_registers.new_texadd\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net6600
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11291_ net3871 net3976 net3774 _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__or4b_2
Xhold6084 net1727 vssd1 vssd1 vccd1 vccd1 net6611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6095 rbzero.spi_registers.new_texadd\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net6622
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5350 net3909 vssd1 vssd1 vccd1 vccd1 net5877 sky130_fd_sc_hd__dlygate4sd3_1
X_13030_ _06205_ net3888 _06202_ net4567 vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__a2bb2o_1
Xhold5361 _01170_ vssd1 vssd1 vccd1 vccd1 net5888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5372 _03649_ vssd1 vssd1 vccd1 vccd1 net5899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5383 gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 net5910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5394 rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 net5921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4660 net863 vssd1 vssd1 vccd1 vccd1 net5187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4671 _00874_ vssd1 vssd1 vccd1 vccd1 net5198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22159_ clknet_leaf_88_i_clk net1094 vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4682 _01243_ vssd1 vssd1 vccd1 vccd1 net5209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4693 net927 vssd1 vssd1 vccd1 vccd1 net5220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3970 net8330 vssd1 vssd1 vccd1 vccd1 net4497 sky130_fd_sc_hd__dlygate4sd3_1
X_14981_ _08088_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
Xhold3981 net3833 vssd1 vssd1 vccd1 vccd1 net4508 sky130_fd_sc_hd__clkbuf_2
Xhold3992 net7808 vssd1 vssd1 vccd1 vccd1 net4519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16720_ net3965 _08194_ vssd1 vssd1 vccd1 vccd1 _09758_ sky130_fd_sc_hd__nor2_1
X_13932_ _06838_ _06849_ _06836_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13863_ _06703_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__nor2_1
X_16651_ net4135 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15602_ _08695_ _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__nand2_2
X_12814_ _05979_ _05982_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__and2b_1
XFILLER_0_202_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19370_ _03205_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__clkbuf_4
X_13794_ _06931_ _06727_ _06758_ _06768_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__a22o_1
X_16582_ _08032_ _09545_ _08421_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18321_ net4733 net4887 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__nor2_1
X_15533_ _08578_ _08583_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__xnor2_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _04468_ _04023_ _05901_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__mux2_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _08555_ _08557_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__and2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ net4413 net3590 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12676_ _05852_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19750__32 clknet_1_0__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17203_ _08948_ _08916_ _09970_ _09976_ vssd1 vssd1 vccd1 vccd1 _10223_ sky130_fd_sc_hd__or4_1
XFILLER_0_53_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14415_ _07543_ _07545_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_182_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11627_ _04814_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or2_4
Xclkbuf_1_1__f__03841_ clknet_0__03841_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03841_
+ sky130_fd_sc_hd__clkbuf_16
X_15395_ _08414_ _08433_ _08489_ _08476_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__a22o_1
X_18183_ _02405_ net3751 _02393_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17134_ _09472_ _09133_ vssd1 vssd1 vccd1 vccd1 _10154_ sky130_fd_sc_hd__and2b_1
Xclkbuf_0__03872_ _03872_ vssd1 vssd1 vccd1 vccd1 clknet_0__03872_ sky130_fd_sc_hd__clkbuf_16
X_14346_ _07514_ _07515_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11558_ _04736_ _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold608 net5506 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ _08880_ _08391_ _09292_ _09411_ vssd1 vssd1 vccd1 vccd1 _10086_ sky130_fd_sc_hd__or4_1
X_10509_ net6259 net6999 _04053_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold619 _03046_ vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ _07446_ _07447_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11489_ net4091 vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__inv_2
X_16016_ _09014_ _08993_ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__or2b_1
X_13228_ _06395_ _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__or2_4
XFILLER_0_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20410__161 clknet_1_1__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__inv_2
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _06270_ _06277_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__and2b_1
Xhold2009 net6889 vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _01502_ vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_17967_ _09040_ _09060_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nor2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1319 net6841 vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
X_19706_ net6076 net3481 _03456_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
X_16918_ _09938_ _09939_ vssd1 vssd1 vccd1 vccd1 _09940_ sky130_fd_sc_hd__and2_1
X_17898_ _02134_ _02135_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__nand2_1
X_19637_ net6434 net3596 _03441_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
X_16849_ net3800 _09871_ _09872_ vssd1 vssd1 vccd1 vccd1 _09873_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_178_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19568_ net6395 net1493 _03403_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18519_ net6017 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19499_ net1622 net6938 _03365_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21530_ clknet_leaf_135_i_clk net5498 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21461_ clknet_leaf_42_i_clk net3004 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21392_ clknet_leaf_39_i_clk net5442 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20274_ net4092 net4071 net4098 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__and3_1
Xhold3200 net7809 vssd1 vssd1 vccd1 vccd1 net3727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22013_ net455 net2157 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold3211 net1334 vssd1 vssd1 vccd1 vccd1 net3738 sky130_fd_sc_hd__buf_2
Xhold3222 net3699 vssd1 vssd1 vccd1 vccd1 net3749 sky130_fd_sc_hd__clkbuf_2
Xhold3233 net4809 vssd1 vssd1 vccd1 vccd1 net3760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3244 _03106_ vssd1 vssd1 vccd1 vccd1 net3771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2510 net4310 vssd1 vssd1 vccd1 vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3255 net7666 vssd1 vssd1 vccd1 vccd1 net3782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2521 net3198 vssd1 vssd1 vccd1 vccd1 net3048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3266 net2046 vssd1 vssd1 vccd1 vccd1 net3793 sky130_fd_sc_hd__clkbuf_2
Xhold3277 net7873 vssd1 vssd1 vccd1 vccd1 net3804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2532 rbzero.pov.spi_buffer\[58\] vssd1 vssd1 vccd1 vccd1 net3059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2543 net7396 vssd1 vssd1 vccd1 vccd1 net3070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3288 rbzero.spi_registers.spi_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net3815 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03861_ clknet_0__03861_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03861_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3299 _01020_ vssd1 vssd1 vccd1 vccd1 net3826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2554 _03029_ vssd1 vssd1 vccd1 vccd1 net3081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1820 _01037_ vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2565 net7321 vssd1 vssd1 vccd1 vccd1 net3092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1831 _04348_ vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2576 _01097_ vssd1 vssd1 vccd1 vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1842 _01294_ vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2587 net5695 vssd1 vssd1 vccd1 vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 net5667 vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 net3095 vssd1 vssd1 vccd1 vccd1 net3125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 _04143_ vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1875 net7170 vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1886 _01137_ vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1897 net6915 vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ net2503 net6587 _04171_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20574__308 clknet_1_0__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__inv_2
XFILLER_0_52_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ net6991 net2408 _04205_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__mux2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ net49 vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__inv_2
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21728_ clknet_leaf_103_i_clk net3714 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ net5 net4 vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and2_1
X_21659_ clknet_leaf_120_i_clk net2905 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_14200_ _07331_ _07332_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__or2_1
X_11412_ _04509_ _04547_ _04551_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15180_ _07917_ net8055 _08112_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__mux2_1
X_12392_ rbzero.tex_b1\[11\] rbzero.tex_b1\[10\] _04951_ vssd1 vssd1 vccd1 vccd1 _05577_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_94 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_94/HI o_rgb[1] sky130_fd_sc_hd__conb_1
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20342__99 clknet_1_0__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__inv_2
X_14131_ _07300_ _07278_ _07301_ _07275_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__o211a_1
X_11343_ rbzero.texu_hot\[4\] _04516_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20468__213 clknet_1_1__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__inv_2
X_14062_ _07232_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__buf_4
X_11274_ _04461_ _04466_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5180 _04122_ vssd1 vssd1 vccd1 vccd1 net5707 sky130_fd_sc_hd__dlygate4sd3_1
X_13013_ net3945 _06172_ _06163_ _06173_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__a2111oi_1
Xhold5191 net2990 vssd1 vssd1 vccd1 vccd1 net5718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18870_ net3026 net7538 _02993_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
Xhold4490 net685 vssd1 vssd1 vccd1 vccd1 net5017 sky130_fd_sc_hd__dlygate4sd3_1
X_17821_ _02057_ _02058_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ _01983_ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__xnor2_1
X_14964_ net4397 _07975_ _08079_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__mux2_1
X_16703_ net971 _09745_ _09746_ net8068 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a22o_1
X_13915_ _07000_ _06813_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__nand2_1
X_17683_ _01919_ _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__xor2_1
XFILLER_0_187_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895_ net3945 _08034_ _08036_ net3932 net4671 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__o221a_1
X_19422_ net3672 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__clkbuf_1
X_16634_ _04496_ _04021_ vssd1 vssd1 vccd1 vccd1 _09722_ sky130_fd_sc_hd__or2_1
X_13846_ _07009_ _07013_ _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20440__187 clknet_1_1__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__inv_2
XFILLER_0_175_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19353_ net6450 _03271_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__or2_1
X_16565_ _08246_ _08430_ _09526_ _09654_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13777_ _06943_ net538 vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ net655 net5640 _04309_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18304_ net6386 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ _08139_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19284_ _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__buf_2
X_12728_ net36 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__inv_2
XFILLER_0_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ _09579_ _09582_ _09580_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235_ net3835 net4524 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nand2_1
X_15447_ _08277_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ net52 _05798_ _05817_ net53 vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6809 net2521 vssd1 vssd1 vccd1 vccd1 net7336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18166_ _02389_ net3666 _02387_ _02381_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__o211a_1
X_15378_ _06119_ net4877 vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17117_ net4657 net4401 vssd1 vssd1 vccd1 vccd1 _10137_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__03855_ _03855_ vssd1 vssd1 vccd1 vccd1 clknet_0__03855_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 net5313 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ _07484_ _07498_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__nor2_1
X_18097_ net3932 net4399 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__nand2_1
Xhold416 net4880 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 net5361 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold438 net6115 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ _08308_ _09165_ vssd1 vssd1 vccd1 vccd1 _10069_ sky130_fd_sc_hd__nor2_1
Xhold449 _04069_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ net3280 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1105 _02490_ vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1116 net6545 vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _01430_ vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1138 net6561 vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 net4800 vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
X_20961_ clknet_leaf_74_i_clk _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20892_ net4928 net6627 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21513_ clknet_leaf_8_i_clk net1491 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20417__167 clknet_1_1__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__inv_2
XFILLER_0_17_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21444_ clknet_leaf_18_i_clk net3335 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21375_ clknet_leaf_45_i_clk net5314 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20326_ net6138 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
Xhold950 net3837 vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 _01460_ vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 net6533 vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20257_ net4025 net6001 _03796_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a21oi_1
Xhold983 _00580_ vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 net6489 vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3030 net7590 vssd1 vssd1 vccd1 vccd1 net3557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3041 _01219_ vssd1 vssd1 vccd1 vccd1 net3568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3063 _02465_ vssd1 vssd1 vccd1 vccd1 net3590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20188_ net4803 _03743_ _03752_ _03732_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__o211a_1
Xhold3074 rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 net3601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2340 _04324_ vssd1 vssd1 vccd1 vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3085 net5956 vssd1 vssd1 vccd1 vccd1 net3612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 net4572 vssd1 vssd1 vccd1 vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3096 net5942 vssd1 vssd1 vccd1 vccd1 net3623 sky130_fd_sc_hd__clkbuf_2
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2362 net7424 vssd1 vssd1 vccd1 vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2373 net7476 vssd1 vssd1 vccd1 vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2384 net7280 vssd1 vssd1 vccd1 vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03844_ clknet_0__03844_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03844_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1650 _04204_ vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2395 _01108_ vssd1 vssd1 vccd1 vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1661 _04159_ vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
X_11961_ net4002 _05135_ _05146_ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a211o_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1672 _02970_ vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1683 _01331_ vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 net6684 vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
X_10912_ net1901 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _06867_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__nand2_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ net7795 _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__nor2_1
X_11892_ _04684_ net4058 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__and2_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ _06766_ _06761_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__or2b_1
X_10843_ net6036 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xsplit32 _06435_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16350_ _09245_ _09313_ _09441_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13562_ net80 _06732_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10774_ net7105 net7381 _04194_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
X_15301_ _08394_ _08395_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__xor2_1
X_12513_ net4149 net4141 net4164 net7727 _05691_ net13 vssd1 vssd1 vccd1 vccd1 _05694_
+ sky130_fd_sc_hd__mux4_1
X_16281_ _08185_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _06522_ _06462_ _06548_ _06499_ _06551_ _06571_ vssd1 vssd1 vccd1 vccd1 _06664_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_192_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18020_ _02062_ _02232_ _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a21oi_1
X_15232_ _08305_ _08318_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ reg_rgb\[23\] _05628_ _05054_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15163_ _08256_ _08257_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__and2_1
X_12375_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _05369_ vssd1 vssd1 vccd1 vccd1 _05560_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ _07268_ _07270_ _07266_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ rbzero.spi_registers.texadd3\[9\] rbzero.spi_registers.texadd1\[9\] rbzero.spi_registers.texadd0\[9\]
+ rbzero.spi_registers.texadd2\[9\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux4_2
X_19971_ net1869 net6665 net2312 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__mux2_1
X_15094_ net3372 _08175_ vssd1 vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18922_ net3277 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
X_14045_ _07211_ _07215_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__nand2_1
X_11257_ net5626 net5566 _04104_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18853_ net3950 net92 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nand2_1
X_11188_ net7089 net6538 _04412_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
X_17804_ _01968_ _02042_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__xnor2_1
X_18784_ net6046 _02931_ _02536_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__mux2_1
X_15996_ _08986_ _08988_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__xor2_4
XFILLER_0_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _09915_ _09612_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__nor2_1
X_14947_ net4353 _07903_ _08068_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20522__262 clknet_1_0__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__inv_2
X_17666_ _01794_ _09664_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__or2_1
X_14878_ _08029_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
X_19405_ net1255 _03302_ net5501 _03299_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16617_ _09704_ _09706_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__nor2_1
X_13829_ net567 _06715_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__nor2_1
X_17597_ _10390_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19336_ net5344 _03235_ _03266_ _03259_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__o211a_1
X_16548_ _09636_ _09637_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__xnor2_1
Xhold8008 _09594_ vssd1 vssd1 vccd1 vccd1 net8535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19267_ net6629 _03217_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__or2_1
X_16479_ _09498_ _09569_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__xnor2_4
Xhold7318 net563 vssd1 vssd1 vccd1 vccd1 net7845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7329 net1138 vssd1 vssd1 vccd1 vccd1 net7856 sky130_fd_sc_hd__dlygate4sd3_1
X_18218_ _02434_ _02435_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__or2b_1
Xhold6606 net2421 vssd1 vssd1 vccd1 vccd1 net7133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6617 rbzero.tex_g0\[60\] vssd1 vssd1 vccd1 vccd1 net7144 sky130_fd_sc_hd__dlygate4sd3_1
X_19198_ net6388 _03183_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6628 net762 vssd1 vssd1 vccd1 vccd1 net7155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6639 rbzero.tex_g0\[41\] vssd1 vssd1 vccd1 vccd1 net7166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5905 net1433 vssd1 vssd1 vccd1 vccd1 net6432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18149_ _02372_ _02375_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__nor2_1
Xhold5916 _04340_ vssd1 vssd1 vccd1 vccd1 net6443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 net5000 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5927 net1631 vssd1 vssd1 vccd1 vccd1 net6454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5938 rbzero.tex_g1\[50\] vssd1 vssd1 vccd1 vccd1 net6465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 net5156 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 net5194 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5949 net1492 vssd1 vssd1 vccd1 vccd1 net6476 sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ clknet_leaf_130_i_clk net3331 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold235 net7154 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold246 net5132 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold257 net5178 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20111_ _03483_ _03694_ _03661_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21oi_1
Xhold268 net5104 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold279 net5243 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21091_ clknet_leaf_47_i_clk net1540 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20042_ net3431 _03642_ _03484_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a21o_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19778__57 clknet_1_0__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21993_ net435 net1126 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20944_ clknet_leaf_70_i_clk net4708 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20875_ net4423 net652 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7830 net4741 vssd1 vssd1 vccd1 vccd1 net8357 sky130_fd_sc_hd__dlygate4sd3_1
X_10490_ net2499 net6975 _04042_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux2_1
Xhold7852 rbzero.wall_tracer.stepDistY\[5\] vssd1 vssd1 vccd1 vccd1 net8379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7863 rbzero.wall_tracer.stepDistX\[-2\] vssd1 vssd1 vccd1 vccd1 net8390 sky130_fd_sc_hd__dlygate4sd3_1
X_21427_ clknet_leaf_35_i_clk net1627 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7885 _08154_ vssd1 vssd1 vccd1 vccd1 net8412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7896 _08180_ vssd1 vssd1 vccd1 vccd1 net8423 sky130_fd_sc_hd__dlygate4sd3_1
X_12160_ _05346_ _05347_ _04938_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__mux2_1
X_21358_ clknet_leaf_14_i_clk net5458 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11111_ net6890 net2578 _04375_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__mux2_1
X_20309_ net6257 net3596 _03825_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__mux2_1
X_12091_ rbzero.tex_r1\[59\] rbzero.tex_r1\[58\] _05220_ vssd1 vssd1 vccd1 vccd1 _05280_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold780 net6473 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
X_21289_ clknet_leaf_27_i_clk net4386 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold791 _01091_ vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net7039 net7218 _04342_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__mux2_1
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _08907_ _08942_ _08943_ _08944_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__o2bb2a_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2170 net5713 vssd1 vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2181 _01315_ vssd1 vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _07963_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__clkbuf_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 net1938 vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _08861_ _08875_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ net3768 vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__inv_2
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _10062_ _01760_ _10433_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1480 net5555 vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 net7229 vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ net7813 _07899_ _07900_ net8354 vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__a31o_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11944_ _04501_ _05092_ _05132_ net3517 _05105_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__o221a_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _09970_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _07815_ _07831_ _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__o21a_1
X_11875_ net3917 _04664_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nor2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _09491_ _09492_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__nor2_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ net2086 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
X_13614_ _06779_ _06784_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17382_ _10398_ _10399_ vssd1 vssd1 vccd1 vccd1 _10400_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ _07758_ _07759_ _07761_ _07750_ _07764_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19121_ _03122_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__buf_4
X_16333_ _09422_ _09424_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10757_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13545_ _06715_ _06697_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19052_ net7615 net3866 net3398 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
X_16264_ _09230_ _09355_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _06645_ _06646_ _06551_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10688_ net6981 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20552__288 clknet_1_0__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__inv_2
X_18003_ net4762 net4388 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__nand2_1
X_12427_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _04924_ vssd1 vssd1 vccd1 vccd1 _05612_
+ sky130_fd_sc_hd__mux2_1
X_15215_ _08255_ _08308_ _08309_ _08280_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_180_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16195_ _08181_ _08450_ _09169_ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15146_ _08240_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__buf_2
X_12358_ _05376_ _05543_ net4140 vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ net5205 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__clkinv_4
X_19954_ net3160 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
X_15077_ _08156_ _08171_ _08148_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__o21a_1
XFILLER_0_205_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _05220_ vssd1 vssd1 vccd1 vccd1 _05475_
+ sky130_fd_sc_hd__mux2_1
X_18905_ net6514 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
X_14028_ _06696_ _07195_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__or3_1
X_19885_ net3234 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18836_ net1547 net3909 net2198 net3935 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20446__193 clknet_1_0__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__inv_2
X_18767_ _02897_ _02900_ _02898_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a21bo_1
X_15979_ _08607_ _08623_ _08606_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17718_ net4723 net4520 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18698_ _02849_ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17649_ _01802_ _01859_ _01887_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20660_ clknet_1_0__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__buf_1
XFILLER_0_147_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19319_ net5177 _03250_ _03257_ _03246_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7104 net3884 vssd1 vssd1 vccd1 vccd1 net7631 sky130_fd_sc_hd__buf_1
Xhold7115 _03735_ vssd1 vssd1 vccd1 vccd1 net7642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7126 net3608 vssd1 vssd1 vccd1 vccd1 net7653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7137 rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1 vccd1 net7664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6403 net1959 vssd1 vssd1 vccd1 vccd1 net6930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7148 _03498_ vssd1 vssd1 vccd1 vccd1 net7675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6414 rbzero.tex_b0\[33\] vssd1 vssd1 vccd1 vccd1 net6941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7159 rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 net7686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6425 net2496 vssd1 vssd1 vccd1 vccd1 net6952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6436 net2122 vssd1 vssd1 vccd1 vccd1 net6963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6447 rbzero.tex_r1\[45\] vssd1 vssd1 vccd1 vccd1 net6974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5702 net1189 vssd1 vssd1 vccd1 vccd1 net6229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6458 net2173 vssd1 vssd1 vccd1 vccd1 net6985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5713 _03585_ vssd1 vssd1 vccd1 vccd1 net6240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5724 net1159 vssd1 vssd1 vccd1 vccd1 net6251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6469 _04400_ vssd1 vssd1 vccd1 vccd1 net6996 sky130_fd_sc_hd__dlygate4sd3_1
X_21212_ clknet_leaf_118_i_clk net2876 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5735 rbzero.spi_registers.new_texadd\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 net6262
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5746 net1226 vssd1 vssd1 vccd1 vccd1 net6273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5757 rbzero.spi_registers.new_texadd\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 net6284
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5768 net1597 vssd1 vssd1 vccd1 vccd1 net6295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5779 rbzero.spi_registers.new_texadd\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net6306
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21143_ clknet_leaf_100_i_clk net4767 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20529__268 clknet_1_0__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__inv_2
X_21074_ clknet_leaf_76_i_clk _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20025_ net3443 _08295_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ net418 net1190 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer50 net3523 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer61 net3607 vssd1 vssd1 vccd1 vccd1 net3634 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ clknet_leaf_75_i_clk net4681 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _04800_ _04814_ _04826_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__nor3_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ net4224 _04001_ _04002_ _09711_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a22o_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ net6189 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ _04777_ _04779_ _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20789_ _03878_ _03957_ net8209 _03883_ net5581 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13330_ _06496_ _06498_ _06500_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__or3_1
XFILLER_0_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ net1913 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ _06428_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__xnor2_2
X_10473_ net6760 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__clkbuf_1
Xhold7671 _01610_ vssd1 vssd1 vccd1 vccd1 net8198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7682 _03958_ vssd1 vssd1 vccd1 vccd1 net8209 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_128_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold7693 net3489 vssd1 vssd1 vccd1 vccd1 net8220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12212_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _04924_ vssd1 vssd1 vccd1 vccd1 _05399_
+ sky130_fd_sc_hd__mux2_1
X_15000_ net4174 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6970 rbzero.pov.spi_buffer\[18\] vssd1 vssd1 vccd1 vccd1 net7497 sky130_fd_sc_hd__dlygate4sd3_1
X_13192_ net8021 _06265_ _06306_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__o21a_1
Xhold6981 net676 vssd1 vssd1 vccd1 vccd1 net7508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6992 rbzero.pov.spi_buffer\[61\] vssd1 vssd1 vccd1 vccd1 net7519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _04955_ _05326_ _05330_ _04824_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a211o_1
X_12074_ _04824_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__clkbuf_8
X_16951_ _08905_ _09970_ _09972_ vssd1 vssd1 vccd1 vccd1 _09973_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ net5669 net5718 _04331_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__mux2_1
X_15902_ _08996_ _08253_ _08545_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__a21bo_1
X_19670_ net1695 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
X_16882_ _09901_ _09902_ vssd1 vssd1 vccd1 vccd1 _09904_ sky130_fd_sc_hd__and2_1
X_18621_ net4635 _02770_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15833_ _08920_ _08927_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__and2_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19757__38 clknet_1_0__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ net7636 net4044 _06242_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
X_15764_ _08826_ _08851_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__xor2_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ net2038 _06039_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17503_ _10406_ _10423_ _10421_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14715_ _07860_ _07804_ _07884_ net7843 vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__a211o_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _02630_ _02648_ _02650_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a21o_1
X_11927_ _05079_ net4108 _05091_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__and3b_1
X_15695_ _08719_ _08788_ _08789_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__nand3_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _01674_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nand2_1
X_14646_ _07814_ _07816_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__xnor2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11858_ net4139 _05041_ net4163 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ net2997 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__clkbuf_1
X_17365_ net4651 net4522 vssd1 vssd1 vccd1 vccd1 _10383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 i_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14577_ _07740_ _07746_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20634__363 clknet_1_0__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__inv_2
X_19104_ net4315 _03125_ net2710 _03128_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ _09402_ _09407_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _06698_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__05742_ clknet_0__05742_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05742_
+ sky130_fd_sc_hd__clkbuf_16
X_17296_ _10217_ _10208_ vssd1 vssd1 vccd1 vccd1 _10315_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19035_ net3397 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__buf_1
X_16247_ _09226_ _09241_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__or2b_1
X_13459_ _06492_ _06591_ _06629_ _06529_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5009 _03137_ vssd1 vssd1 vccd1 vccd1 net5536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16178_ _09246_ _09270_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4308 _03424_ vssd1 vssd1 vccd1 vccd1 net4835 sky130_fd_sc_hd__buf_1
Xhold4319 net1045 vssd1 vssd1 vccd1 vccd1 net4846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15129_ net4415 _08123_ _08148_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3607 _09730_ vssd1 vssd1 vccd1 vccd1 net4134 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_92_i_clk clknet_4_5__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold3618 net4088 vssd1 vssd1 vccd1 vccd1 net4145 sky130_fd_sc_hd__clkbuf_4
Xhold3629 _05053_ vssd1 vssd1 vccd1 vccd1 net4156 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__03506_ clknet_0__03506_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03506_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_195_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19937_ net3313 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
Xhold2906 net8206 vssd1 vssd1 vccd1 vccd1 net3433 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2917 net5870 vssd1 vssd1 vccd1 vccd1 net3444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2928 rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 net3455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2939 net8321 vssd1 vssd1 vccd1 vccd1 net3466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19868_ net3023 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18819_ net3770 _02472_ _02948_ _02955_ _02950_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a311o_1
X_19799_ clknet_1_1__leaf__03506_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__buf_1
XFILLER_0_207_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21830_ net272 net2511 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21761_ clknet_leaf_111_i_clk net4130 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20712_ net5400 _03877_ _03874_ net8232 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21692_ clknet_leaf_114_i_clk net5901 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_45_i_clk clknet_4_8__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6200 net1903 vssd1 vssd1 vccd1 vccd1 net6727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6211 rbzero.spi_registers.new_leak\[5\] vssd1 vssd1 vccd1 vccd1 net6738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6222 rbzero.tex_g1\[15\] vssd1 vssd1 vccd1 vccd1 net6749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6233 net2132 vssd1 vssd1 vccd1 vccd1 net6760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6244 rbzero.tex_g1\[49\] vssd1 vssd1 vccd1 vccd1 net6771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6255 net1722 vssd1 vssd1 vccd1 vccd1 net6782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5510 gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 net6037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6266 _03115_ vssd1 vssd1 vccd1 vccd1 net6793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5521 net3602 vssd1 vssd1 vccd1 vccd1 net6048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6277 net1819 vssd1 vssd1 vccd1 vccd1 net6804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5532 _03873_ vssd1 vssd1 vccd1 vccd1 net6059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5543 net2076 vssd1 vssd1 vccd1 vccd1 net6070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6288 rbzero.spi_registers.new_vinf vssd1 vssd1 vccd1 vccd1 net6815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6299 net1517 vssd1 vssd1 vccd1 vccd1 net6826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5554 _03837_ vssd1 vssd1 vccd1 vccd1 net6081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5565 net803 vssd1 vssd1 vccd1 vccd1 net6092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4820 rbzero.spi_registers.texadd0\[21\] vssd1 vssd1 vccd1 vccd1 net5347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5576 net938 vssd1 vssd1 vccd1 vccd1 net6103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4831 net847 vssd1 vssd1 vccd1 vccd1 net5358 sky130_fd_sc_hd__dlygate4sd3_1
X_22175_ clknet_leaf_68_i_clk net1100 vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5587 net964 vssd1 vssd1 vccd1 vccd1 net6114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4842 _00829_ vssd1 vssd1 vccd1 vccd1 net5369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4853 net854 vssd1 vssd1 vccd1 vccd1 net5380 sky130_fd_sc_hd__buf_1
Xhold5598 net735 vssd1 vssd1 vccd1 vccd1 net6125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4864 rbzero.mapdyw\[1\] vssd1 vssd1 vccd1 vccd1 net5391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21126_ clknet_leaf_33_i_clk net4056 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_1
Xhold4875 net873 vssd1 vssd1 vccd1 vccd1 net5402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4886 _00826_ vssd1 vssd1 vccd1 vccd1 net5413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4897 net1036 vssd1 vssd1 vccd1 vccd1 net5424 sky130_fd_sc_hd__dlygate4sd3_1
X_21057_ clknet_leaf_71_i_clk _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20008_ net3543 _08218_ _03614_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _06004_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__xnor2_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ net50 _05912_ _05916_ net49 _05905_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21959_ net401 net1937 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _07660_ _07661_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__or2_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ net4145 _04887_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nor2_1
X_15480_ _08384_ _08458_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__nor2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _05850_ _05851_ _05869_ _05854_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a31o_1
XFILLER_0_194_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11643_ net1136 _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__or2_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14431_ _07583_ _07600_ _07601_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_182_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17150_ _10164_ _10065_ _10169_ vssd1 vssd1 vccd1 vccd1 _10170_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _04761_ _04762_ net2753 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14362_ _07519_ _07528_ _07530_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dlymetal6s2s_1
X_16101_ _09153_ _09194_ vssd1 vssd1 vccd1 vccd1 _09195_ sky130_fd_sc_hd__xnor2_2
Xinput28 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_4
Xinput39 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
X_10525_ net5698 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__clkbuf_1
X_13313_ _06478_ _06467_ net574 _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17081_ _09673_ _09971_ vssd1 vssd1 vccd1 vccd1 _10102_ sky130_fd_sc_hd__and2_1
X_14293_ _07306_ _06796_ _07303_ _07280_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__or4_4
XFILLER_0_126_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16032_ _09012_ _09110_ _09125_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__a21oi_1
Xhold7490 net4248 vssd1 vssd1 vccd1 vccd1 net8017 sky130_fd_sc_hd__dlygate4sd3_1
X_13244_ _06263_ _06414_ _06306_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o21a_1
X_10456_ net2549 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _06343_ _06345_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__or2_4
XFILLER_0_21_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12126_ _05204_ _05311_ _05313_ _05213_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__o211a_1
X_17983_ _02188_ _02219_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__xor2_1
X_19722_ net7655 net7648 net7673 net4944 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__and4bb_1
X_16934_ _09665_ _09670_ _09955_ vssd1 vssd1 vccd1 vccd1 _09956_ sky130_fd_sc_hd__a21o_1
X_12057_ rbzero.tex_r1\[37\] rbzero.tex_r1\[36\] _05220_ vssd1 vssd1 vccd1 vccd1 _05246_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ net6548 net7101 _04320_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19653_ net6401 net3478 _03429_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__mux2_1
X_16865_ _09475_ _09592_ vssd1 vssd1 vccd1 vccd1 _09887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ _02763_ _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__or2b_1
X_15816_ _08904_ _08910_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19584_ net6482 net3838 net1779 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16796_ net4541 net4630 vssd1 vssd1 vccd1 vccd1 _09825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18535_ net5954 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__clkbuf_1
X_15747_ _08836_ _08841_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__xnor2_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ net3893 _06039_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18466_ net8085 _02643_ net4820 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__or3_1
X_15678_ _08200_ _08280_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17417_ _10433_ _10434_ vssd1 vssd1 vccd1 vccd1 _10435_ sky130_fd_sc_hd__xnor2_1
X_20558__294 clknet_1_1__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__inv_2
X_14629_ _07451_ _07799_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18397_ net5884 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ _10311_ _10366_ vssd1 vssd1 vccd1 vccd1 _10367_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ _10189_ _10191_ _10188_ vssd1 vssd1 vccd1 vccd1 _10298_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19018_ _03080_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20290_ net6409 net4074 _03814_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4105 _09832_ vssd1 vssd1 vccd1 vccd1 net4632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4116 _06096_ vssd1 vssd1 vccd1 vccd1 net4643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4127 net7973 vssd1 vssd1 vccd1 vccd1 net4654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4138 net3392 vssd1 vssd1 vccd1 vccd1 net4665 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3404 net4874 vssd1 vssd1 vccd1 vccd1 net3931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4149 _00432_ vssd1 vssd1 vccd1 vccd1 net4676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3415 _00747_ vssd1 vssd1 vccd1 vccd1 net3942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3426 _01241_ vssd1 vssd1 vccd1 vccd1 net3953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3437 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 net3964 sky130_fd_sc_hd__buf_1
Xhold2703 net3350 vssd1 vssd1 vccd1 vccd1 net3230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3448 net3451 vssd1 vssd1 vccd1 vccd1 net3975 sky130_fd_sc_hd__buf_1
Xhold2714 net5678 vssd1 vssd1 vccd1 vccd1 net3241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3459 _08101_ vssd1 vssd1 vccd1 vccd1 net3986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2725 net7470 vssd1 vssd1 vccd1 vccd1 net3252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2736 net7483 vssd1 vssd1 vccd1 vccd1 net3263 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2747 _03031_ vssd1 vssd1 vccd1 vccd1 net3274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _01143_ vssd1 vssd1 vccd1 vccd1 net3285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2769 net4739 vssd1 vssd1 vccd1 vccd1 net3296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21813_ net255 net2276 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21744_ clknet_leaf_98_i_clk net4827 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21675_ clknet_leaf_124_i_clk net3201 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6030 rbzero.spi_registers.new_texadd\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net6557
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6041 net1629 vssd1 vssd1 vccd1 vccd1 net6568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6052 rbzero.pov.spi_buffer\[60\] vssd1 vssd1 vccd1 vccd1 net6579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11290_ net4862 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__buf_2
Xhold6063 rbzero.tex_g0\[19\] vssd1 vssd1 vccd1 vccd1 net6590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6074 net1785 vssd1 vssd1 vccd1 vccd1 net6601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6085 rbzero.spi_registers.new_vshift\[0\] vssd1 vssd1 vccd1 vccd1 net6612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5340 rbzero.pov.ready_buffer\[68\] vssd1 vssd1 vccd1 vccd1 net5867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6096 net1697 vssd1 vssd1 vccd1 vccd1 net6623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5351 _02971_ vssd1 vssd1 vccd1 vccd1 net5878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5362 net3371 vssd1 vssd1 vccd1 vccd1 net5889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5373 _01179_ vssd1 vssd1 vccd1 vccd1 net5900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5384 net4105 vssd1 vssd1 vccd1 vccd1 net5911 sky130_fd_sc_hd__buf_1
Xhold4650 net783 vssd1 vssd1 vccd1 vccd1 net5177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5395 net3870 vssd1 vssd1 vccd1 vccd1 net5922 sky130_fd_sc_hd__dlygate4sd3_1
X_20386__139 clknet_1_1__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__inv_2
Xhold4661 rbzero.spi_registers.texadd3\[18\] vssd1 vssd1 vccd1 vccd1 net5188 sky130_fd_sc_hd__dlygate4sd3_1
X_22158_ clknet_leaf_88_i_clk net4934 vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4672 net881 vssd1 vssd1 vccd1 vccd1 net5199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4683 net3643 vssd1 vssd1 vccd1 vccd1 net5210 sky130_fd_sc_hd__dlygate4sd3_1
X_21109_ clknet_leaf_94_i_clk net4885 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4694 _00802_ vssd1 vssd1 vccd1 vccd1 net5221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3960 net8186 vssd1 vssd1 vccd1 vccd1 net4487 sky130_fd_sc_hd__dlygate4sd3_1
X_22089_ net151 net2013 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
Xhold3971 net1791 vssd1 vssd1 vccd1 vccd1 net4498 sky130_fd_sc_hd__dlygate4sd3_1
X_14980_ net4520 _08025_ _08079_ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__mux2_1
Xhold3982 _00419_ vssd1 vssd1 vccd1 vccd1 net4509 sky130_fd_sc_hd__dlygate4sd3_1
X_19814__89 clknet_1_1__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__inv_2
Xhold3993 net3727 vssd1 vssd1 vccd1 vccd1 net4520 sky130_fd_sc_hd__clkbuf_2
X_13931_ _06828_ _06850_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16650_ net5949 _09727_ net4134 vssd1 vssd1 vccd1 vccd1 _09731_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13862_ net3579 vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__clkbuf_4
X_15601_ _08686_ _08683_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__or2b_1
X_12813_ _05987_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__nand2_1
X_16581_ _09665_ _09670_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__xor2_2
XFILLER_0_97_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13793_ net575 _06755_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18320_ net4501 net4852 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15532_ _08626_ _08592_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__xnor2_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12744_ _04648_ net4133 _04461_ net4089 net36 _05901_ vssd1 vssd1 vccd1 vccd1 _05921_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _06162_ net3589 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__xnor2_1
X_15463_ _08555_ _08557_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03509_ clknet_0__03509_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03509_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ net31 net30 vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17202_ _08948_ _09970_ _09976_ _08916_ vssd1 vssd1 vccd1 vccd1 _10222_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ _07570_ _07576_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03840_ clknet_0__03840_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03840_
+ sky130_fd_sc_hd__clkbuf_16
X_11626_ _04803_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__xnor2_2
X_18182_ _02245_ _02403_ _02404_ _10133_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15394_ _08427_ _08428_ net8042 _08475_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__nand4_1
XFILLER_0_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17133_ _10030_ _10149_ _10152_ vssd1 vssd1 vccd1 vccd1 _10153_ sky130_fd_sc_hd__o21a_1
Xclkbuf_0__03871_ _03871_ vssd1 vssd1 vccd1 vccd1 clknet_0__03871_ sky130_fd_sc_hd__clkbuf_16
X_14345_ _06832_ _07194_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11557_ _04739_ _04741_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__or3b_1
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ net2791 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__clkbuf_1
X_17064_ _09537_ _09664_ _09967_ vssd1 vssd1 vccd1 vccd1 _10085_ sky130_fd_sc_hd__nor3_1
Xhold609 net5459 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ _07359_ _07366_ _07368_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__o21a_1
X_11488_ net3990 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _09076_ _09078_ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__or2_4
XFILLER_0_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ _06396_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__xnor2_2
X_10439_ net6038 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ net8051 _06006_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__o21ai_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _05297_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17966_ _02078_ _02079_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a21bo_1
X_13089_ _06244_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nand2_1
Xhold1309 rbzero.tex_b0\[0\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16917_ _08661_ _08616_ _09937_ vssd1 vssd1 vccd1 vccd1 _09939_ sky130_fd_sc_hd__o21ai_1
X_19705_ net6070 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__clkbuf_1
X_17897_ _02096_ _02133_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16848_ _09818_ _09577_ vssd1 vssd1 vccd1 vccd1 _09872_ sky130_fd_sc_hd__nand2_1
X_19636_ net1924 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__clkbuf_1
X_19567_ net1998 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
X_16779_ _09809_ _09094_ vssd1 vssd1 vccd1 vccd1 _09810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18518_ net6015 _02693_ _02664_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19498_ _08092_ _03364_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nand2_4
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18449_ _02625_ _02628_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20491__234 clknet_1_0__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__inv_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21460_ clknet_leaf_41_i_clk net1321 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21391_ clknet_leaf_19_i_clk net4978 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20273_ net4071 net4098 _03807_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22012_ net454 net2392 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold3201 net8082 vssd1 vssd1 vccd1 vccd1 net3728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3212 _03095_ vssd1 vssd1 vccd1 vccd1 net3739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3223 net7983 vssd1 vssd1 vccd1 vccd1 net3750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3234 rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 net3761 sky130_fd_sc_hd__clkbuf_2
Xhold2500 _03526_ vssd1 vssd1 vccd1 vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3245 _00746_ vssd1 vssd1 vccd1 vccd1 net3772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2511 net6060 vssd1 vssd1 vccd1 vccd1 net3038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3256 _00521_ vssd1 vssd1 vccd1 vccd1 net3783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2522 _03601_ vssd1 vssd1 vccd1 vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3267 _03105_ vssd1 vssd1 vccd1 vccd1 net3794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 net2940 vssd1 vssd1 vccd1 vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03860_ clknet_0__03860_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03860_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3278 _09789_ vssd1 vssd1 vccd1 vccd1 net3805 sky130_fd_sc_hd__buf_1
Xhold2544 _04274_ vssd1 vssd1 vccd1 vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3289 net2598 vssd1 vssd1 vccd1 vccd1 net3816 sky130_fd_sc_hd__buf_2
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1810 net6899 vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 _00679_ vssd1 vssd1 vccd1 vccd1 net3082 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2566 _04365_ vssd1 vssd1 vccd1 vccd1 net3093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1821 net6901 vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1832 _01314_ vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2577 rbzero.tex_g1\[1\] vssd1 vssd1 vccd1 vccd1 net3104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2588 net5697 vssd1 vssd1 vccd1 vccd1 net3115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1843 net7323 vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1854 net7247 vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2599 _03558_ vssd1 vssd1 vccd1 vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1865 _01499_ vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1876 net7172 vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1887 net6075 vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1898 _01510_ vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10790_ net6458 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkbuf_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21727_ clknet_leaf_102_i_clk net4489 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21658_ clknet_leaf_121_i_clk net3062 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_12460_ net5 _05633_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11411_ net71 _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12391_ _05204_ _05575_ _04955_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__o21a_1
X_21589_ net223 net1501 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_95 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_95/HI o_rgb[2] sky130_fd_sc_hd__conb_1
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14130_ _07245_ _07228_ _07277_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__a21o_1
X_11342_ _04521_ _04531_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ _07191_ _07231_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__xnor2_1
X_11273_ _04461_ _04466_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5170 _04070_ vssd1 vssd1 vccd1 vccd1 net5697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5181 net1439 vssd1 vssd1 vccd1 vccd1 net5708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13012_ _06176_ _06183_ _06186_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__or4b_1
Xhold5192 _04335_ vssd1 vssd1 vccd1 vccd1 net5719 sky130_fd_sc_hd__dlygate4sd3_1
X_17820_ _01956_ _01959_ _01957_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4480 net698 vssd1 vssd1 vccd1 vccd1 net5007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4491 _00855_ vssd1 vssd1 vccd1 vccd1 net5018 sky130_fd_sc_hd__dlygate4sd3_1
X_17751_ _01988_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__nor2_1
Xhold3790 net2711 vssd1 vssd1 vccd1 vccd1 net4317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14963_ _08067_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__buf_4
X_16702_ net1015 _09745_ _09746_ net8002 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a22o_1
X_13914_ _07072_ _07082_ _07084_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__o21a_1
X_17682_ _01920_ _01921_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14894_ rbzero.wall_tracer.visualWallDist\[-9\] _08037_ _08038_ vssd1 vssd1 vccd1
+ vccd1 _08041_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19421_ _08093_ net3671 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__and2_1
X_16633_ _08092_ vssd1 vssd1 vccd1 vccd1 _09721_ sky130_fd_sc_hd__buf_4
X_13845_ _07014_ _07015_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19352_ net5113 _03269_ _03277_ _03275_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16564_ _09527_ _09528_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__and2_1
X_13776_ _06922_ _06946_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__xnor2_1
X_10988_ net7214 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18303_ net6384 net3556 _02493_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
X_15515_ _08602_ _08597_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__or2b_1
XFILLER_0_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19283_ net4842 _03123_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__nand2_4
X_12727_ net35 vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16495_ net4769 _08115_ _09584_ _09585_ _01633_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__o221a_1
X_18234_ net3835 net4524 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__or2_1
X_15446_ _08358_ _08514_ _08515_ _08517_ _08512_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__a32o_1
X_12658_ net25 _05814_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11609_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__inv_2
X_18165_ _02381_ _02387_ net3666 _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15377_ net3453 _08405_ net8501 vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12589_ _05760_ _05768_ net19 vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_170_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ net4657 net4401 vssd1 vssd1 vccd1 vccd1 _10136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03854_ _03854_ vssd1 vssd1 vccd1 vccd1 clknet_0__03854_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _07484_ _07498_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__xor2_4
X_18096_ net3932 net4399 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold406 net6087 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 net5319 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold428 net5347 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _08309_ _09025_ vssd1 vssd1 vccd1 vccd1 _10068_ sky130_fd_sc_hd__nor2_1
Xhold439 _01443_ vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14259_ _07394_ _07409_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ net5988 net5868 _03058_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _00579_ vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 _03367_ vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1128 net3561 vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ _02068_ _02092_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a21o_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 net6563 vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20960_ clknet_leaf_74_i_clk _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19619_ net1248 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
X_20891_ net4928 net63 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21512_ clknet_leaf_12_i_clk net1513 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21443_ clknet_leaf_17_i_clk net3369 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21374_ clknet_leaf_48_i_clk net5398 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20325_ net6136 net3478 _03813_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__mux2_1
Xhold940 _01259_ vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold951 _03414_ vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold962 net6416 vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 net6535 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
X_20256_ net4024 net4103 net4122 _04459_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a31o_1
Xhold984 net6350 vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 _01488_ vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3020 net7721 vssd1 vssd1 vccd1 vccd1 net3547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3031 _00738_ vssd1 vssd1 vccd1 vccd1 net3558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3042 net7736 vssd1 vssd1 vccd1 vccd1 net3569 sky130_fd_sc_hd__dlygate4sd3_1
X_20187_ _05155_ _03744_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__or2_1
Xhold3053 net7642 vssd1 vssd1 vccd1 vccd1 net3580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3064 _02466_ vssd1 vssd1 vccd1 vccd1 net3591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2330 rbzero.tex_g0\[3\] vssd1 vssd1 vccd1 vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3075 net6047 vssd1 vssd1 vccd1 vccd1 net3602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2341 _01336_ vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3086 _00639_ vssd1 vssd1 vccd1 vccd1 net3613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2352 rbzero.tex_r1\[13\] vssd1 vssd1 vccd1 vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3097 net5944 vssd1 vssd1 vccd1 vccd1 net3624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2363 _03602_ vssd1 vssd1 vccd1 vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03843_ clknet_0__03843_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03843_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2374 net7478 vssd1 vssd1 vccd1 vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1640 net6994 vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2385 net7282 vssd1 vssd1 vccd1 vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2396 net7354 vssd1 vssd1 vccd1 vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 _01444_ vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1662 _01484_ vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ rbzero.debug_overlay.facingY\[-8\] _05113_ _05147_ _05148_ vssd1 vssd1 vccd1
+ vccd1 _05149_ sky130_fd_sc_hd__a211o_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1673 net5846 vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1684 net7058 vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_10911_ net6762 net6235 _04265_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1695 _01273_ vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _05074_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nor2_4
XFILLER_0_168_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13630_ _06792_ _06800_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__xnor2_1
X_10842_ net2023 net6034 _04238_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xsplit33 _06533_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13561_ _06683_ _06692_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__xor2_2
X_10773_ net6814 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15300_ _08211_ _08266_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _05691_ net7571 vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16280_ _09274_ _09281_ _09283_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_165_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _06618_ _06634_ net79 net80 _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15231_ _08308_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ net4139 _05627_ _05545_ net4172 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15162_ net3433 _08230_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__nand2_1
X_12374_ _05557_ _05558_ _04949_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _06832_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11325_ rbzero.texu_hot\[4\] _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nand2_1
X_19970_ net6329 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
X_15093_ net3372 _08175_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11256_ net2896 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__clkbuf_1
X_18921_ net7516 net7550 _03025_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
X_14044_ _07168_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11187_ net2842 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__clkbuf_1
X_18852_ net3697 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17803_ _02040_ _02041_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__xor2_2
X_18783_ _02922_ _02923_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__o22ai_1
X_15995_ net5859 net7765 _08111_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__mux2_1
X_17734_ _01971_ _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__xnor2_1
X_14946_ _08070_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17665_ _01903_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__xnor2_1
X_14877_ net4524 _08028_ _07976_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__mux2_1
X_16616_ _09464_ _09573_ _09705_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__a21oi_1
X_19404_ net5500 _03303_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or2_1
X_13828_ _06706_ _06832_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__nor2_1
X_17596_ _01835_ _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ _08338_ _08383_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__nor2_1
X_19335_ net6331 _03237_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13759_ _06719_ _06755_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19266_ net5109 _03216_ _03226_ _03219_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16478_ _09567_ _09568_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__and2b_1
XFILLER_0_183_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7308 net8434 vssd1 vssd1 vccd1 vccd1 net7835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7319 _07924_ vssd1 vssd1 vccd1 vccd1 net7846 sky130_fd_sc_hd__clkbuf_2
X_18217_ net4575 net4428 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15429_ _08522_ _08523_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__xnor2_1
Xhold6607 rbzero.tex_r0\[57\] vssd1 vssd1 vccd1 vccd1 net7134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ net5244 _03182_ _03186_ _03176_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__o211a_1
Xhold6618 net2291 vssd1 vssd1 vccd1 vccd1 net7145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6629 rbzero.tex_b1\[54\] vssd1 vssd1 vccd1 vccd1 net7156 sky130_fd_sc_hd__dlygate4sd3_1
X_18148_ _02373_ _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__or2b_1
Xhold5906 rbzero.spi_registers.new_texadd\[0\]\[12\] vssd1 vssd1 vccd1 vccd1 net6433
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5917 net1353 vssd1 vssd1 vccd1 vccd1 net6444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5928 rbzero.tex_g1\[33\] vssd1 vssd1 vccd1 vccd1 net6455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold203 net5002 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 net5158 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5939 net1450 vssd1 vssd1 vccd1 vccd1 net6466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold225 net5124 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _02314_ net4742 _10260_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_4
Xhold236 net4700 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold247 net5134 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 net5152 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ net6061 _03631_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nor2_1
Xhold269 net5106 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21090_ clknet_leaf_46_i_clk net1421 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20041_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__inv_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21992_ net434 net2124 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ clknet_leaf_70_i_clk net4721 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ net4852 _02508_ _02559_ _04009_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7820 net4639 vssd1 vssd1 vccd1 vccd1 net8347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7831 rbzero.texu_hot\[3\] vssd1 vssd1 vccd1 vccd1 net8358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7842 _06687_ vssd1 vssd1 vccd1 vccd1 net8369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7853 net4439 vssd1 vssd1 vccd1 vccd1 net8380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7864 net4470 vssd1 vssd1 vccd1 vccd1 net8391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21426_ clknet_leaf_40_i_clk net1566 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7875 _08120_ vssd1 vssd1 vccd1 vccd1 net8402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7886 _08156_ vssd1 vssd1 vccd1 vccd1 net8413 sky130_fd_sc_hd__buf_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21357_ clknet_leaf_5_i_clk net5318 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11110_ net6639 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
X_20308_ net1786 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
X_12090_ rbzero.tex_r1\[57\] rbzero.tex_r1\[56\] _05220_ vssd1 vssd1 vccd1 vccd1 _05279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21288_ clknet_leaf_27_i_clk net4395 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold770 _00972_ vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold781 _03458_ vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ net7198 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
Xhold792 net6394 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
X_20239_ net3952 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _01399_ vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2171 net5715 vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
X_20506__247 clknet_1_1__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__inv_2
XFILLER_0_157_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14800_ net4390 _07962_ _07872_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__mux2_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 net7557 vssd1 vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
X_15780_ _08868_ _08873_ _08874_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__a21oi_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2193 _04074_ vssd1 vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ _06162_ net4742 net4762 _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__o22a_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1470 net6799 vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1481 net6771 vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ net7843 _07845_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__or2_1
Xhold1492 _01357_ vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ net4108 _05084_ _05073_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17450_ _10106_ _10351_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nand2_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14662_ _07822_ _07812_ _07826_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__a21o_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11874_ net5205 net5911 _04666_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__or3_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _09350_ _09362_ _09360_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__a21oi_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _06780_ _06783_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and2_1
X_17381_ _09612_ _09249_ vssd1 vssd1 vccd1 vccd1 _10399_ sky130_fd_sc_hd__and2b_1
X_10825_ net6750 net6774 _04227_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ _07753_ _07755_ _07760_ _07763_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19120_ net3996 _05730_ net4097 _03120_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__nand4b_4
X_16332_ _09293_ _09298_ _09423_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__a21o_1
X_13544_ net80 vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__buf_2
X_10756_ _04029_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19051_ net7591 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__clkbuf_1
X_16263_ _09133_ _09354_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13475_ _06472_ _06558_ _06580_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__a21oi_1
X_10687_ net6979 net2728 _04149_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18002_ _02236_ _02237_ net90 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a21oi_2
X_15214_ _08306_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__buf_4
X_12426_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _05258_ vssd1 vssd1 vccd1 vccd1 _05611_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _08401_ _08402_ _09165_ _09170_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15145_ _08148_ _08234_ _08235_ _08239_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__a2bb2o_2
X_12357_ _05040_ _05540_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11308_ _04462_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__buf_4
X_19953_ net3159 net2927 _03583_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__mux2_1
X_15076_ _08169_ _08170_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__nand2_1
X_12288_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _05237_ vssd1 vssd1 vccd1 vccd1 _05474_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14027_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__clkbuf_4
X_18904_ net6512 net1057 _03014_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
X_11239_ net7320 net6215 _04445_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__mux2_1
X_19884_ net3302 net7516 _03550_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ net5879 net1548 net4063 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _09056_ _09072_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__xnor2_2
X_18766_ _02913_ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17717_ net4723 net4520 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__nor2_1
X_14929_ net3875 _08050_ _08052_ net4575 net4719 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18697_ net3678 net4528 _02848_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17648_ _01802_ _01859_ _01887_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a21o_1
X_17579_ _01814_ _01818_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19318_ net1444 _03251_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7105 _02750_ vssd1 vssd1 vccd1 vccd1 net7632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7116 net3580 vssd1 vssd1 vccd1 vccd1 net7643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7127 rbzero.pov.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 net7654 sky130_fd_sc_hd__dlygate4sd3_1
X_19249_ _03202_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__buf_2
XFILLER_0_171_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7138 net3781 vssd1 vssd1 vccd1 vccd1 net7665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6404 rbzero.tex_b0\[9\] vssd1 vssd1 vccd1 vccd1 net6931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7149 net3709 vssd1 vssd1 vccd1 vccd1 net7676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6415 net1773 vssd1 vssd1 vccd1 vccd1 net6942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6426 rbzero.pov.ready_buffer\[25\] vssd1 vssd1 vccd1 vccd1 net6953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20611__342 clknet_1_1__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__inv_2
Xhold6437 _04166_ vssd1 vssd1 vccd1 vccd1 net6964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6448 net2229 vssd1 vssd1 vccd1 vccd1 net6975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5703 rbzero.pov.spi_buffer\[13\] vssd1 vssd1 vccd1 vccd1 net6230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6459 rbzero.tex_b0\[31\] vssd1 vssd1 vccd1 vccd1 net6986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21211_ clknet_leaf_117_i_clk net3325 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5714 net1166 vssd1 vssd1 vccd1 vccd1 net6241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5725 rbzero.spi_registers.new_texadd\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 net6252
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5736 net1247 vssd1 vssd1 vccd1 vccd1 net6263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5747 rbzero.spi_registers.new_texadd\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net6274
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5758 net1377 vssd1 vssd1 vccd1 vccd1 net6285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5769 rbzero.spi_registers.new_texadd\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 net6296
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21142_ clknet_leaf_99_i_clk net3500 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_4
X_21073_ clknet_leaf_75_i_clk _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20024_ net2898 _03609_ net5827 _03316_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21975_ net417 net2246 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer40 _06618_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer51 _06980_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ clknet_leaf_60_i_clk net4545 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ net4219 _04001_ _04002_ _09577_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ net6187 net2247 _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__mux2_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ net2494 _04774_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20788_ _03954_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__nand3_1
XFILLER_0_135_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net6088 net6752 _04075_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7650 _03739_ vssd1 vssd1 vccd1 vccd1 net8177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7661 _08041_ vssd1 vssd1 vccd1 vccd1 net8188 sky130_fd_sc_hd__dlygate4sd3_1
X_13260_ _06385_ _06418_ _06386_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10472_ net2780 net6758 _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7672 rbzero.traced_texa\[8\] vssd1 vssd1 vccd1 vccd1 net8199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7683 _01615_ vssd1 vssd1 vccd1 vccd1 net8210 sky130_fd_sc_hd__dlygate4sd3_1
X_12211_ _05263_ _05385_ _05389_ _05397_ _04817_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__o311a_1
Xhold7694 rbzero.traced_texa\[7\] vssd1 vssd1 vccd1 vccd1 net8221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6960 _04284_ vssd1 vssd1 vccd1 vccd1 net7487 sky130_fd_sc_hd__dlygate4sd3_1
X_21409_ clknet_leaf_36_i_clk net4958 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6971 net3155 vssd1 vssd1 vccd1 vccd1 net7498 sky130_fd_sc_hd__dlygate4sd3_1
X_13191_ _05976_ _05998_ net8051 vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__a21o_1
Xhold6982 rbzero.pov.spi_buffer\[72\] vssd1 vssd1 vccd1 vccd1 net7509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6993 net3286 vssd1 vssd1 vccd1 vccd1 net7520 sky130_fd_sc_hd__dlygate4sd3_1
X_12142_ _04847_ _05327_ _05329_ _04829_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12073_ _04943_ _05259_ _05261_ _04947_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__o211a_1
X_16950_ net4877 _08494_ _09673_ _09971_ vssd1 vssd1 vccd1 vccd1 _09972_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11024_ net2668 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
X_15901_ _06122_ net4918 vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__nor2_2
X_16881_ _09901_ _09902_ vssd1 vssd1 vccd1 vccd1 _09903_ sky130_fd_sc_hd__nor2_1
X_15832_ _08925_ _08926_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__nor2_1
X_18620_ net4635 _02770_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__nand2_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _08854_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__and2_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ net7635 _02720_ _02245_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12975_ net4347 net3999 vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__xnor2_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17502_ _01741_ _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nor2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14714_ net7795 _07853_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _02658_ _02659_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__nand2_1
X_11926_ net4118 _05094_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__nor2_1
X_15694_ _08716_ _08718_ _08717_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__a21o_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _01663_ _01673_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__or2_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14645_ _07511_ _07787_ _07803_ _07815_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__o31a_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _04664_ _04660_ net4162 net4139 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__o31ai_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ net7250 net7429 _04216_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__mux2_1
X_17364_ _10382_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__clkbuf_1
X_14576_ _07740_ _07746_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11788_ _04835_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16315_ _09405_ _09406_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19103_ net2709 _03126_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__or2_1
X_13527_ _06697_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__buf_2
X_17295_ _10210_ _10216_ vssd1 vssd1 vccd1 vccd1 _10314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ net6912 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19034_ net3403 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__clkbuf_1
X_16246_ _09123_ _09121_ _09243_ _09337_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_126_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13458_ _06498_ _06558_ _06594_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12409_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _05369_ vssd1 vssd1 vccd1 vccd1 _05594_
+ sky130_fd_sc_hd__mux2_1
X_16177_ _09248_ _09269_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ _06441_ _06558_ _06559_ _06550_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4309 _00963_ vssd1 vssd1 vccd1 vccd1 net4836 sky130_fd_sc_hd__dlygate4sd3_1
X_15128_ _07938_ net8393 _08113_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__mux2_2
XFILLER_0_142_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3608 _09731_ vssd1 vssd1 vccd1 vccd1 net4135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3619 _05049_ vssd1 vssd1 vccd1 vccd1 net4146 sky130_fd_sc_hd__dlygate4sd3_1
X_19936_ net7560 net3312 _03572_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
X_15059_ _06361_ _06314_ net8411 vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__nor3_1
Xhold2907 net4329 vssd1 vssd1 vccd1 vccd1 net3434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2918 net8224 vssd1 vssd1 vccd1 vccd1 net3445 sky130_fd_sc_hd__clkbuf_4
Xhold2929 net4839 vssd1 vssd1 vccd1 vccd1 net3456 sky130_fd_sc_hd__dlygate4sd3_1
X_19867_ net7443 net6512 _03539_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18818_ net5845 _02960_ _02961_ _02962_ net1547 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18749_ _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21760_ clknet_leaf_111_i_clk net7683 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20711_ _03889_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21691_ clknet_leaf_114_i_clk net4457 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6201 _03450_ vssd1 vssd1 vccd1 vccd1 net6728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6212 net2146 vssd1 vssd1 vccd1 vccd1 net6739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6223 net2029 vssd1 vssd1 vccd1 vccd1 net6750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6234 rbzero.tex_g0\[39\] vssd1 vssd1 vccd1 vccd1 net6761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5500 _04393_ vssd1 vssd1 vccd1 vccd1 net6027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6245 net2008 vssd1 vssd1 vccd1 vccd1 net6772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5511 net3641 vssd1 vssd1 vccd1 vccd1 net6038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6256 rbzero.tex_g1\[27\] vssd1 vssd1 vccd1 vccd1 net6783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6267 net2183 vssd1 vssd1 vccd1 vccd1 net6794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5522 rbzero.spi_registers.new_floor\[1\] vssd1 vssd1 vccd1 vccd1 net6049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6278 _04396_ vssd1 vssd1 vccd1 vccd1 net6805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5533 rbzero.pov.ready_buffer\[57\] vssd1 vssd1 vccd1 vccd1 net6060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5544 rbzero.tex_g0\[32\] vssd1 vssd1 vccd1 vccd1 net6071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6289 net636 vssd1 vssd1 vccd1 vccd1 net6816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4810 _00803_ vssd1 vssd1 vccd1 vccd1 net5337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5555 net1591 vssd1 vssd1 vccd1 vccd1 net6082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5566 _04260_ vssd1 vssd1 vccd1 vccd1 net6093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4821 net955 vssd1 vssd1 vccd1 vccd1 net5348 sky130_fd_sc_hd__dlygate4sd3_1
X_22174_ clknet_leaf_68_i_clk net4938 vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4832 rbzero.spi_registers.texadd3\[5\] vssd1 vssd1 vccd1 vccd1 net5359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5577 _04404_ vssd1 vssd1 vccd1 vccd1 net6104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5588 _04206_ vssd1 vssd1 vccd1 vccd1 net6115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4843 net947 vssd1 vssd1 vccd1 vccd1 net5370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4854 _01604_ vssd1 vssd1 vccd1 vccd1 net5381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5599 _03540_ vssd1 vssd1 vccd1 vccd1 net6126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4865 net951 vssd1 vssd1 vccd1 vccd1 net5392 sky130_fd_sc_hd__dlygate4sd3_1
X_21125_ clknet_leaf_33_i_clk net3895 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_1
Xhold4876 rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 net5403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4887 net990 vssd1 vssd1 vccd1 vccd1 net5414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4898 _00818_ vssd1 vssd1 vccd1 vccd1 net5425 sky130_fd_sc_hd__dlygate4sd3_1
X_21056_ clknet_leaf_73_i_clk _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_20007_ net5887 _03607_ _03621_ _03339_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ net4147 _05912_ _05935_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a211o_1
X_21958_ net400 net2535 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ net4145 _04887_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20909_ clknet_leaf_81_i_clk _00396_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12691_ net6111 _05853_ _05863_ net54 vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a22o_1
X_21889_ net331 net3178 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20618__348 clknet_1_1__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__inv_2
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _07584_ _07599_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11642_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__buf_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14361_ _07482_ _07499_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ net2753 _04761_ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16100_ _09192_ _09193_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__and2b_1
Xinput18 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
X_13312_ _06459_ _06479_ _06480_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__a31o_1
X_17080_ _10097_ _10100_ vssd1 vssd1 vccd1 vccd1 _10101_ sky130_fd_sc_hd__xor2_1
X_10524_ net5547 net5696 _04064_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__mux2_1
Xinput29 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14292_ _07394_ _07462_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__nand2_1
X_16031_ _09121_ _09124_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__xor2_1
Xhold7480 net4737 vssd1 vssd1 vccd1 vccd1 net8007 sky130_fd_sc_hd__buf_1
X_13243_ net7837 _06266_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__nor2_1
X_10455_ net6940 net7121 _04031_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__mux2_1
Xhold7491 net4550 vssd1 vssd1 vccd1 vccd1 net8018 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6790 _04292_ vssd1 vssd1 vccd1 vccd1 net7317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ rbzero.wall_tracer.rayAddendX\[-2\] _06344_ _06305_ vssd1 vssd1 vccd1 vccd1
+ _06345_ sky130_fd_sc_hd__mux2_4
XFILLER_0_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ _04921_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _02217_ _02218_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__nor2_1
X_19721_ net973 net7273 net3703 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a21o_1
X_12056_ rbzero.tex_r1\[39\] rbzero.tex_r1\[38\] _04838_ vssd1 vssd1 vccd1 vccd1 _05245_
+ sky130_fd_sc_hd__mux2_1
X_16933_ _09668_ _09669_ vssd1 vssd1 vccd1 vccd1 _09955_ sky130_fd_sc_hd__and2b_1
XFILLER_0_205_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20363__118 clknet_1_0__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__inv_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ net3164 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
X_19652_ net6518 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16864_ _09876_ _09878_ _09883_ _09884_ vssd1 vssd1 vccd1 vccd1 _09886_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ net3619 net1002 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__nand2_1
X_15815_ _08906_ _08908_ _08909_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a21o_1
X_16795_ net4541 net4630 vssd1 vssd1 vccd1 vccd1 _09824_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19583_ net6289 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15746_ _08204_ _08573_ _08837_ _08838_ _08840_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__a32o_1
X_18534_ net5952 _02707_ _02664_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12958_ net3965 net3999 _06060_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__and3_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11909_ _04465_ _05083_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nand2_2
XFILLER_0_185_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15677_ _08245_ _08433_ _08770_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__a31o_1
X_18465_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _02617_
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _04686_ net3964 _06030_ net3469 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17416_ _10062_ _08461_ vssd1 vssd1 vccd1 vccd1 _10434_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14628_ _07796_ _07798_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18396_ rbzero.wall_tracer.rayAddendX\[0\] _02579_ _02537_ vssd1 vssd1 vccd1 vccd1
+ _02580_ sky130_fd_sc_hd__mux2_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17347_ _10364_ _10365_ vssd1 vssd1 vccd1 vccd1 _10366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14559_ _07726_ _07729_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17278_ _10295_ _10296_ vssd1 vssd1 vccd1 vccd1 _10297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16229_ _09217_ _09320_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19017_ net3899 net4030 _03078_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4106 _09840_ vssd1 vssd1 vccd1 vccd1 net4633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4117 _06102_ vssd1 vssd1 vccd1 vccd1 net4644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4128 net3855 vssd1 vssd1 vccd1 vccd1 net4655 sky130_fd_sc_hd__clkbuf_2
Xhold4139 net8344 vssd1 vssd1 vccd1 vccd1 net4666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3405 net3729 vssd1 vssd1 vccd1 vccd1 net3932 sky130_fd_sc_hd__clkbuf_2
Xhold3416 net8274 vssd1 vssd1 vccd1 vccd1 net3943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3427 net7677 vssd1 vssd1 vccd1 vccd1 net3954 sky130_fd_sc_hd__clkbuf_2
Xhold3438 _06107_ vssd1 vssd1 vccd1 vccd1 net3965 sky130_fd_sc_hd__clkbuf_4
Xhold2704 _03520_ vssd1 vssd1 vccd1 vccd1 net3231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3449 _04474_ vssd1 vssd1 vccd1 vccd1 net3976 sky130_fd_sc_hd__buf_2
Xhold2715 _01572_ vssd1 vssd1 vccd1 vccd1 net3242 sky130_fd_sc_hd__dlygate4sd3_1
X_19919_ net6744 net2801 _03561_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__mux2_1
Xhold2726 _03044_ vssd1 vssd1 vccd1 vccd1 net3253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2737 _04288_ vssd1 vssd1 vccd1 vccd1 net3264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2748 _00681_ vssd1 vssd1 vccd1 vccd1 net3275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2759 net7519 vssd1 vssd1 vccd1 vccd1 net3286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21812_ net254 net3094 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_127_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21743_ clknet_leaf_99_i_clk net4593 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21674_ clknet_leaf_124_i_clk net1810 vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6020 rbzero.tex_b1\[56\] vssd1 vssd1 vccd1 vccd1 net6547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6031 net1859 vssd1 vssd1 vccd1 vccd1 net6558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6042 rbzero.spi_registers.new_texadd\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net6569
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6053 rbzero.tex_r1\[60\] vssd1 vssd1 vccd1 vccd1 net6580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6064 net1739 vssd1 vssd1 vccd1 vccd1 net6591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5330 _00631_ vssd1 vssd1 vccd1 vccd1 net5857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6075 rbzero.spi_registers.new_texadd\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net6602
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6086 net1033 vssd1 vssd1 vccd1 vccd1 net6613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5341 net3279 vssd1 vssd1 vccd1 vccd1 net5868 sky130_fd_sc_hd__buf_1
Xhold6097 _03476_ vssd1 vssd1 vccd1 vccd1 net6624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5352 _02976_ vssd1 vssd1 vccd1 vccd1 net5879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5374 net3432 vssd1 vssd1 vccd1 vccd1 net5901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4640 net908 vssd1 vssd1 vccd1 vccd1 net5167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5385 _05067_ vssd1 vssd1 vccd1 vccd1 net5912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4651 _00846_ vssd1 vssd1 vccd1 vccd1 net5178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22157_ clknet_leaf_55_i_clk _01644_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5396 _03989_ vssd1 vssd1 vccd1 vccd1 net5923 sky130_fd_sc_hd__buf_1
Xhold4662 net882 vssd1 vssd1 vccd1 vccd1 net5189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4673 rbzero.spi_registers.texadd2\[4\] vssd1 vssd1 vccd1 vccd1 net5200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4684 rbzero.spi_registers.texadd0\[10\] vssd1 vssd1 vccd1 vccd1 net5211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4695 net928 vssd1 vssd1 vccd1 vccd1 net5222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3950 net8184 vssd1 vssd1 vccd1 vccd1 net4477 sky130_fd_sc_hd__dlygate4sd3_1
X_21108_ clknet_leaf_17_i_clk net1391 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3961 _01214_ vssd1 vssd1 vccd1 vccd1 net4488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22088_ net150 net2659 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3972 net7947 vssd1 vssd1 vccd1 vccd1 net4499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3983 net3410 vssd1 vssd1 vccd1 vccd1 net4510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _06851_ _06862_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__nor2_1
Xhold3994 net7874 vssd1 vssd1 vccd1 vccd1 net4521 sky130_fd_sc_hd__dlygate4sd3_1
X_21039_ clknet_leaf_56_i_clk net5724 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ net536 _07031_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15600_ _08685_ _08684_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__or2b_1
X_12812_ _05986_ _05982_ _05980_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nand3b_1
X_16580_ _09668_ _09669_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__xnor2_2
X_13792_ _06933_ _06932_ _06930_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a21o_1
X_15531_ _08593_ _08586_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ net37 net36 _05914_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__o31a_2
XFILLER_0_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_91_i_clk clknet_4_7__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18250_ net3588 _02460_ _02457_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a21bo_1
X_15462_ _08280_ _08323_ _08524_ _08556_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__o31a_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12674_ _05850_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__03508_ clknet_0__03508_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03508_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _09537_ _10220_ vssd1 vssd1 vccd1 vccd1 _10221_ sky130_fd_sc_hd__nor2_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _07536_ _07547_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__xnor2_2
X_11625_ _04804_ _04769_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and2b_1
X_18181_ _02401_ _02402_ _02396_ _02398_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15393_ _08403_ _08458_ _08477_ _08476_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__or4b_1
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17132_ _10028_ _10151_ vssd1 vssd1 vccd1 vccd1 _10152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03870_ _03870_ vssd1 vssd1 vccd1 vccd1 clknet_0__03870_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ _07306_ _07281_ _07513_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_108_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11556_ _04742_ _04467_ _04744_ _04022_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__o221a_1
X_17063_ _09965_ _09966_ vssd1 vssd1 vccd1 vccd1 _10084_ sky130_fd_sc_hd__and2_1
X_10507_ net6999 net2790 _04053_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14275_ _07441_ _07445_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ net3443 _04464_ _04501_ net3431 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a22o_1
X_16014_ _08992_ _09083_ _09081_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__a21bo_1
X_13226_ _06378_ _06367_ _06385_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ net4268 rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__or2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ reg_rgb\[7\] _05296_ _05054_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__mux2_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _01784_ _09410_ _02076_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__or3_1
X_13088_ net5408 _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__xnor2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19704_ net6068 net3478 _03456_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16916_ _08661_ _08616_ _09937_ vssd1 vssd1 vccd1 vccd1 _09938_ sky130_fd_sc_hd__or3_1
X_12039_ _05204_ _05225_ _05227_ _04955_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17896_ _02096_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_44_i_clk clknet_4_9__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19635_ net6647 net3745 _03441_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__mux2_1
X_16847_ net3799 _09867_ _09868_ _06057_ vssd1 vssd1 vccd1 vccd1 _09871_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19566_ net6800 net1396 _03403_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
X_16778_ _08103_ vssd1 vssd1 vccd1 vccd1 _09809_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18517_ _02684_ _02685_ _02691_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_193_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15729_ _08821_ _08822_ _08823_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19497_ _03344_ _03363_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_59_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18448_ _02627_ rbzero.wall_tracer.rayAddendX\[3\] _02623_ vssd1 vssd1 vccd1 vccd1
+ _02628_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18379_ net8048 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21390_ clknet_leaf_21_i_clk net5274 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20272_ _03689_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22011_ net453 net1208 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3202 net4875 vssd1 vssd1 vccd1 vccd1 net3729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3213 _00736_ vssd1 vssd1 vccd1 vccd1 net3740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3224 net2196 vssd1 vssd1 vccd1 vccd1 net3751 sky130_fd_sc_hd__clkbuf_2
Xhold3235 _02918_ vssd1 vssd1 vccd1 vccd1 net3762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2501 _01094_ vssd1 vssd1 vccd1 vccd1 net3028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3246 net4082 vssd1 vssd1 vccd1 vccd1 net3773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2512 _03056_ vssd1 vssd1 vccd1 vccd1 net3039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3257 net4898 vssd1 vssd1 vccd1 vccd1 net3784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 _01163_ vssd1 vssd1 vccd1 vccd1 net3050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3268 _00745_ vssd1 vssd1 vccd1 vccd1 net3795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3279 net7962 vssd1 vssd1 vccd1 vccd1 net3806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 _03582_ vssd1 vssd1 vccd1 vccd1 net3061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1800 net7066 vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2545 _01381_ vssd1 vssd1 vccd1 vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1811 _01539_ vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2556 net4831 vssd1 vssd1 vccd1 vccd1 net3083 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1822 _04037_ vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2567 _01299_ vssd1 vssd1 vccd1 vccd1 net3094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 net2647 vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 net5701 vssd1 vssd1 vccd1 vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2589 _01562_ vssd1 vssd1 vccd1 vccd1 net3116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _04092_ vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1855 _04417_ vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1866 net3066 vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1877 _01427_ vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1888 net6077 vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1899 net4900 vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21726_ clknet_leaf_102_i_clk net4469 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21657_ clknet_leaf_121_i_clk net2862 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ _04500_ _04501_ _04599_ _04601_ _04466_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__o32a_1
XFILLER_0_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _04838_ vssd1 vssd1 vccd1 vccd1 _05575_
+ sky130_fd_sc_hd__mux2_1
X_21588_ net222 net2989 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_96 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_96/HI o_rgb[3] sky130_fd_sc_hd__conb_1
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11341_ _04519_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14060_ _07200_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__xor2_2
X_11272_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__buf_4
Xhold5160 rbzero.tex_r0\[11\] vssd1 vssd1 vccd1 vccd1 net5687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ net4506 _06175_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__or2_1
Xhold5171 net3115 vssd1 vssd1 vccd1 vccd1 net5698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5182 rbzero.pov.spi_buffer\[50\] vssd1 vssd1 vccd1 vccd1 net5709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5193 net2991 vssd1 vssd1 vccd1 vccd1 net5720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4470 net670 vssd1 vssd1 vccd1 vccd1 net4997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4481 rbzero.spi_registers.texadd3\[11\] vssd1 vssd1 vccd1 vccd1 net5008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4492 net686 vssd1 vssd1 vccd1 vccd1 net5019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3780 _00764_ vssd1 vssd1 vccd1 vccd1 net4307 sky130_fd_sc_hd__dlygate4sd3_1
X_17750_ _01896_ _01900_ _01987_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__and3_1
X_14962_ _08078_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__clkbuf_1
X_16701_ net969 _09745_ _09746_ net8015 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__a22o_1
X_13913_ _07061_ _07083_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__or2b_1
X_17681_ _08918_ _10211_ _01693_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a21oi_1
X_14893_ net4506 _08034_ _08036_ net4518 net4679 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19420_ net1724 net3670 _03310_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__mux2_1
X_13844_ _07009_ _07013_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__xnor2_1
X_16632_ _04021_ net4124 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19351_ net6510 _03271_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__or2_1
X_16563_ _09634_ _09652_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13775_ _06707_ _06925_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10987_ net2857 net7212 _04309_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__mux2_1
X_20475__219 clknet_1_1__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__inv_2
X_18302_ net6382 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__clkbuf_1
X_15514_ _08601_ _08599_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__or2b_1
X_12726_ net37 net36 _05900_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or4b_1
XFILLER_0_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19282_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__clkbuf_4
X_16494_ _09581_ _09583_ net3454 vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _08526_ _08527_ _08539_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18233_ _02449_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__clkbuf_1
X_12657_ _05814_ _05833_ _05834_ _05835_ net27 vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11608_ _04781_ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ _08456_ _08466_ _08459_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__a21o_1
X_18164_ net3790 net3777 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12588_ net51 net41 net40 _05203_ _05747_ _05749_ vssd1 vssd1 vccd1 vccd1 _05768_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03853_ _03853_ vssd1 vssd1 vccd1 vccd1 clknet_0__03853_ sky130_fd_sc_hd__clkbuf_16
X_17115_ _10135_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14327_ _07485_ _07496_ _07497_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18095_ net3700 _02324_ _02323_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__o21a_1
X_11539_ net4127 net4366 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold407 net6089 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 net5321 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ _10065_ _10066_ vssd1 vssd1 vccd1 vccd1 _10067_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold429 net5349 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ _07385_ _07428_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20369__124 clknet_1_1__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__inv_2
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13209_ _06266_ _05987_ _05988_ _06379_ net8217 vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__a311o_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _07342_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ net1704 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1107 net5499 vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _00919_ vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ _02162_ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__xnor2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 _03417_ vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17879_ _02115_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19618_ net6263 net1426 _03430_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20890_ _03312_ net679 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19549_ net1743 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21511_ clknet_leaf_12_i_clk net1554 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21442_ clknet_leaf_26_i_clk net1702 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21373_ clknet_leaf_44_i_clk net5362 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20324_ net6685 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold930 _02496_ vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 net6314 vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold952 _00955_ vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _03469_ vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20255_ net4103 _03794_ net6001 _03765_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold974 _01076_ vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3010 net5819 vssd1 vssd1 vccd1 vccd1 net3537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 net6352 vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3021 _03327_ vssd1 vssd1 vccd1 vccd1 net3548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 net6206 vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3032 net4873 vssd1 vssd1 vccd1 vccd1 net3559 sky130_fd_sc_hd__dlygate4sd3_1
X_20580__314 clknet_1_1__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__inv_2
X_20186_ net3567 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
Xhold3043 _03313_ vssd1 vssd1 vccd1 vccd1 net3570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3054 _03736_ vssd1 vssd1 vccd1 vccd1 net3581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2320 _01341_ vssd1 vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3065 net7620 vssd1 vssd1 vccd1 vccd1 net3592 sky130_fd_sc_hd__buf_2
Xhold2331 net7213 vssd1 vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3076 _00637_ vssd1 vssd1 vccd1 vccd1 net3603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2342 net7541 vssd1 vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3087 rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 net3614 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2353 net2767 vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3098 _00935_ vssd1 vssd1 vccd1 vccd1 net3625 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03842_ clknet_0__03842_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03842_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2364 _01164_ vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2375 _01389_ vssd1 vssd1 vccd1 vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1630 _01500_ vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1641 net6996 vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 _01033_ vssd1 vssd1 vccd1 vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2397 _04257_ vssd1 vssd1 vccd1 vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1652 net3172 vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1663 net7174 vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1674 net7134 vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1685 net7060 vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_10910_ net3071 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1696 net6959 vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _05070_ _05077_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__a21o_4
XFILLER_0_168_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _04193_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xsplit23 _06503_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_1
X_13560_ _06721_ _06728_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_17_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xsplit34 _06531_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10772_ net2533 net6812 _04194_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _05691_ net4156 vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21709_ clknet_leaf_119_i_clk net3471 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13491_ _06658_ _06659_ _06632_ _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__o2bb2a_2
X_15230_ _08311_ _08324_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ _04706_ _05625_ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15161_ net3433 _08230_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__or2_2
X_12373_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _05250_ vssd1 vssd1 vccd1 vccd1 _05558_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14112_ _07241_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__nor2_2
XFILLER_0_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ rbzero.spi_registers.texadd3\[10\] rbzero.spi_registers.texadd1\[10\] rbzero.spi_registers.texadd0\[10\]
+ rbzero.spi_registers.texadd2\[10\] _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04516_
+ sky130_fd_sc_hd__mux4_2
X_15092_ _08161_ _08168_ _08180_ _08186_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18920_ net3208 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
X_14043_ _07212_ _07213_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__xor2_1
X_11255_ net7375 net5626 _04445_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__mux2_1
X_18851_ _02969_ net3696 _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__and3_1
X_11186_ net7147 net7089 _04412_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17802_ _01891_ _01934_ _01932_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18782_ _02914_ _02924_ _02928_ _04480_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a31o_1
X_15994_ _08989_ _08991_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__xor2_4
X_17733_ _10163_ net4908 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__nor2_1
X_14945_ net4535 _07892_ _08068_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _10327_ _10220_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__nor2_1
X_14876_ net7794 _07979_ _08027_ _08020_ _07869_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__a221o_1
X_19403_ net5484 _03302_ _03306_ _03299_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__o211a_1
X_16615_ _09570_ _09572_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__nor2_1
X_13827_ _06956_ _06957_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__xnor2_1
X_17595_ _10392_ _01713_ _01711_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a21oi_1
X_19334_ net5304 _03235_ _03265_ _03259_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__o211a_1
X_16546_ _08323_ _08418_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__or2_2
X_13758_ _06889_ _06888_ _06887_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12709_ net43 _05852_ _05864_ net44 _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a221o_1
X_19265_ net6623 _03217_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__or2_1
X_16477_ _09565_ _09566_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__nand2_1
X_13689_ _06855_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__xnor2_1
Xhold7309 _08668_ vssd1 vssd1 vccd1 vccd1 net7836 sky130_fd_sc_hd__buf_2
XFILLER_0_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18216_ net4575 net4428 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nor2_1
X_15428_ _08255_ _08306_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19196_ net6434 _03183_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__or2_1
Xhold6608 net2201 vssd1 vssd1 vccd1 vccd1 net7135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6619 rbzero.tex_b0\[36\] vssd1 vssd1 vccd1 vccd1 net7146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15359_ _08428_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__inv_2
X_18147_ net3785 net4390 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__nand2_1
Xhold5907 net1483 vssd1 vssd1 vccd1 vccd1 net6434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5918 rbzero.spi_registers.new_texadd\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net6445
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5929 net1313 vssd1 vssd1 vccd1 vccd1 net6456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 net5120 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold215 net5100 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 net5126 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _02250_ _02251_ _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold237 net5148 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold248 net7082 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _09908_ _09920_ _09918_ vssd1 vssd1 vccd1 vccd1 _10050_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold259 net5154 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ net3431 _03642_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21991_ net433 net2145 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ clknet_leaf_70_i_clk net4754 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_20423__173 clknet_1_0__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__inv_2
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _02517_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7810 net4621 vssd1 vssd1 vccd1 vccd1 net8337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7821 rbzero.wall_tracer.stepDistY\[-2\] vssd1 vssd1 vccd1 vccd1 net8348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7832 net3501 vssd1 vssd1 vccd1 vccd1 net8359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7843 net7783 vssd1 vssd1 vccd1 vccd1 net8370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7854 rbzero.wall_tracer.stepDistX\[-1\] vssd1 vssd1 vccd1 vccd1 net8381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21425_ clknet_leaf_35_i_clk net1595 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7876 net4895 vssd1 vssd1 vccd1 vccd1 net8403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7887 _08209_ vssd1 vssd1 vccd1 vccd1 net8414 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7898 _08193_ vssd1 vssd1 vccd1 vccd1 net8425 sky130_fd_sc_hd__buf_1
X_21356_ clknet_leaf_8_i_clk net5302 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20307_ net6601 net3745 _03825_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__mux2_1
X_21287_ clknet_leaf_27_i_clk net4368 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold760 _02478_ vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 net6344 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold782 _00990_ vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net2777 net7196 _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__mux2_1
X_20238_ _02993_ net3951 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and2_1
Xhold793 net6396 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ rbzero.debug_overlay.facingY\[-3\] _03711_ vssd1 vssd1 vccd1 vccd1 _03740_
+ sky130_fd_sc_hd__or2_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2150 _04121_ vssd1 vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 net7122 vssd1 vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2172 _01342_ vssd1 vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2183 _03130_ vssd1 vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12991_ net3926 vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__inv_2
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _01558_ vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1460 _01432_ vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11942_ _05100_ _05109_ _05110_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__or3_1
X_14730_ _07821_ _07830_ _07839_ net7811 vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__a211o_1
Xhold1471 _03405_ vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1482 _04192_ vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 net6871 vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _07511_ _07787_ _07803_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__or4_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11873_ _04667_ net4116 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__or2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _09478_ _09490_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20398__150 clknet_1_1__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__inv_2
X_13612_ _06780_ _06781_ _06782_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__nand3_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ net2784 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__clkbuf_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _10395_ _10396_ _10397_ vssd1 vssd1 vccd1 vccd1 _10398_ sky130_fd_sc_hd__a21oi_1
X_14592_ net77 _07146_ _07756_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__and3_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16331_ _09177_ _09297_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13543_ _06708_ _06695_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or2_1
X_10755_ net2009 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _06122_ _09060_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__nor2_2
X_19050_ net7589 net3674 net3398 vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
X_13474_ _06441_ _06558_ _06559_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o21a_1
X_10686_ net2451 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15213_ _08294_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18001_ _02236_ _02237_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__or2_1
X_12425_ _04943_ _05609_ _04947_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__o21a_1
X_16193_ _08666_ _08430_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15144_ _08156_ _08238_ _06118_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12356_ _04706_ _04750_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__or3b_1
XFILLER_0_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ _04494_ _04496_ _04497_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__a22o_1
X_19952_ net2713 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
X_15075_ net3536 net4168 net3348 vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12287_ _05465_ _05468_ _05472_ _04942_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a211o_1
X_14026_ _07148_ _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__nand2_2
X_18903_ net7445 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
X_11238_ net7283 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__clkbuf_1
X_19883_ net3303 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
X_18834_ net1547 _02973_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nand2_1
X_11169_ net7447 net7417 _04401_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _02865_ net3678 net4560 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__or3b_2
X_15977_ _09070_ _09071_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ _01955_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14928_ net8264 _06237_ _04482_ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__o21a_1
X_18696_ net3678 net4528 _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _01871_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14859_ net8491 _07934_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19783__62 clknet_1_1__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17578_ _01814_ _01818_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19317_ net5456 _03250_ _03256_ _03246_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16529_ _09506_ _09617_ _09618_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7106 net3885 vssd1 vssd1 vccd1 vccd1 net7633 sky130_fd_sc_hd__dlygate4sd3_1
X_19248_ _03200_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7128 net3823 vssd1 vssd1 vccd1 vccd1 net7655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7139 _09748_ vssd1 vssd1 vccd1 vccd1 net7666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6405 net2072 vssd1 vssd1 vccd1 vccd1 net6932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6416 _04422_ vssd1 vssd1 vccd1 vccd1 net6943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19179_ net5081 _03168_ _03175_ _03176_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__o211a_1
Xhold6427 net2485 vssd1 vssd1 vccd1 vccd1 net6954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6438 net2144 vssd1 vssd1 vccd1 vccd1 net6965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20453__199 clknet_1_1__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__inv_2
Xhold6449 _04052_ vssd1 vssd1 vccd1 vccd1 net6976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5704 net1168 vssd1 vssd1 vccd1 vccd1 net6231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5715 rbzero.tex_g1\[46\] vssd1 vssd1 vccd1 vccd1 net6242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21210_ clknet_leaf_117_i_clk net2195 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5726 net1211 vssd1 vssd1 vccd1 vccd1 net6253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5737 rbzero.spi_registers.new_texadd\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net6264
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5748 net1340 vssd1 vssd1 vccd1 vccd1 net6275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5759 rbzero.spi_registers.new_mapd\[9\] vssd1 vssd1 vccd1 vccd1 net6286 sky130_fd_sc_hd__dlygate4sd3_1
X_21141_ clknet_leaf_99_i_clk net4774 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21072_ clknet_leaf_78_i_clk _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20023_ net5826 _03631_ _03606_ _03632_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21974_ net416 net2702 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer30 _06900_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer41 net567 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer52 _06694_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ clknet_leaf_88_i_clk _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20856_ net4215 _04001_ _04002_ _09450_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a22o_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20787_ _03954_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10540_ net1992 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7640 rbzero.map_overlay.i_mapdy\[1\] vssd1 vssd1 vccd1 vccd1 net8167 sky130_fd_sc_hd__dlygate4sd3_1
X_10471_ _04030_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7673 _03982_ vssd1 vssd1 vccd1 vccd1 net8200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12210_ _04947_ _05392_ _05394_ _05396_ net84 vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21408_ clknet_leaf_36_i_clk net3647 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6950 net2900 vssd1 vssd1 vccd1 vccd1 net7477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7695 _03974_ vssd1 vssd1 vccd1 vccd1 net8222 sky130_fd_sc_hd__dlygate4sd3_1
X_13190_ _06359_ _06360_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__xnor2_2
Xhold6961 net3108 vssd1 vssd1 vccd1 vccd1 net7488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6972 rbzero.tex_g0\[47\] vssd1 vssd1 vccd1 vccd1 net7499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6983 net1869 vssd1 vssd1 vccd1 vccd1 net7510 sky130_fd_sc_hd__dlygate4sd3_1
X_12141_ _04832_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__or2_1
Xhold6994 rbzero.spi_registers.new_mapd\[6\] vssd1 vssd1 vccd1 vccd1 net7521 sky130_fd_sc_hd__dlygate4sd3_1
X_21339_ clknet_leaf_6_i_clk net5414 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ _04930_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold590 _01544_ vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net5718 net7451 _04331_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__mux2_1
X_15900_ _08131_ _08277_ _08142_ _08253_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__or4b_1
X_16880_ _09479_ _09603_ _09605_ vssd1 vssd1 vccd1 vccd1 _09902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15831_ _08924_ _08914_ _08923_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__and3_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_15__f_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _06046_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__xnor2_1
X_15762_ _08808_ _08813_ _08853_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__a21o_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ net1817 _06061_ _06043_ net4324 _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a221oi_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17501_ _10425_ _01739_ _01740_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__and3_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 net8162 vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__clkbuf_2
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ net7811 _07881_ _07882_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__or3_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _02626_ net4698 net3494 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__or3b_1
X_11925_ _05107_ _05077_ net4108 _05091_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__and4_4
X_15693_ _08773_ _08776_ _08775_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__a21bo_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _01663_ _01673_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nand2_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _07790_ _07788_ _07802_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__o21ai_1
X_11856_ _04658_ net4161 _05044_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__and4b_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10807_ net6645 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17363_ _10381_ net4610 _10260_ vssd1 vssd1 vccd1 vccd1 _10382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14575_ _07741_ _07744_ _07745_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__a21boi_1
X_11787_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19102_ net4309 _03125_ net3036 _03128_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16314_ _08948_ _09292_ _09404_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10738_ net6910 net2244 _04182_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__mux2_1
X_13526_ _06576_ _06694_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17294_ _10199_ _10201_ _10312_ vssd1 vssd1 vccd1 vccd1 _10313_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19033_ net3402 net7698 _03078_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
X_16245_ _09150_ _09221_ _09242_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__a21o_1
X_13457_ _06564_ _06627_ _06505_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10669_ net2626 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ _05591_ _05592_ _05204_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__mux2_1
X_16176_ _09258_ _09268_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__xor2_2
X_13388_ _06406_ _06464_ _06525_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12339_ _05517_ _05522_ _05524_ _05465_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15127_ _06006_ _06331_ net4180 vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3609 _00480_ vssd1 vssd1 vccd1 vccd1 net4136 sky130_fd_sc_hd__dlygate4sd3_1
X_19935_ net3122 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
X_15058_ _06364_ _06321_ _06317_ net8410 vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__or4_1
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2908 rbzero.pov.ready_buffer\[37\] vssd1 vssd1 vccd1 vccd1 net3435 sky130_fd_sc_hd__dlygate4sd3_1
X_14009_ _07120_ _07125_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__nand2_1
Xhold2919 net5773 vssd1 vssd1 vccd1 vccd1 net3446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19866_ net2921 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18817_ net3909 net5845 _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nor3_1
X_20641__369 clknet_1_0__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__inv_2
X_18748_ _02865_ net4686 net3678 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18679_ _02832_ _02833_ rbzero.wall_tracer.rayAddendY\[1\] _09735_ vssd1 vssd1 vccd1
+ vccd1 _02834_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_204_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20710_ _03890_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21690_ clknet_leaf_28_i_clk net3994 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20572_ clknet_1_1__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__buf_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20535__274 clknet_1_0__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__inv_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6202 net1904 vssd1 vssd1 vccd1 vccd1 net6729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6213 _03371_ vssd1 vssd1 vccd1 vccd1 net6740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6224 rbzero.tex_r1\[21\] vssd1 vssd1 vccd1 vccd1 net6751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6235 net1900 vssd1 vssd1 vccd1 vccd1 net6762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5501 net624 vssd1 vssd1 vccd1 vccd1 net6028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6246 rbzero.tex_g1\[16\] vssd1 vssd1 vccd1 vccd1 net6773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6257 net1985 vssd1 vssd1 vccd1 vccd1 net6784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5512 _04020_ vssd1 vssd1 vccd1 vccd1 net6039 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_147_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6268 rbzero.tex_g1\[59\] vssd1 vssd1 vccd1 vccd1 net6795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5523 net1593 vssd1 vssd1 vccd1 vccd1 net6050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5534 net3038 vssd1 vssd1 vccd1 vccd1 net6061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6279 net1820 vssd1 vssd1 vccd1 vccd1 net6806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4800 rbzero.wall_tracer.mapX\[10\] vssd1 vssd1 vccd1 vccd1 net5327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5545 net642 vssd1 vssd1 vccd1 vccd1 net6072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5556 rbzero.tex_r0\[24\] vssd1 vssd1 vccd1 vccd1 net6083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4811 net914 vssd1 vssd1 vccd1 vccd1 net5338 sky130_fd_sc_hd__dlygate4sd3_1
X_22173_ clknet_4_7__leaf_i_clk net2615 vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5567 net804 vssd1 vssd1 vccd1 vccd1 net6094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4822 _00804_ vssd1 vssd1 vccd1 vccd1 net5349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5578 net939 vssd1 vssd1 vccd1 vccd1 net6105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4833 net953 vssd1 vssd1 vccd1 vccd1 net5360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5589 net965 vssd1 vssd1 vccd1 vccd1 net6116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4844 rbzero.spi_registers.texadd0\[13\] vssd1 vssd1 vccd1 vccd1 net5371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4855 net855 vssd1 vssd1 vccd1 vccd1 net5382 sky130_fd_sc_hd__dlygate4sd3_1
X_21124_ clknet_leaf_107_i_clk net3780 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4866 _00782_ vssd1 vssd1 vccd1 vccd1 net5393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4877 net830 vssd1 vssd1 vccd1 vccd1 net5404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4888 rbzero.mapdxw\[1\] vssd1 vssd1 vccd1 vccd1 net5415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4899 net1037 vssd1 vssd1 vccd1 vccd1 net5426 sky130_fd_sc_hd__dlygate4sd3_1
X_21055_ clknet_leaf_74_i_clk _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20006_ _03609_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21957_ net399 net2178 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ net4132 _04889_ _04898_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ clknet_leaf_81_i_clk _00395_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ net3 _05865_ _05864_ clknet_1_1__leaf__05645_ vssd1 vssd1 vccd1 vccd1 _05868_
+ sky130_fd_sc_hd__a22o_2
X_21888_ net330 net2733 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19762__43 clknet_1_1__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
X_11641_ _04796_ _04814_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__or3_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _03996_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__buf_1
XFILLER_0_193_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ _07519_ _07528_ _07530_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__a21oi_4
X_11572_ net1105 net1156 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _06392_ _06481_ _06473_ _06401_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10523_ net976 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_4
X_14291_ net8355 _07393_ _07387_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16030_ _09122_ _09123_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__nand2_1
X_13242_ _06409_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xnor2_1
Xhold7470 rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1 vccd1 net7997 sky130_fd_sc_hd__dlygate4sd3_1
X_10454_ net3068 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__clkbuf_1
Xhold7481 _08533_ vssd1 vssd1 vccd1 vccd1 net8008 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7492 _00508_ vssd1 vssd1 vccd1 vccd1 net8019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6780 _04368_ vssd1 vssd1 vccd1 vccd1 net7307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13173_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__mux2_4
Xhold6791 net2301 vssd1 vssd1 vccd1 vccd1 net7318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12124_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _04837_ vssd1 vssd1 vccd1 vccd1 _05312_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17981_ _02189_ _02216_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19720_ net7685 net5280 net7273 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__and3_1
X_16932_ _09657_ _09659_ _09658_ vssd1 vssd1 vccd1 vccd1 _09954_ sky130_fd_sc_hd__o21bai_2
X_12055_ _04967_ _05228_ _05232_ _04991_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__o311a_1
X_11006_ net7101 net3163 _04320_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
X_19651_ net6516 net1447 _03441_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
X_16863_ _09883_ _09884_ _09876_ _09878_ vssd1 vssd1 vccd1 vccd1 _09885_ sky130_fd_sc_hd__a211o_1
X_18602_ net3619 net1002 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__nor2_1
X_15814_ _08494_ _08277_ _08253_ _08464_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__and4bb_1
X_19582_ net6287 net2953 _03403_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__mux2_1
X_16794_ _09823_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__clkbuf_1
X_18533_ _04490_ _02704_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15745_ _08839_ _08837_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__xnor2_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _06039_ net3848 net4044 net3807 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__and4_1
XFILLER_0_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _02623_ _02625_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__and2_1
X_11908_ net3461 _05080_ _05090_ net3348 _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a221o_1
X_15676_ _08185_ _08204_ _08464_ _08573_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ net4048 vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17415_ _08140_ _10432_ vssd1 vssd1 vccd1 vccd1 _10433_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _07446_ _07447_ _07797_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__o21a_1
X_11839_ net4335 net4259 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__nand2_1
X_18395_ _02573_ _02578_ _04480_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17346_ _10360_ _10363_ vssd1 vssd1 vccd1 vccd1 _10365_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ _07704_ _07728_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _06676_ _06677_ _06679_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__a21bo_1
X_17277_ _08661_ _09116_ vssd1 vssd1 vccd1 vccd1 _10296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ _07657_ _07659_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20666__12 clknet_1_0__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XFILLER_0_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19016_ net3900 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
X_16228_ _09217_ _09320_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__nand2_2
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4107 _09844_ vssd1 vssd1 vccd1 vccd1 net4634 sky130_fd_sc_hd__dlygate4sd3_1
X_16159_ _08996_ _09249_ _08864_ _09135_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__a22o_1
Xhold4118 _06115_ vssd1 vssd1 vccd1 vccd1 net4645 sky130_fd_sc_hd__buf_1
Xhold4129 net7975 vssd1 vssd1 vccd1 vccd1 net4656 sky130_fd_sc_hd__dlygate4sd3_1
X_20681__26 clknet_1_0__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3406 net8357 vssd1 vssd1 vccd1 vccd1 net3933 sky130_fd_sc_hd__buf_1
Xhold3417 net4872 vssd1 vssd1 vccd1 vccd1 net3944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3428 _04597_ vssd1 vssd1 vccd1 vccd1 net3955 sky130_fd_sc_hd__clkbuf_2
Xhold3439 net5919 vssd1 vssd1 vccd1 vccd1 net3966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2705 _01088_ vssd1 vssd1 vccd1 vccd1 net3232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2716 net7529 vssd1 vssd1 vccd1 vccd1 net3243 sky130_fd_sc_hd__dlygate4sd3_1
X_19918_ net3135 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
Xhold2727 _00693_ vssd1 vssd1 vccd1 vccd1 net3254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 _01369_ vssd1 vssd1 vccd1 vccd1 net3265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2749 net7549 vssd1 vssd1 vccd1 vccd1 net3276 sky130_fd_sc_hd__buf_1
X_19849_ net1183 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21811_ net253 net2109 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21742_ clknet_leaf_100_i_clk net5478 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21673_ clknet_leaf_124_i_clk net1868 vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6010 rbzero.tex_b0\[34\] vssd1 vssd1 vccd1 vccd1 net6537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6021 net1526 vssd1 vssd1 vccd1 vccd1 net6548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6032 rbzero.pov.ready_buffer\[4\] vssd1 vssd1 vccd1 vccd1 net6559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6043 net1685 vssd1 vssd1 vccd1 vccd1 net6570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6054 net1605 vssd1 vssd1 vccd1 vccd1 net6581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6065 rbzero.tex_g0\[57\] vssd1 vssd1 vccd1 vccd1 net6592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5320 net2200 vssd1 vssd1 vccd1 vccd1 net5847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6076 net1718 vssd1 vssd1 vccd1 vccd1 net6603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5331 rbzero.debug_overlay.playerY\[-7\] vssd1 vssd1 vccd1 vccd1 net5858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6087 rbzero.tex_g1\[55\] vssd1 vssd1 vccd1 vccd1 net6614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5342 _03637_ vssd1 vssd1 vccd1 vccd1 net5869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5353 _00642_ vssd1 vssd1 vccd1 vccd1 net5880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6098 net1698 vssd1 vssd1 vccd1 vccd1 net6625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5364 _02665_ vssd1 vssd1 vccd1 vccd1 net5891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5375 _06757_ vssd1 vssd1 vccd1 vccd1 net5902 sky130_fd_sc_hd__clkbuf_4
Xhold4630 net740 vssd1 vssd1 vccd1 vccd1 net5157 sky130_fd_sc_hd__dlygate4sd3_1
X_22156_ clknet_leaf_55_i_clk _01643_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4641 rbzero.spi_registers.texadd1\[13\] vssd1 vssd1 vccd1 vccd1 net5168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5386 _05069_ vssd1 vssd1 vccd1 vccd1 net5913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5397 rbzero.wall_tracer.rayAddendY\[-4\] vssd1 vssd1 vccd1 vccd1 net5924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4652 net784 vssd1 vssd1 vccd1 vccd1 net5179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4663 _00873_ vssd1 vssd1 vccd1 vccd1 net5190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4674 net844 vssd1 vssd1 vccd1 vccd1 net5201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3940 net8177 vssd1 vssd1 vccd1 vccd1 net4467 sky130_fd_sc_hd__dlygate4sd3_1
X_21107_ clknet_leaf_20_i_clk net1601 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4685 net824 vssd1 vssd1 vccd1 vccd1 net5212 sky130_fd_sc_hd__dlygate4sd3_1
X_22087_ net149 net2261 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
Xhold3951 _01198_ vssd1 vssd1 vccd1 vccd1 net4478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4696 rbzero.spi_registers.texadd3\[15\] vssd1 vssd1 vccd1 vccd1 net5223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3962 net1056 vssd1 vssd1 vccd1 vccd1 net4489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3973 net3655 vssd1 vssd1 vccd1 vccd1 net4500 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3984 rbzero.row_render.size\[6\] vssd1 vssd1 vccd1 vccd1 net4511 sky130_fd_sc_hd__dlygate4sd3_1
X_21038_ clknet_leaf_31_i_clk net5474 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3995 net3726 vssd1 vssd1 vccd1 vccd1 net4522 sky130_fd_sc_hd__buf_1
XFILLER_0_22_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _07025_ _07024_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12811_ _05980_ _05982_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13791_ _06933_ _06930_ _06932_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15530_ _08595_ _08603_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__xnor2_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12742_ net37 _05905_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__or3b_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _08522_ _08523_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ net28 vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__03507_ clknet_0__03507_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03507_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _10219_ vssd1 vssd1 vccd1 vccd1 _10220_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11624_ net4450 _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__nor2_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _07580_ _07582_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__nor2_1
X_18180_ _02396_ _02398_ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a211o_1
X_15392_ _08479_ _08482_ _08481_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17131_ _10150_ vssd1 vssd1 vccd1 vccd1 _10151_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14343_ _07306_ _07280_ _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__or3b_4
X_11555_ net4354 _04464_ _04501_ net4431 vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ net5600 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__clkbuf_1
X_17062_ _09958_ _09960_ _09957_ vssd1 vssd1 vccd1 vccd1 _10083_ sky130_fd_sc_hd__a21bo_1
X_14274_ _07443_ _07444_ _07339_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ net4138 _04674_ net3443 _04464_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16013_ net4559 _08115_ _09106_ _09107_ _01633_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__o221a_1
X_13225_ _06306_ _06370_ _06380_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ _06324_ _06326_ _06306_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__mux2_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _02115_ _02116_ _02118_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a21bo_1
X_13087_ net2058 _06244_ _06258_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__a21oi_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19703_ net6564 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__clkbuf_1
X_16915_ _09934_ _09936_ vssd1 vssd1 vccd1 vccd1 _09937_ sky130_fd_sc_hd__nand2_1
X_12038_ _05206_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or2_1
X_17895_ _02097_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19634_ net1469 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__clkbuf_1
X_16846_ _09867_ _09868_ net3799 vssd1 vssd1 vccd1 vccd1 _09870_ sky130_fd_sc_hd__a21oi_1
X_19565_ net1430 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
X_16777_ _09804_ _09807_ vssd1 vssd1 vccd1 vccd1 _09808_ sky130_fd_sc_hd__xnor2_1
X_13989_ _07159_ _06793_ _06757_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ _02676_ _02686_ _02690_ _04480_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a31o_1
X_15728_ _08819_ _08820_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19496_ net1879 _02472_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18447_ _02626_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__clkbuf_4
X_15659_ _08708_ _08753_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18378_ _02554_ _02560_ net4784 net8047 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ _08948_ _08916_ _09970_ vssd1 vssd1 vccd1 vccd1 _10348_ sky130_fd_sc_hd__or3_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20271_ net4071 net4098 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22010_ net452 net2142 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3203 _02330_ vssd1 vssd1 vccd1 vccd1 net3730 sky130_fd_sc_hd__dlygate4sd3_1
X_20647__375 clknet_1_1__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__inv_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3236 net4859 vssd1 vssd1 vccd1 vccd1 net3763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2502 net7472 vssd1 vssd1 vccd1 vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3247 _04484_ vssd1 vssd1 vccd1 vccd1 net3774 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2513 _00704_ vssd1 vssd1 vccd1 vccd1 net3040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3258 net3428 vssd1 vssd1 vccd1 vccd1 net3785 sky130_fd_sc_hd__clkbuf_2
X_20346__103 clknet_1_1__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__inv_2
Xhold2524 rbzero.pov.spi_buffer\[52\] vssd1 vssd1 vccd1 vccd1 net3051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3269 net7996 vssd1 vssd1 vccd1 vccd1 net3796 sky130_fd_sc_hd__buf_1
Xhold2535 _01145_ vssd1 vssd1 vccd1 vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1801 net7068 vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2546 net3255 vssd1 vssd1 vccd1 vccd1 net3073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1812 net6978 vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2557 _02949_ vssd1 vssd1 vccd1 vccd1 net3084 sky130_fd_sc_hd__clkbuf_2
Xhold1823 _01592_ vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 net3124 vssd1 vssd1 vccd1 vccd1 net3095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _04391_ vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 _01407_ vssd1 vssd1 vccd1 vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1845 _01542_ vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1856 _01059_ vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 _04032_ vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 net6917 vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 _01011_ vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21725_ clknet_leaf_110_i_clk net3883 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21656_ clknet_leaf_121_i_clk net3285 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20392__145 clknet_1_0__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__inv_2
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21587_ net221 net2169 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11340_ rbzero.texu_hot\[3\] _04518_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or2_1
X_20538_ clknet_1_0__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__buf_1
Xtop_ew_algofoogle_97 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_97/HI o_rgb[4] sky130_fd_sc_hd__conb_1
XFILLER_0_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ net5205 vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5150 net5598 vssd1 vssd1 vccd1 vccd1 net5677 sky130_fd_sc_hd__dlygate4sd3_1
X_13010_ net3749 _06174_ _06184_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__a211o_1
Xhold5161 net1124 vssd1 vssd1 vccd1 vccd1 net5688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5172 rbzero.tex_g1\[2\] vssd1 vssd1 vccd1 vccd1 net5699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5183 net2193 vssd1 vssd1 vccd1 vccd1 net5710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5194 rbzero.wall_tracer.mapX\[9\] vssd1 vssd1 vccd1 vccd1 net5721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4460 rbzero.spi_registers.texadd3\[20\] vssd1 vssd1 vccd1 vccd1 net4987 sky130_fd_sc_hd__dlygate4sd3_1
X_22139_ clknet_leaf_37_i_clk _01626_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold4471 _01014_ vssd1 vssd1 vccd1 vccd1 net4998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4482 net727 vssd1 vssd1 vccd1 vccd1 net5009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4493 rbzero.spi_registers.texadd3\[10\] vssd1 vssd1 vccd1 vccd1 net5020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3770 net7921 vssd1 vssd1 vccd1 vccd1 net4297 sky130_fd_sc_hd__dlygate4sd3_1
X_14961_ net4471 _07968_ _08068_ vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__mux2_1
Xhold3781 net1078 vssd1 vssd1 vccd1 vccd1 net4308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3792 net7925 vssd1 vssd1 vccd1 vccd1 net4319 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ net1038 _09745_ _09746_ net8009 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_3__f_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13912_ _07058_ _07060_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17680_ _08918_ _10211_ _09970_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__or3_1
XFILLER_0_199_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14892_ rbzero.wall_tracer.visualWallDist\[-10\] _08037_ _08038_ vssd1 vssd1 vccd1
+ vccd1 _08040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16631_ net4123 vssd1 vssd1 vccd1 vccd1 _09720_ sky130_fd_sc_hd__clkbuf_2
X_13843_ _06999_ _07001_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19350_ net4992 _03269_ _03276_ _03275_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__o211a_1
X_16562_ _09650_ _09651_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__nand2_1
X_10986_ net6876 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
X_13774_ _06943_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18301_ net6380 net3592 _02493_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
X_15513_ _08606_ _08607_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__and2b_2
XFILLER_0_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19281_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__buf_2
X_12725_ net35 _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nor2_2
X_16493_ _09581_ _09583_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__nor2_1
X_18232_ _02448_ net3820 _02393_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
X_15444_ _08537_ _08538_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ net25 net24 net26 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_111_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11607_ _04780_ _04777_ _04779_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__and3_1
X_18163_ net3790 net3777 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15375_ _08420_ _08469_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__xnor2_2
X_12587_ net4066 _05744_ _05763_ net71 _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a221o_1
X_17114_ _10134_ net4589 net4649 vssd1 vssd1 vccd1 vccd1 _10135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03852_ _03852_ vssd1 vssd1 vccd1 vccd1 clknet_0__03852_ sky130_fd_sc_hd__clkbuf_16
X_14326_ _07486_ _07495_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18094_ _02327_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__clkbuf_1
X_11538_ net4384 vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 _01553_ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17045_ _09915_ _08616_ _10064_ vssd1 vssd1 vccd1 vccd1 _10066_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold419 net5367 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ _07410_ _07426_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__a21oi_1
X_11469_ _04657_ _04658_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_126_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13208_ net8261 _06266_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _07357_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__or2b_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _06264_ _06309_ _06307_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a21oi_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ net3009 net5826 _03058_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _03369_ vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ _02164_ _02183_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__xnor2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1119 net3297 vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17878_ _09040_ _08612_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19617_ net6255 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
X_16829_ _09818_ _09326_ vssd1 vssd1 vccd1 vccd1 _09855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19548_ net6544 net4016 _03388_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _03352_ net3903 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21510_ clknet_leaf_48_i_clk net1802 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21441_ clknet_leaf_26_i_clk net1428 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21372_ clknet_leaf_44_i_clk net5115 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20323_ net6683 net1447 _03825_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold920 net7584 vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold931 _00584_ vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold942 _03442_ vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 net6018 vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
X_20254_ net4103 net4122 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__nand2_1
Xhold964 _01000_ vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3000 net5808 vssd1 vssd1 vccd1 vccd1 net3527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 net6469 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3011 net4527 vssd1 vssd1 vccd1 vccd1 net3538 sky130_fd_sc_hd__clkbuf_2
Xhold986 _00999_ vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3022 _03328_ vssd1 vssd1 vccd1 vccd1 net3549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3033 net4672 vssd1 vssd1 vccd1 vccd1 net3560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 net6208 vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
X_20185_ _03728_ net3566 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3044 _03314_ vssd1 vssd1 vccd1 vccd1 net3571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2310 _01023_ vssd1 vssd1 vccd1 vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3055 _01211_ vssd1 vssd1 vccd1 vccd1 net3582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 rbzero.tex_g1\[11\] vssd1 vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3066 _03096_ vssd1 vssd1 vccd1 vccd1 net3593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 _01344_ vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3077 rbzero.wall_tracer.rayAddendX\[2\] vssd1 vssd1 vccd1 vccd1 net3604 sky130_fd_sc_hd__buf_2
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2343 _03531_ vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3088 _02680_ vssd1 vssd1 vccd1 vccd1 net3615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03841_ clknet_0__03841_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03841_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2354 _04088_ vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3099 net8447 vssd1 vssd1 vccd1 vccd1 net3626 sky130_fd_sc_hd__buf_1
Xhold2365 net7319 vssd1 vssd1 vccd1 vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 net6740 vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 net6905 vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2376 net7454 vssd1 vssd1 vccd1 vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1642 _01074_ vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2387 net7414 vssd1 vssd1 vccd1 vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2398 _01396_ vssd1 vssd1 vccd1 vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1653 _03544_ vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1664 net7176 vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1675 _04113_ vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1686 _01058_ vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1697 net6961 vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10840_ net2966 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ net2433 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20400__152 clknet_1_1__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__inv_2
XFILLER_0_17_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ net10 vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13490_ _06660_ _06552_ _06547_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__mux2_1
X_21708_ clknet_leaf_119_i_clk net3555 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ _04706_ _04751_ _05541_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__or3_1
X_21639_ clknet_leaf_127_i_clk net3322 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ rbzero.tex_b1\[31\] rbzero.tex_b1\[30\] _05250_ vssd1 vssd1 vccd1 vccd1 _05557_
+ sky130_fd_sc_hd__mux2_1
X_15160_ _08253_ _08254_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__nand2_2
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_i_clk clknet_4_8__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14111_ _07242_ _07233_ _07281_ _07033_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__o22a_1
X_11323_ rbzero.texu_hot\[5\] _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nand2_1
X_15091_ net3637 _08181_ _08185_ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ net7115 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__clkbuf_1
X_14042_ _06729_ _06923_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18850_ net3695 net5800 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_58_i_clk clknet_4_15__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11185_ net7061 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17801_ _02000_ _02039_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__xnor2_2
Xhold4290 _00965_ vssd1 vssd1 vccd1 vccd1 net4817 sky130_fd_sc_hd__dlygate4sd3_1
X_18781_ _02914_ _02924_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15993_ _09086_ _09087_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__nand2_1
X_17732_ _10408_ _09345_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__nor2_1
X_14944_ _08069_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _08799_ _10096_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__nor2_1
X_14875_ net7811 _07995_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19402_ net2256 _03303_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__or2_1
X_16614_ _09596_ _09703_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13826_ _06992_ _06996_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__or2_4
X_17594_ _01743_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19333_ net1599 _03237_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__or2_1
X_16545_ _09532_ _09523_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__or2b_1
XFILLER_0_175_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13757_ _06889_ _06887_ _06888_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__nand3_1
X_10969_ net6199 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19264_ net5284 _03216_ _03225_ _03219_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__o211a_1
X_12708_ net46 _05865_ _05853_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a21bo_1
X_16476_ _09565_ _09566_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__nor2_1
X_13688_ _06857_ _06858_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18215_ _02433_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__clkbuf_1
X_15427_ _08229_ _08294_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19195_ net5292 _03182_ _03185_ _03176_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__o211a_1
X_12639_ net22 net23 vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__and2b_1
XFILLER_0_182_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6609 rbzero.tex_g1\[43\] vssd1 vssd1 vccd1 vccd1 net7136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ net3785 net4390 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _08434_ _08452_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__xor2_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5908 rbzero.pov.spi_buffer\[33\] vssd1 vssd1 vccd1 vccd1 net6435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14309_ _07463_ _07478_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__and2_1
Xhold5919 net1474 vssd1 vssd1 vccd1 vccd1 net6446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 net5122 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
X_18077_ _02254_ _02309_ _02310_ _02312_ net90 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a311o_1
X_15289_ net4471 _06121_ _08383_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__a21boi_4
Xhold216 net5102 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 net8231 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold238 net5150 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _10039_ _10048_ vssd1 vssd1 vccd1 vccd1 _10049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold249 net4448 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ net2873 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__clkbuf_4
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21990_ net432 net2663 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
X_20941_ clknet_leaf_77_i_clk net4760 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20872_ _02509_ _02518_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__and2b_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20458__204 clknet_1_0__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__inv_2
XFILLER_0_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7800 net4484 vssd1 vssd1 vccd1 vccd1 net8327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7811 rbzero.wall_tracer.stepDistX\[6\] vssd1 vssd1 vccd1 vccd1 net8338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7822 net4460 vssd1 vssd1 vccd1 vccd1 net8349 sky130_fd_sc_hd__dlygate4sd3_1
X_21424_ clknet_leaf_36_i_clk net1482 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7855 net4396 vssd1 vssd1 vccd1 vccd1 net8382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7866 _08222_ vssd1 vssd1 vccd1 vccd1 net8393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7877 rbzero.wall_tracer.stepDistX\[5\] vssd1 vssd1 vccd1 vccd1 net8404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7888 rbzero.wall_tracer.stepDistX\[-6\] vssd1 vssd1 vccd1 vccd1 net8415 sky130_fd_sc_hd__dlygate4sd3_1
X_21355_ clknet_leaf_10_i_clk net5087 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20306_ net1475 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold750 _01534_ vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21286_ clknet_leaf_27_i_clk net5616 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold761 _00572_ vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _04321_ vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
X_20237_ net2310 net7273 _03492_ net3950 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a31o_1
Xhold783 net6312 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _00947_ vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20168_ net7552 _03707_ net4467 _03732_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__o211a_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 net7450 vssd1 vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2151 _01519_ vssd1 vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2162 _04045_ vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
X_19769__49 clknet_1_1__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_0_196_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2173 net6909 vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _06164_ net3787 _06165_ net3932 vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__a22o_1
X_20099_ net4052 _03682_ net4436 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__o21ai_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2184 net4316 vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2195 net7231 vssd1 vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1450 net6837 vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1461 net2238 vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ net3433 _05095_ _05128_ _05129_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a211o_1
Xhold1472 _00946_ vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1483 _01454_ vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 _04083_ vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14660_ _07814_ _07827_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__nand2_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ net4115 _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and2b_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13611_ _06575_ _06702_ _06692_ _06754_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ net6774 net7340 _04227_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
X_14591_ _07750_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__nand2_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16330_ _09412_ _09421_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__xnor2_1
X_13542_ _06709_ _06710_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__nand2_1
X_10754_ net6203 net6772 _04182_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _08542_ _09062_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10685_ net7208 net6979 _04149_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__mux2_1
X_13473_ _06343_ _06459_ _06639_ _06498_ _06549_ _06492_ vssd1 vssd1 vccd1 vccd1 _06644_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18000_ _02150_ _02153_ _02148_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a21bo_1
X_15212_ _08255_ _08280_ _08294_ _08306_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__or4_1
X_12424_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _04951_ vssd1 vssd1 vccd1 vccd1 _05609_
+ sky130_fd_sc_hd__mux2_1
X_16192_ _09283_ _09284_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ _08236_ _08237_ vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__nand2_1
X_12355_ _05189_ _05198_ _05456_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ _04494_ _04496_ _04021_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__o21ai_1
X_12286_ _05276_ _05469_ _05471_ _04928_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19951_ net7449 net3159 _03583_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__mux2_1
X_15074_ net3348 net3536 net4168 vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11237_ net7281 net2892 _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__mux2_1
X_14025_ _07142_ _07147_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__or2_1
X_18902_ net7443 net3182 _03014_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19882_ net3342 net3302 _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__mux2_1
X_11168_ net6790 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__clkbuf_1
X_18833_ net5878 net1547 _02968_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or3b_1
XFILLER_0_208_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18764_ _02911_ _02912_ _02895_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15976_ _09057_ _09058_ _09069_ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__and3_1
X_11099_ net5588 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20407__158 clknet_1_0__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__inv_2
XFILLER_0_136_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17715_ _01954_ net3875 _10260_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14927_ net4659 _08050_ _08052_ net3803 net4752 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__o221a_1
X_18695_ _02846_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nand2_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17646_ _01884_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _07913_ _07985_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ _06976_ _06978_ _06979_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__a21oi_1
X_17577_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14789_ net7846 _07935_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19316_ net1380 _03251_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__or2_1
X_16528_ _09373_ _09254_ _09351_ _09249_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7107 rbzero.debug_overlay.playerY\[3\] vssd1 vssd1 vccd1 vccd1 net7634 sky130_fd_sc_hd__dlygate4sd3_1
X_19247_ net5061 _03201_ _03215_ _03206_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__o211a_1
X_16459_ _09547_ _09549_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__xnor2_2
Xhold7118 _03741_ vssd1 vssd1 vccd1 vccd1 net7645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7129 _03502_ vssd1 vssd1 vccd1 vccd1 net7656 sky130_fd_sc_hd__buf_1
Xhold6406 _04449_ vssd1 vssd1 vccd1 vccd1 net6933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6417 net1774 vssd1 vssd1 vccd1 vccd1 net6944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19178_ _09721_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__buf_4
XFILLER_0_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6428 rbzero.tex_b1\[5\] vssd1 vssd1 vccd1 vccd1 net6955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6439 rbzero.tex_r1\[5\] vssd1 vssd1 vccd1 vccd1 net6966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5705 _03008_ vssd1 vssd1 vccd1 vccd1 net6232 sky130_fd_sc_hd__dlygate4sd3_1
X_18129_ net3757 net4379 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__nor2_1
Xhold5716 net1191 vssd1 vssd1 vccd1 vccd1 net6243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5727 _03433_ vssd1 vssd1 vccd1 vccd1 net6254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5738 net1214 vssd1 vssd1 vccd1 vccd1 net6265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5749 rbzero.tex_r0\[29\] vssd1 vssd1 vccd1 vccd1 net6276 sky130_fd_sc_hd__dlygate4sd3_1
X_21140_ clknet_leaf_95_i_clk net3525 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21071_ clknet_leaf_78_i_clk _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20022_ _08297_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21973_ net415 net1488 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer20 net546 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer31 net3463 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer42 _06913_ vssd1 vssd1 vccd1 vccd1 net3513 sky130_fd_sc_hd__clkbuf_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer53 net579 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_1
X_20924_ clknet_leaf_69_i_clk _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20855_ net4213 _04001_ _04002_ _09326_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a22o_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20786_ _03949_ _03952_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7630 rbzero.map_overlay.i_otherx\[4\] vssd1 vssd1 vccd1 vccd1 net8157 sky130_fd_sc_hd__dlygate4sd3_1
X_10470_ net6691 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7641 rbzero.map_overlay.i_mapdy\[3\] vssd1 vssd1 vccd1 vccd1 net8168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7652 _03714_ vssd1 vssd1 vccd1 vccd1 net8179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7663 _08039_ vssd1 vssd1 vccd1 vccd1 net8190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7685 _03722_ vssd1 vssd1 vccd1 vccd1 net8212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6940 net2830 vssd1 vssd1 vccd1 vccd1 net7467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21407_ clknet_leaf_35_i_clk net4954 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6951 _04266_ vssd1 vssd1 vccd1 vccd1 net7478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7696 rbzero.traced_texa\[3\] vssd1 vssd1 vccd1 vccd1 net8223 sky130_fd_sc_hd__dlygate4sd3_1
X_20512__253 clknet_1_0__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__inv_2
Xhold6962 rbzero.pov.ready_buffer\[8\] vssd1 vssd1 vccd1 vccd1 net7489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6973 net3202 vssd1 vssd1 vccd1 vccd1 net7500 sky130_fd_sc_hd__dlygate4sd3_1
X_12140_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _04836_ vssd1 vssd1 vccd1 vccd1 _05328_
+ sky130_fd_sc_hd__mux2_1
Xhold6984 _03072_ vssd1 vssd1 vccd1 vccd1 net7511 sky130_fd_sc_hd__dlygate4sd3_1
X_21338_ clknet_leaf_6_i_clk net5310 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6995 net1830 vssd1 vssd1 vccd1 vccd1 net7522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ rbzero.tex_r1\[43\] rbzero.tex_r1\[42\] _04923_ vssd1 vssd1 vccd1 vccd1 _05260_
+ sky130_fd_sc_hd__mux2_1
X_21269_ clknet_leaf_25_i_clk net5757 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold580 net4281 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 net5455 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net6896 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15830_ _08914_ _08923_ _08924_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__a21oi_2
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _08854_ _08855_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__nor2_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ net4152 _06104_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__xor2_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _10425_ _01739_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a21oi_2
Xhold1280 _01398_ vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 net5528 vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ net8442 _07850_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__nor2_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _02626_ net4698 _02656_ _02657_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a2bb2o_1
X_11924_ _04501_ _05088_ _05092_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nor3_4
X_15692_ _08782_ _08785_ _08786_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__o21ai_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17431_ _01670_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__xor2_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14643_ _07812_ _07813_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__and2_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11855_ _05043_ net4127 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__nand2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ net2996 net6643 _04216_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
X_17362_ _09809_ _10264_ _10265_ _10380_ vssd1 vssd1 vccd1 vccd1 _10381_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_32_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14574_ _07489_ _07327_ _07742_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__or3_1
X_11786_ _04846_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19101_ net3333 _03126_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or2_1
X_16313_ _08948_ _09403_ _09404_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__nor3_1
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _06695_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__clkbuf_4
X_17293_ _10192_ _10202_ vssd1 vssd1 vccd1 vccd1 _10312_ sky130_fd_sc_hd__or2b_1
XFILLER_0_166_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10737_ net6229 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19032_ net3817 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__clkbuf_1
X_16244_ _09318_ _09319_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__or2_2
XFILLER_0_67_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _06492_ _06625_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10668_ net7222 net6703 _04138_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12407_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _05250_ vssd1 vssd1 vccd1 vccd1 _05592_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _09266_ _09267_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__nor2_1
X_10599_ net6983 net6906 _04105_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__mux2_1
X_13387_ _06528_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__buf_2
XFILLER_0_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ _08220_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__buf_2
X_12338_ _05276_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__or2_1
X_20487__230 clknet_1_1__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__inv_2
XFILLER_0_121_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19934_ net3121 net7560 _03572_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__mux2_1
X_15057_ _06334_ _06331_ _06324_ net8409 vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__or4_1
X_12269_ _04736_ _05176_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2909 net7659 vssd1 vssd1 vccd1 vccd1 net3436 sky130_fd_sc_hd__dlygate4sd3_1
X_14008_ _07177_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__nand2_1
X_19865_ net3056 net7443 _03539_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18816_ _02955_ _02951_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15959_ _09051_ _09053_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__nor2_1
X_18747_ _02865_ net4686 _02895_ _02896_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18678_ _02830_ _02831_ _04481_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17629_ _01867_ _01868_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6203 rbzero.pov.spi_buffer\[37\] vssd1 vssd1 vccd1 vccd1 net6730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6214 rbzero.spi_registers.new_mapd\[13\] vssd1 vssd1 vccd1 vccd1 net6741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6225 net1912 vssd1 vssd1 vccd1 vccd1 net6752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6236 rbzero.tex_b1\[45\] vssd1 vssd1 vccd1 vccd1 net6763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5502 rbzero.tex_b0\[20\] vssd1 vssd1 vccd1 vccd1 net6029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6247 net2085 vssd1 vssd1 vccd1 vccd1 net6774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6258 _04218_ vssd1 vssd1 vccd1 vccd1 net6785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5513 gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5524 rbzero.tex_b1\[6\] vssd1 vssd1 vccd1 vccd1 net6051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6269 net1994 vssd1 vssd1 vccd1 vccd1 net6796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5535 _03702_ vssd1 vssd1 vccd1 vccd1 net6062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5546 _04283_ vssd1 vssd1 vccd1 vccd1 net6073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4801 net832 vssd1 vssd1 vccd1 vccd1 net5328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22172_ clknet_leaf_67_i_clk net4930 vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5557 net766 vssd1 vssd1 vccd1 vccd1 net6084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4812 rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 net5339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4823 net956 vssd1 vssd1 vccd1 vccd1 net5350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5568 rbzero.tex_b0\[30\] vssd1 vssd1 vccd1 vccd1 net6095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5579 rbzero.tex_g0\[22\] vssd1 vssd1 vccd1 vccd1 net6106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4834 _00860_ vssd1 vssd1 vccd1 vccd1 net5361 sky130_fd_sc_hd__dlygate4sd3_1
X_21123_ clknet_leaf_92_i_clk net4830 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4845 net980 vssd1 vssd1 vccd1 vccd1 net5372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4856 rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 net5383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4867 net952 vssd1 vssd1 vccd1 vccd1 net5394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4878 _01605_ vssd1 vssd1 vccd1 vccd1 net5405 sky130_fd_sc_hd__dlygate4sd3_1
X_21054_ clknet_leaf_74_i_clk _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4889 net1004 vssd1 vssd1 vccd1 vccd1 net5416 sky130_fd_sc_hd__dlygate4sd3_1
X_20005_ net3269 _08198_ _03615_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21956_ net398 net966 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ clknet_leaf_81_i_clk _00394_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ net329 net2618 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__and2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20838_ _03320_ clknet_1_1__leaf__05742_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__and2_2
X_11571_ net1105 net1156 vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nand2_1
X_20769_ _03878_ _03940_ _03941_ _03883_ net5492 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _06378_ _06393_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10522_ net5696 net2797 _04064_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__mux2_1
X_14290_ _07459_ _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__nand2_2
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7460 rbzero.wall_tracer.trackDistX\[-6\] vssd1 vssd1 vccd1 vccd1 net7987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10453_ net7121 net3067 _04031_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__mux2_1
X_13241_ _06411_ _06388_ _06404_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o21a_1
Xhold7471 net3925 vssd1 vssd1 vccd1 vccd1 net7998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7482 net4757 vssd1 vssd1 vccd1 vccd1 net8009 sky130_fd_sc_hd__buf_2
XFILLER_0_161_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7493 net4240 vssd1 vssd1 vccd1 vccd1 net8020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6770 net2479 vssd1 vssd1 vccd1 vccd1 net7297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6781 net2695 vssd1 vssd1 vccd1 vccd1 net7308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13172_ rbzero.wall_tracer.rayAddendX\[-3\] _06342_ _06305_ vssd1 vssd1 vccd1 vccd1
+ _06343_ sky130_fd_sc_hd__mux2_4
XFILLER_0_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6792 rbzero.tex_b0\[11\] vssd1 vssd1 vccd1 vccd1 net7319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _04838_ vssd1 vssd1 vccd1 vccd1 _05311_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17980_ _02189_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__and2_1
X_16931_ _09931_ _09952_ vssd1 vssd1 vccd1 vccd1 _09953_ sky130_fd_sc_hd__xnor2_1
X_12054_ _05233_ _05236_ _05242_ _04825_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a211o_1
XFILLER_0_202_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11005_ net2867 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
X_16862_ net4669 net4373 vssd1 vssd1 vccd1 vccd1 _09884_ sky130_fd_sc_hd__nand2_1
X_19650_ net6729 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15813_ _08253_ _08573_ _08907_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__a21o_1
X_18601_ net3618 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19581_ net2004 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
X_16793_ _09821_ net4569 net4649 vssd1 vssd1 vccd1 vccd1 _09823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18532_ _02705_ _02691_ _04480_ _02627_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15744_ _08204_ _08573_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__nand2_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12956_ _06126_ _06128_ net4008 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ net8084 _02641_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__and2_1
X_11907_ net3443 _05093_ _05095_ net3457 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a22o_1
X_15675_ _08204_ _08464_ _08573_ _08185_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__a22o_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12887_ net3326 _06061_ _06062_ net3389 vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17414_ _08427_ _08428_ vssd1 vssd1 vccd1 vccd1 _10432_ sky130_fd_sc_hd__nand2_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14626_ _07448_ _07436_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__or2b_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11838_ net4335 net4259 _04824_ _05027_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__or4_1
X_18394_ _02574_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20519__259 clknet_1_0__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__inv_2
X_17345_ _10360_ _10363_ vssd1 vssd1 vccd1 vccd1 _10364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _07726_ _07727_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__nand2_1
X_11769_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _04950_ vssd1 vssd1 vccd1 vccd1 _04959_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _06493_ _06565_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__o21ai_1
X_17276_ _10293_ _10294_ vssd1 vssd1 vccd1 vccd1 _10295_ sky130_fd_sc_hd__and2b_1
X_14488_ _07308_ _07326_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19015_ net3793 net3899 _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
X_16227_ _09318_ _09319_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__xor2_1
X_13439_ _06394_ _06558_ _06609_ _06550_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _08864_ _09250_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4108 net8262 vssd1 vssd1 vccd1 vccd1 net4635 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4119 _06116_ vssd1 vssd1 vccd1 vccd1 net4646 sky130_fd_sc_hd__dlygate4sd3_1
X_15109_ _08118_ _08202_ _08203_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__a21o_4
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3407 net7815 vssd1 vssd1 vccd1 vccd1 net3934 sky130_fd_sc_hd__buf_1
X_16089_ _08450_ _08464_ _09182_ _09038_ _09032_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__a32o_1
Xhold3418 net3559 vssd1 vssd1 vccd1 vccd1 net3945 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3429 _09724_ vssd1 vssd1 vccd1 vccd1 net3956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2706 net7515 vssd1 vssd1 vccd1 vccd1 net3233 sky130_fd_sc_hd__dlygate4sd3_1
X_19917_ net7453 net6744 _03561_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__mux2_1
Xhold2717 _04367_ vssd1 vssd1 vccd1 vccd1 net3244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2728 rbzero.pov.spi_buffer\[32\] vssd1 vssd1 vccd1 vccd1 net3255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2739 net5848 vssd1 vssd1 vccd1 vccd1 net3266 sky130_fd_sc_hd__dlygate4sd3_1
X_19848_ net6231 net6247 _03528_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21810_ net252 net3245 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21741_ clknet_leaf_100_i_clk net4606 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21672_ clknet_leaf_123_i_clk net1871 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6000 rbzero.spi_registers.new_texadd\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net6527
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6011 net1712 vssd1 vssd1 vccd1 vccd1 net6538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6022 _04327_ vssd1 vssd1 vccd1 vccd1 net6549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6033 net1573 vssd1 vssd1 vccd1 vccd1 net6560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6044 _03831_ vssd1 vssd1 vccd1 vccd1 net6571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6055 _04036_ vssd1 vssd1 vccd1 vccd1 net6582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5310 _03619_ vssd1 vssd1 vccd1 vccd1 net5837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5321 rbzero.pov.ready_buffer\[65\] vssd1 vssd1 vccd1 vccd1 net5848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6066 net1805 vssd1 vssd1 vccd1 vccd1 net6593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6077 _02501_ vssd1 vssd1 vccd1 vccd1 net6604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5332 net3315 vssd1 vssd1 vccd1 vccd1 net5859 sky130_fd_sc_hd__clkbuf_2
Xhold6088 net1486 vssd1 vssd1 vccd1 vccd1 net6615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5343 _01176_ vssd1 vssd1 vccd1 vccd1 net5870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5354 net1549 vssd1 vssd1 vccd1 vccd1 net5881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6099 gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5365 net3891 vssd1 vssd1 vccd1 vccd1 net5892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4620 net772 vssd1 vssd1 vccd1 vccd1 net5147 sky130_fd_sc_hd__dlygate4sd3_1
X_22155_ clknet_leaf_55_i_clk _01642_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5376 rbzero.debug_overlay.playerX\[-5\] vssd1 vssd1 vccd1 vccd1 net5903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4631 _00779_ vssd1 vssd1 vccd1 vccd1 net5158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4642 net812 vssd1 vssd1 vccd1 vccd1 net5169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5387 rbzero.debug_overlay.playerX\[2\] vssd1 vssd1 vccd1 vccd1 net5914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5398 net3308 vssd1 vssd1 vccd1 vccd1 net5925 sky130_fd_sc_hd__buf_1
Xhold4653 rbzero.spi_registers.texadd2\[16\] vssd1 vssd1 vccd1 vccd1 net5180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4664 net883 vssd1 vssd1 vccd1 vccd1 net5191 sky130_fd_sc_hd__dlygate4sd3_1
X_21106_ clknet_leaf_20_i_clk net1507 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3930 net3390 vssd1 vssd1 vccd1 vccd1 net4457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4675 _00835_ vssd1 vssd1 vccd1 vccd1 net5202 sky130_fd_sc_hd__dlygate4sd3_1
X_22086_ net528 net586 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
Xhold3941 _01213_ vssd1 vssd1 vccd1 vccd1 net4468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4686 _00793_ vssd1 vssd1 vccd1 vccd1 net5213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3952 net2243 vssd1 vssd1 vccd1 vccd1 net4479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4697 net820 vssd1 vssd1 vccd1 vccd1 net5224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3963 rbzero.pov.ready_buffer\[66\] vssd1 vssd1 vccd1 vccd1 net4490 sky130_fd_sc_hd__buf_1
X_21037_ clknet_leaf_56_i_clk net5668 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3974 net8268 vssd1 vssd1 vccd1 vccd1 net4501 sky130_fd_sc_hd__clkbuf_4
Xhold3985 net3014 vssd1 vssd1 vccd1 vccd1 net4512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20624__354 clknet_1_0__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__inv_2
XFILLER_0_96_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3996 net8334 vssd1 vssd1 vccd1 vccd1 net4523 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__05742_ clknet_0__05742_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05742_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_199_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12810_ _05984_ _05981_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__or2_1
X_13790_ _06937_ _06938_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net54 _05912_ _05915_ net53 _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a221o_1
X_21939_ net381 net2523 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _08553_ _08554_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__xnor2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ net29 vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__buf_2
Xclkbuf_1_0__f__03506_ clknet_0__03506_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03506_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _07568_ _07577_ _07579_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__and3_1
X_11623_ _04755_ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__xnor2_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15391_ _08400_ _08485_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17130_ _09249_ net4914 vssd1 vssd1 vccd1 vccd1 _10150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14342_ _07308_ _07233_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__nor2_1
X_11554_ net1024 _04743_ net3983 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17061_ _10059_ _10081_ vssd1 vssd1 vccd1 vccd1 _10082_ sky130_fd_sc_hd__xnor2_1
X_10505_ net2790 net5598 _04053_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__mux2_1
X_14273_ _07336_ _07337_ _07290_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__a21o_1
X_11485_ net4126 net4748 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7290 net8535 vssd1 vssd1 vccd1 vccd1 net7817 sky130_fd_sc_hd__dlygate4sd3_1
X_16012_ _09101_ net7779 net3454 vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__a21o_1
X_13224_ _06392_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__or2_4
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13155_ _06265_ _06000_ _06001_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a31o_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ net3774 net2 net4067 _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a211o_1
X_17963_ _02198_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__xnor2_1
X_13086_ net2058 _06244_ _06255_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__o21ba_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19702_ net6562 net1447 _03468_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
X_16914_ _08338_ _08383_ _09935_ vssd1 vssd1 vccd1 vccd1 _09936_ sky130_fd_sc_hd__or3_1
X_12037_ rbzero.tex_r1\[23\] rbzero.tex_r1\[22\] _04979_ vssd1 vssd1 vccd1 vccd1 _05226_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17894_ _02130_ _02131_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19633_ net6315 net3838 _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
X_20599__331 clknet_1_0__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__inv_2
X_16845_ _09858_ _09859_ net3798 vssd1 vssd1 vccd1 vccd1 _09869_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16776_ _09805_ _09806_ vssd1 vssd1 vccd1 vccd1 _09807_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19564_ net6411 net1622 _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
X_13988_ net581 _07158_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15727_ _08341_ _08329_ _08246_ _08244_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__and4bb_1
X_18515_ _02676_ _02686_ _02690_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ net4644 net3985 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__or2b_2
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _03352_ net3521 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__nor2_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15658_ _08725_ _08751_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_186_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18446_ _02617_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__buf_2
XFILLER_0_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ _07608_ _07653_ _07655_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__a22o_1
X_18377_ net4554 rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _02562_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_29_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _08666_ _08245_ _08671_ _08670_ _08669_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _09537_ _10346_ vssd1 vssd1 vccd1 vccd1 _10347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ _09373_ net4909 vssd1 vssd1 vccd1 vccd1 _10278_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20270_ _03805_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3204 _02335_ vssd1 vssd1 vccd1 vccd1 net3731 sky130_fd_sc_hd__buf_1
XFILLER_0_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3215 net5841 vssd1 vssd1 vccd1 vccd1 net3742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3226 net5855 vssd1 vssd1 vccd1 vccd1 net3753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3237 net7950 vssd1 vssd1 vccd1 vccd1 net3764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2503 _04302_ vssd1 vssd1 vccd1 vccd1 net3030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3248 _07871_ vssd1 vssd1 vccd1 vccd1 net3775 sky130_fd_sc_hd__clkbuf_2
Xhold3259 net4925 vssd1 vssd1 vccd1 vccd1 net3786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 net5862 vssd1 vssd1 vccd1 vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2525 net2542 vssd1 vssd1 vccd1 vccd1 net3052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2536 net7539 vssd1 vssd1 vccd1 vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1802 _01525_ vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2547 _03554_ vssd1 vssd1 vccd1 vccd1 net3074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1813 net6980 vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 _03373_ vssd1 vssd1 vccd1 vccd1 net3085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 rbzero.tex_b1\[1\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 _03557_ vssd1 vssd1 vccd1 vccd1 net3096 sky130_fd_sc_hd__dlygate4sd3_1
X_19804__81 clknet_1_1__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__inv_2
Xhold1835 _01083_ vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1846 net7456 vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1857 net7140 vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 _01597_ vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1879 net6919 vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ clknet_leaf_103_i_clk net3582 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_91_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21655_ clknet_leaf_121_i_clk net3314 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21586_ net220 net2389 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_98 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_98/HI o_rgb[5] sky130_fd_sc_hd__conb_1
X_11270_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__nor2_2
Xhold5140 _00524_ vssd1 vssd1 vccd1 vccd1 net5667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5151 _04059_ vssd1 vssd1 vccd1 vccd1 net5678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5162 _04164_ vssd1 vssd1 vccd1 vccd1 net5689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5173 net5662 vssd1 vssd1 vccd1 vccd1 net5700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5184 _03049_ vssd1 vssd1 vccd1 vccd1 net5711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5195 net2968 vssd1 vssd1 vccd1 vccd1 net5722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4450 _00878_ vssd1 vssd1 vccd1 vccd1 net4977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4461 net715 vssd1 vssd1 vccd1 vccd1 net4988 sky130_fd_sc_hd__dlygate4sd3_1
X_22138_ clknet_leaf_85_i_clk net3873 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4472 net671 vssd1 vssd1 vccd1 vccd1 net4999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4483 _00866_ vssd1 vssd1 vccd1 vccd1 net5010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4494 net748 vssd1 vssd1 vccd1 vccd1 net5021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3771 net7923 vssd1 vssd1 vccd1 vccd1 net4298 sky130_fd_sc_hd__dlygate4sd3_1
X_14960_ _08077_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__clkbuf_1
X_22069_ net511 net2175 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold3782 net8160 vssd1 vssd1 vccd1 vccd1 net4309 sky130_fd_sc_hd__clkbuf_2
Xhold3793 net7927 vssd1 vssd1 vccd1 vccd1 net4320 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ _07047_ _07081_ _06706_ _07035_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a2bb2o_1
X_14891_ net4667 _08034_ _08036_ net3749 net4543 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__o221a_1
X_16630_ _04458_ net4122 vssd1 vssd1 vccd1 vccd1 _09719_ sky130_fd_sc_hd__or2_1
X_13842_ _07010_ _07011_ _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ _09530_ _09635_ _09649_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13773_ _06897_ _06898_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__xor2_1
X_10985_ net6874 net2857 _04309_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__mux2_1
X_15512_ _08605_ _08564_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__nand2_2
X_18300_ net1381 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
X_19280_ net4842 _03140_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__and2_1
X_12724_ net34 vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16492_ net7779 _09582_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18231_ _02446_ _02447_ _02052_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o21ai_1
X_15443_ _08526_ _08527_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ net26 _05809_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__nor2_1
X_18162_ _02382_ _02380_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15374_ _08453_ _08468_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__xor2_2
XFILLER_0_68_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12586_ net49 _05764_ _05765_ _05760_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17113_ _09788_ _10015_ _10016_ _10133_ vssd1 vssd1 vccd1 vccd1 _10134_ sky130_fd_sc_hd__a31o_1
Xclkbuf_0__03851_ _03851_ vssd1 vssd1 vccd1 vccd1 clknet_0__03851_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14325_ _07486_ _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__xor2_4
XFILLER_0_163_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18093_ _02326_ net4518 _02320_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ _04679_ net4357 net4393 _04657_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17044_ _09915_ _08616_ _10064_ vssd1 vssd1 vccd1 vccd1 _10065_ sky130_fd_sc_hd__or3_1
Xhold409 net5235 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ _07411_ _07425_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__nor2_1
X_11468_ net4126 net4160 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ net8217 _06374_ _06375_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__a31o_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14187_ _06726_ _07342_ _07344_ net8355 vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__a211o_1
X_11399_ _04553_ _04556_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__and2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ net8267 _06266_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ net5814 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17946_ _02181_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__nor2_1
X_13069_ _06028_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__buf_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 _00921_ vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17877_ _01760_ _09060_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19616_ net6253 net1493 _03430_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
X_16828_ _09850_ _09853_ vssd1 vssd1 vccd1 vccd1 _09854_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19547_ net2099 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
X_16759_ _09791_ _08978_ net89 vssd1 vssd1 vccd1 vccd1 _09792_ sky130_fd_sc_hd__a21oi_1
X_19478_ net5940 _03139_ _03344_ _02954_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18429_ net3494 net4501 _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20653__380 clknet_1_0__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__inv_2
X_21440_ clknet_leaf_26_i_clk net1495 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21371_ clknet_leaf_10_i_clk net4994 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20322_ net6319 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold910 _00582_ vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 net6427 vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 net6509 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold943 _00976_ vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
X_20253_ net4122 net7619 vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__and2_1
Xhold954 _03355_ vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3001 net5810 vssd1 vssd1 vccd1 vccd1 net3528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 net6475 vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _03829_ vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3012 _03769_ vssd1 vssd1 vccd1 vccd1 net3539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 net6362 vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3023 _00893_ vssd1 vssd1 vccd1 vccd1 net3550 sky130_fd_sc_hd__dlygate4sd3_1
X_20184_ net3565 net2943 _03723_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__mux2_1
Xhold998 _01013_ vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3034 rbzero.spi_registers.spi_buffer\[13\] vssd1 vssd1 vccd1 vccd1 net3561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2300 _04250_ vssd1 vssd1 vccd1 vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3045 _00886_ vssd1 vssd1 vccd1 vccd1 net3572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2311 net3137 vssd1 vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3056 net7600 vssd1 vssd1 vccd1 vccd1 net3583 sky130_fd_sc_hd__clkbuf_2
Xhold2322 net7006 vssd1 vssd1 vccd1 vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3067 _00737_ vssd1 vssd1 vccd1 vccd1 net3594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3078 net5971 vssd1 vssd1 vccd1 vccd1 net3605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2333 net3282 vssd1 vssd1 vccd1 vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03840_ clknet_0__03840_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03840_
+ sky130_fd_sc_hd__clkbuf_16
Xhold2344 _01098_ vssd1 vssd1 vccd1 vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3089 net4870 vssd1 vssd1 vccd1 vccd1 net3616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2355 _01546_ vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 net6131 vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2366 _04447_ vssd1 vssd1 vccd1 vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1621 _00923_ vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 net6907 vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2377 _03584_ vssd1 vssd1 vccd1 vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2388 _04109_ vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 net7118 vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1654 _01110_ vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2399 rbzero.pov.spi_buffer\[64\] vssd1 vssd1 vccd1 vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1665 _01152_ vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1676 _01526_ vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1687 net2631 vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1698 _00941_ vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ net6812 net7091 _04194_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xsplit47 _06433_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_1
XFILLER_0_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21707_ clknet_leaf_119_i_clk net4377 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12440_ net7726 _05624_ net7570 vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__mux2_1
X_21638_ clknet_leaf_127_i_clk net1153 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12371_ _05306_ _05551_ _05555_ _04967_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_164_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21569_ net203 net2727 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__clkbuf_4
X_11322_ rbzero.spi_registers.texadd3\[11\] rbzero.spi_registers.texadd1\[11\] rbzero.spi_registers.texadd0\[11\]
+ rbzero.spi_registers.texadd2\[11\] _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04514_
+ sky130_fd_sc_hd__mux4_2
X_15090_ _08118_ _08183_ _08184_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__a21o_4
XFILLER_0_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14041_ _06673_ _06695_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__or2_1
X_11253_ net7113 net2895 _04445_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11184_ net7059 net2841 _04412_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
Xhold4280 _02883_ vssd1 vssd1 vccd1 vccd1 net4807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17800_ _02037_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4291 net1022 vssd1 vssd1 vccd1 vccd1 net4818 sky130_fd_sc_hd__dlygate4sd3_1
X_20481__225 clknet_1_0__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__inv_2
X_15992_ _09084_ net7769 vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__or2_1
X_18780_ _02911_ _02927_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__xnor2_1
Xhold3590 _05062_ vssd1 vssd1 vccd1 vccd1 net4117 sky130_fd_sc_hd__dlygate4sd3_1
X_17731_ _01916_ _01892_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__or2b_1
X_14943_ net3822 _07870_ _08068_ vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__mux2_1
X_17662_ _01900_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14874_ _08026_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19401_ net5460 _03302_ _03305_ _03299_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__o211a_1
X_16613_ _09701_ _09702_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__xor2_1
X_13825_ _06993_ _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__xnor2_2
X_17593_ _01831_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16544_ _09507_ _09517_ _09515_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__a21o_1
X_19332_ net5069 _03235_ _03264_ _03259_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__o211a_1
X_13756_ _06893_ _06895_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ net6197 net1715 _04298_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12707_ _05862_ _05884_ net31 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21bo_1
X_16475_ _09390_ _09434_ _09433_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__a21oi_1
X_19263_ net6347 _03217_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13687_ _06813_ _06698_ _06856_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__o21ai_1
X_10899_ net7279 net7057 _04265_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__mux2_1
X_15426_ _08486_ _08520_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__xor2_1
X_18214_ _02432_ net3803 _02393_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19194_ net1923 _03183_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__or2_1
X_12638_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__and2b_1
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15357_ _08444_ _08451_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__xor2_2
X_18145_ _02365_ _02366_ _02367_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__o21a_1
X_12569_ net16 vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5909 net1244 vssd1 vssd1 vccd1 vccd1 net6436 sky130_fd_sc_hd__dlygate4sd3_1
X_14308_ _07463_ _07478_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18076_ _02150_ _02153_ _02236_ _02253_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a311oi_1
X_15288_ _08119_ _08381_ _08382_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__a21o_4
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold206 net5096 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 net8347 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 net7926 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ _10046_ _10047_ vssd1 vssd1 vccd1 vccd1 _10048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 net6083 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ _07394_ _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ net5735 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _10062_ _09666_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__or2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20940_ clknet_leaf_77_i_clk net4740 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20871_ net4887 _02508_ _02559_ _04007_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7801 rbzero.wall_tracer.stepDistX\[1\] vssd1 vssd1 vccd1 vccd1 net8328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7812 net4623 vssd1 vssd1 vccd1 vccd1 net8339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7823 rbzero.wall_tracer.stepDistX\[-7\] vssd1 vssd1 vccd1 vccd1 net8350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7834 _06632_ vssd1 vssd1 vccd1 vccd1 net8361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7845 _08163_ vssd1 vssd1 vccd1 vccd1 net8372 sky130_fd_sc_hd__dlygate4sd3_1
X_21423_ clknet_leaf_18_i_clk net3904 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_sky
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7856 _09886_ vssd1 vssd1 vccd1 vccd1 net8383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7867 rbzero.wall_tracer.stepDistY\[0\] vssd1 vssd1 vccd1 vccd1 net8394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7878 net4652 vssd1 vssd1 vccd1 vccd1 net8405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7889 net4582 vssd1 vssd1 vccd1 vccd1 net8416 sky130_fd_sc_hd__dlygate4sd3_1
X_21354_ clknet_leaf_10_i_clk net5262 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20305_ net6446 net3838 _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
X_21285_ clknet_leaf_24_i_clk net5434 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold740 net6322 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_20430__179 clknet_1_1__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__inv_2
Xhold751 net6280 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 net6481 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold773 _01339_ vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
X_20236_ net5045 _03706_ _03780_ _03765_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__o211a_1
Xhold784 _03459_ vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 net6308 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167_ rbzero.debug_overlay.facingY\[-4\] _03711_ vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__or2_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2130 rbzero.tex_r1\[42\] vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2141 _04334_ vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2152 net7124 vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2163 _01585_ vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
X_20098_ net4436 net4748 _03682_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_110_i_clk clknet_4_6__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2174 _04185_ vssd1 vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1440 net6903 vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2185 net7448 vssd1 vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 _01590_ vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2196 _04289_ vssd1 vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ net4436 _05110_ _05116_ net3552 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1462 net5593 vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1473 net6763 vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1484 net7160 vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _01550_ vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ net5911 _04666_ net5205 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__o21ai_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13610_ net555 _06759_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and2_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ net6480 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_125_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _07751_ _07757_ _07760_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__o21ai_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13541_ _06707_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__nor2_1
X_10753_ net6468 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16260_ _09133_ _09351_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _06436_ _06637_ _06638_ _06642_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_164_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ net6490 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _08305_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ _04922_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16191_ _09156_ _09273_ _09282_ vssd1 vssd1 vccd1 vccd1 _09284_ sky130_fd_sc_hd__nand3_1
XFILLER_0_164_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15142_ net3419 _08196_ net3339 vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__o21ai_1
X_12354_ net7720 _05539_ net7570 vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ net3954 _04495_ net3641 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__or3_1
X_15073_ net4776 _08162_ _08167_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19950_ net3287 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
X_12285_ _04976_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18901_ net3057 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
X_14024_ _06699_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__or2_1
X_11236_ _04103_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__clkbuf_4
X_19881_ net2312 vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__clkbuf_4
X_18832_ net3911 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__clkbuf_1
X_11167_ net6788 net2804 _04401_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__mux2_1
X_18763_ _02865_ net4560 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _09057_ _09058_ _09069_ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_175_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11098_ net2978 net5586 _04364_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
X_17714_ _01851_ _01852_ _01953_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14926_ net8270 _08047_ _04482_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18694_ net4560 net3619 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17645_ _01882_ _01883_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__and2_1
X_14857_ net7846 _07987_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _06961_ _06975_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17576_ _01815_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and2_1
X_14788_ _07881_ _07884_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19315_ net5316 _03250_ _03255_ _03246_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__o211a_1
X_16527_ _08185_ _09351_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__and2_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ _06883_ _06908_ _06909_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246_ net6351 _03203_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__or2_1
X_16458_ _09548_ _09417_ _08474_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7108 net3473 vssd1 vssd1 vccd1 vccd1 net7635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7119 net3712 vssd1 vssd1 vccd1 vccd1 net7646 sky130_fd_sc_hd__dlygate4sd3_1
X_15409_ _08502_ _08503_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__xor2_1
Xhold6407 net2073 vssd1 vssd1 vccd1 vccd1 net6934 sky130_fd_sc_hd__dlygate4sd3_1
X_16389_ _08226_ _08614_ _09355_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19177_ net6448 _03170_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or2_1
Xhold6418 rbzero.tex_b0\[62\] vssd1 vssd1 vccd1 vccd1 net6945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6429 net2149 vssd1 vssd1 vccd1 vccd1 net6956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18128_ _02350_ _02351_ _02352_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__o21a_1
Xhold5706 net1169 vssd1 vssd1 vccd1 vccd1 net6233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5717 _04197_ vssd1 vssd1 vccd1 vccd1 net6244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5728 net1212 vssd1 vssd1 vccd1 vccd1 net6255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5739 rbzero.tex_b1\[0\] vssd1 vssd1 vccd1 vccd1 net6266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18059_ _08612_ _09410_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21070_ clknet_leaf_80_i_clk _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20021_ _03615_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21972_ net414 net2419 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer10 _06987_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 _06978_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_i_clk clknet_4_9__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xrebuffer32 _06902_ vssd1 vssd1 vccd1 vccd1 net3463 sky130_fd_sc_hd__buf_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20923_ clknet_leaf_69_i_clk _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer43 _06395_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__dlygate4sd3_1
Xrebuffer54 _06694_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20854_ net4211 _04001_ _04002_ _09209_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a22o_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20785_ net1038 net5581 vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_i_clk clknet_4_14__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7620 rbzero.spi_registers.vshift\[2\] vssd1 vssd1 vccd1 vccd1 net8147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7631 rbzero.map_overlay.i_otherx\[2\] vssd1 vssd1 vccd1 vccd1 net8158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7642 rbzero.map_overlay.i_mapdy\[2\] vssd1 vssd1 vccd1 vccd1 net8169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7653 rbzero.traced_texa\[0\] vssd1 vssd1 vccd1 vccd1 net8180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7664 rbzero.traced_texa\[-10\] vssd1 vssd1 vccd1 vccd1 net8191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6930 net2373 vssd1 vssd1 vccd1 vccd1 net7457 sky130_fd_sc_hd__dlygate4sd3_1
X_21406_ clknet_leaf_36_i_clk net3550 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7675 _08040_ vssd1 vssd1 vccd1 vccd1 net8202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6941 rbzero.tex_r0\[46\] vssd1 vssd1 vccd1 vccd1 net7468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7686 net8519 vssd1 vssd1 vccd1 vccd1 net8213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6952 net2901 vssd1 vssd1 vccd1 vccd1 net7479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7697 rbzero.debug_overlay.playerY\[-2\] vssd1 vssd1 vccd1 vccd1 net8224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6963 net645 vssd1 vssd1 vccd1 vccd1 net7490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6974 rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net7501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6985 net3346 vssd1 vssd1 vccd1 vccd1 net7512 sky130_fd_sc_hd__dlygate4sd3_1
X_21337_ clknet_leaf_6_i_clk net5111 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6996 rbzero.spi_registers.new_other\[9\] vssd1 vssd1 vccd1 vccd1 net7523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12070_ rbzero.tex_r1\[41\] rbzero.tex_r1\[40\] _05258_ vssd1 vssd1 vccd1 vccd1 _05259_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21268_ clknet_leaf_122_i_clk net3043 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold570 _01656_ vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 net5475 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 net5457 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net2667 net6894 _04331_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20219_ net3540 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21199_ clknet_leaf_127_i_clk net1934 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _08763_ _08809_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__xnor2_4
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _04718_ net4034 net3807 _04721_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__o221a_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 net6656 vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1281 net1865 vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ net4168 _05106_ _05108_ net3419 _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a221o_1
X_14711_ net7795 _07854_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1292 net6803 vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _08783_ _08784_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__nand2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _10327_ _09403_ _10322_ _01671_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__o31a_1
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _07800_ _07811_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__or2_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _05043_ net4127 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__or2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20593__326 clknet_1_0__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__inv_2
XFILLER_0_200_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ net2516 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _10266_ _10268_ _10377_ _10379_ vssd1 vssd1 vccd1 vccd1 _10380_ sky130_fd_sc_hd__a31o_2
X_14573_ _07742_ _07743_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__xnor2_1
X_11785_ _04971_ _04974_ _04955_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19100_ net5755 _03125_ net2629 _03128_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16312_ _08180_ _09288_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__nand2_1
X_13524_ _06577_ _06694_ net83 vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__a21o_2
X_17292_ _10276_ _10310_ vssd1 vssd1 vccd1 vccd1 _10311_ sky130_fd_sc_hd__xnor2_2
X_10736_ net2244 net6227 _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16243_ _09323_ _09325_ _09321_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__o21ai_4
X_19031_ net3816 net3402 _03078_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
X_13455_ _06550_ _06612_ _06613_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__and3_1
X_10667_ net6842 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _05250_ vssd1 vssd1 vccd1 vccd1 _05591_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16174_ _09264_ _09265_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13386_ _06538_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__buf_2
X_10598_ net1843 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15125_ _06119_ _08216_ _08217_ _08219_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__a2bb2o_2
X_12337_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _05249_ vssd1 vssd1 vccd1 vccd1 _05523_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19933_ net1111 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
X_15056_ rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\] _06349_
+ _06340_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12268_ net7734 _05454_ net7570 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14007_ _07151_ _07128_ _07176_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__nand3_1
X_11219_ net1825 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__clkbuf_1
X_19864_ net3187 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
X_12199_ rbzero.tex_g1\[9\] rbzero.tex_g1\[8\] _04924_ vssd1 vssd1 vccd1 vccd1 _05386_
+ sky130_fd_sc_hd__mux2_1
X_18815_ net3084 _02955_ _02956_ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a31o_1
XFILLER_0_208_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ _02865_ net3678 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nand2_1
X_15958_ _08521_ _08563_ _09052_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__a21oi_1
X_14909_ net3888 _08034_ _08036_ net3785 net4730 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18677_ _02830_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nor2_1
X_15889_ _08810_ _08856_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17628_ _01865_ _01866_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17559_ _01798_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19229_ net5264 _03201_ _03204_ _03206_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__o211a_1
Xhold6204 net1618 vssd1 vssd1 vccd1 vccd1 net6731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6215 net1238 vssd1 vssd1 vccd1 vccd1 net6742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6226 rbzero.tex_r1\[22\] vssd1 vssd1 vccd1 vccd1 net6753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6237 net2000 vssd1 vssd1 vccd1 vccd1 net6764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5503 net633 vssd1 vssd1 vccd1 vccd1 net6030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6248 rbzero.tex_g0\[17\] vssd1 vssd1 vccd1 vccd1 net6775 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__05898_ _05898_ vssd1 vssd1 vccd1 vccd1 clknet_0__05898_ sky130_fd_sc_hd__clkbuf_16
Xhold6259 net1986 vssd1 vssd1 vccd1 vccd1 net6786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5514 net678 vssd1 vssd1 vccd1 vccd1 net6041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5525 net660 vssd1 vssd1 vccd1 vccd1 net6052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5536 net3554 vssd1 vssd1 vccd1 vccd1 net6063 sky130_fd_sc_hd__dlygate4sd3_1
X_22171_ clknet_leaf_89_i_clk net680 vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold5547 net643 vssd1 vssd1 vccd1 vccd1 net6074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4802 _00527_ vssd1 vssd1 vccd1 vccd1 net5329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5558 _04150_ vssd1 vssd1 vccd1 vccd1 net6085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4813 net915 vssd1 vssd1 vccd1 vccd1 net5340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5569 net904 vssd1 vssd1 vccd1 vccd1 net6096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4824 rbzero.spi_registers.texadd1\[3\] vssd1 vssd1 vccd1 vccd1 net5351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4835 net954 vssd1 vssd1 vccd1 vccd1 net5362 sky130_fd_sc_hd__dlygate4sd3_1
X_21122_ clknet_leaf_106_i_clk net3736 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4846 _00796_ vssd1 vssd1 vccd1 vccd1 net5373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4857 net848 vssd1 vssd1 vccd1 vccd1 net5384 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold4868 rbzero.spi_registers.texadd3\[6\] vssd1 vssd1 vccd1 vccd1 net5395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4879 net831 vssd1 vssd1 vccd1 vccd1 net5406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21053_ clknet_leaf_74_i_clk _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20004_ net3348 _03607_ net5837 _03339_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21955_ net397 net2431 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ clknet_leaf_61_i_clk _00393_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ net328 net644 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _03995_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__buf_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ net3189 _04758_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a21boi_1
X_20768_ _03936_ _03937_ _03938_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ net2798 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20699_ _03109_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__clkbuf_4
X_20436__185 clknet_1_0__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__inv_2
Xhold7450 rbzero.wall_tracer.trackDistX\[0\] vssd1 vssd1 vccd1 vccd1 net7977 sky130_fd_sc_hd__dlygate4sd3_1
X_13240_ _06385_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__nor2_1
X_10452_ net2394 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__clkbuf_1
Xhold7461 net4546 vssd1 vssd1 vccd1 vccd1 net7988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7472 net4690 vssd1 vssd1 vccd1 vccd1 net7999 sky130_fd_sc_hd__clkbuf_2
Xhold7483 _00514_ vssd1 vssd1 vccd1 vccd1 net8010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7494 net4576 vssd1 vssd1 vccd1 vccd1 net8021 sky130_fd_sc_hd__buf_2
Xhold6760 net2786 vssd1 vssd1 vccd1 vccd1 net7287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13171_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__mux2_4
Xhold6771 rbzero.tex_r0\[31\] vssd1 vssd1 vccd1 vccd1 net7298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6782 rbzero.pov.spi_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net7309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6793 net2892 vssd1 vssd1 vccd1 vccd1 net7320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12122_ _05308_ _05309_ _04911_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16930_ _09933_ _09951_ vssd1 vssd1 vccd1 vccd1 _09952_ sky130_fd_sc_hd__xor2_1
X_12053_ _04911_ _05238_ _05241_ _04919_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__o211a_1
X_11004_ net3163 net7389 _04320_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
X_16861_ net4669 net4373 vssd1 vssd1 vccd1 vccd1 _09883_ sky130_fd_sc_hd__or2_1
X_18600_ _02751_ _02759_ net4529 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__o21a_1
XFILLER_0_205_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15812_ _08277_ _08474_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__nor2_1
X_19580_ net7085 net3402 _03403_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
X_16792_ net4648 vssd1 vssd1 vccd1 vccd1 _09822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20601__333 clknet_1_1__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__inv_2
X_18531_ net4603 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__inv_2
X_15743_ _08253_ _08254_ _08433_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__and3_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _06068_ net4007 _06129_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and4_1
XFILLER_0_198_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _05079_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor2_4
XFILLER_0_169_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18462_ _02617_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02641_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15674_ _08243_ _08433_ _08768_ _08732_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__a22o_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ net3964 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__inv_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _10344_ _10337_ vssd1 vssd1 vccd1 vccd1 _10431_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11837_ net1822 net4271 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__nand2_1
X_14625_ _07793_ _07795_ _07339_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__o21a_1
X_18393_ _02575_ _02576_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__nand2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _10361_ _10362_ _10233_ _10235_ vssd1 vssd1 vccd1 vccd1 _10363_ sky130_fd_sc_hd__o31a_1
X_14556_ _07725_ _07723_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__or2b_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _04921_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ net5601 net2793 _04171_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux2_1
X_13507_ _06493_ _06572_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__nand2_1
X_17275_ _10190_ _08383_ _08614_ _09062_ vssd1 vssd1 vccd1 vccd1 _10294_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ _07308_ _07327_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__or3_1
X_11699_ _04886_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19014_ net3397 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__buf_4
X_16226_ _09070_ _09202_ _09201_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__a21oi_1
X_13438_ _06398_ net82 _06525_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer1 _06536_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_1
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16157_ _08996_ _09135_ _09249_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13369_ _06538_ net81 vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__xnor2_4
Xhold4109 _03768_ vssd1 vssd1 vccd1 vccd1 net4636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ net4379 _08123_ _08148_ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__a21o_1
X_16088_ net8033 _09181_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__nor2_1
Xhold3408 net7694 vssd1 vssd1 vccd1 vccd1 net3935 sky130_fd_sc_hd__clkbuf_2
X_19916_ net3139 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
X_15039_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] net4181
+ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2707 _03552_ vssd1 vssd1 vccd1 vccd1 net3234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2718 _01297_ vssd1 vssd1 vccd1 vccd1 net3245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2729 net3073 vssd1 vssd1 vccd1 vccd1 net3256 sky130_fd_sc_hd__dlygate4sd3_1
X_19847_ net2772 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ _02856_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20576__310 clknet_1_0__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__inv_2
X_21740_ clknet_leaf_99_i_clk net4557 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21671_ clknet_leaf_123_i_clk net1262 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6001 net1602 vssd1 vssd1 vccd1 vccd1 net6528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6012 _04421_ vssd1 vssd1 vccd1 vccd1 net6539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6023 net1527 vssd1 vssd1 vccd1 vccd1 net6550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6034 rbzero.spi_registers.new_texadd\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net6561
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6045 net1686 vssd1 vssd1 vccd1 vccd1 net6572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5300 _03633_ vssd1 vssd1 vccd1 vccd1 net5827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6056 net1606 vssd1 vssd1 vccd1 vccd1 net6583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5311 _01169_ vssd1 vssd1 vccd1 vccd1 net5838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6067 _04255_ vssd1 vssd1 vccd1 vccd1 net6594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5322 net3266 vssd1 vssd1 vccd1 vccd1 net5849 sky130_fd_sc_hd__buf_1
Xhold6078 net1719 vssd1 vssd1 vccd1 vccd1 net6605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5333 _01184_ vssd1 vssd1 vccd1 vccd1 net5860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5344 net3444 vssd1 vssd1 vccd1 vccd1 net5871 sky130_fd_sc_hd__dlygate4sd3_1
X_20672__17 clknet_1_1__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
Xhold6089 _04186_ vssd1 vssd1 vccd1 vccd1 net6616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4610 net787 vssd1 vssd1 vccd1 vccd1 net5137 sky130_fd_sc_hd__dlygate4sd3_1
X_22154_ clknet_leaf_54_i_clk _01641_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5366 _00607_ vssd1 vssd1 vccd1 vccd1 net5893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4621 rbzero.spi_registers.texadd0\[17\] vssd1 vssd1 vccd1 vccd1 net5148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5377 net3419 vssd1 vssd1 vccd1 vccd1 net5904 sky130_fd_sc_hd__buf_1
Xhold4632 net741 vssd1 vssd1 vccd1 vccd1 net5159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4643 _00820_ vssd1 vssd1 vccd1 vccd1 net5170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5388 net3389 vssd1 vssd1 vccd1 vccd1 net5915 sky130_fd_sc_hd__buf_1
XFILLER_0_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5399 _02778_ vssd1 vssd1 vccd1 vccd1 net5926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4654 net828 vssd1 vssd1 vccd1 vccd1 net5181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3920 _03727_ vssd1 vssd1 vccd1 vccd1 net4447 sky130_fd_sc_hd__dlygate4sd3_1
X_21105_ clknet_leaf_4_i_clk net1345 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4665 rbzero.spi_registers.texadd3\[2\] vssd1 vssd1 vccd1 vccd1 net5192 sky130_fd_sc_hd__dlygate4sd3_1
X_22085_ net527 net3242 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
Xhold3931 net7879 vssd1 vssd1 vccd1 vccd1 net4458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4676 net845 vssd1 vssd1 vccd1 vccd1 net5203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3942 net1060 vssd1 vssd1 vccd1 vccd1 net4469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4687 net825 vssd1 vssd1 vccd1 vccd1 net5214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3953 net7826 vssd1 vssd1 vccd1 vccd1 net4480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4698 _00870_ vssd1 vssd1 vccd1 vccd1 net5225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3964 _03629_ vssd1 vssd1 vccd1 vccd1 net4491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3975 _03754_ vssd1 vssd1 vccd1 vccd1 net4502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21036_ clknet_leaf_31_i_clk net5556 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3986 rbzero.debug_overlay.facingX\[0\] vssd1 vssd1 vccd1 vccd1 net4513 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3997 net3724 vssd1 vssd1 vccd1 vccd1 net4524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ net52 _05902_ _05916_ net55 vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a22o_1
X_21938_ net380 net1963 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ net32 net33 vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor2_1
X_21869_ net311 net3031 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _07534_ _07550_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _04757_ _04760_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15390_ _08470_ _08484_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14341_ _07503_ _07502_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__xor2_1
X_11553_ net4431 net4420 net4369 net4354 vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17060_ _10079_ _10080_ vssd1 vssd1 vccd1 vccd1 _10081_ sky130_fd_sc_hd__nand2_1
X_10504_ net5679 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__clkbuf_1
X_14272_ _06696_ _07281_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__nor3b_1
X_11484_ net3473 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__inv_2
X_16011_ _09101_ net7779 vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7280 net8441 vssd1 vssd1 vccd1 vccd1 net7807 sky130_fd_sc_hd__dlygate4sd3_1
X_13223_ _06378_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__xnor2_4
Xhold7291 net4891 vssd1 vssd1 vccd1 vccd1 net7818 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6590 net2747 vssd1 vssd1 vccd1 vccd1 net7117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13154_ net4236 net8051 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ net4172 _05293_ _04656_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17962_ _10190_ net7818 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__nand2_1
X_13085_ _06241_ _06256_ _06257_ _06242_ net5618 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__a32o_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19701_ net6631 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__clkbuf_1
X_16913_ _08142_ _08374_ vssd1 vssd1 vccd1 vccd1 _09935_ sky130_fd_sc_hd__or2_1
X_12036_ rbzero.tex_r1\[21\] rbzero.tex_r1\[20\] _04838_ vssd1 vssd1 vccd1 vccd1 _05225_
+ sky130_fd_sc_hd__mux2_1
X_17893_ _02031_ _02098_ _02129_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19632_ _03429_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__buf_4
X_16844_ net4665 net4471 vssd1 vssd1 vccd1 vccd1 _09868_ sky130_fd_sc_hd__nand2_2
X_19563_ net1779 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__clkbuf_4
X_16775_ net3945 net4353 vssd1 vssd1 vccd1 vccd1 _09806_ sky130_fd_sc_hd__nand2_1
X_13987_ _07152_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__xnor2_2
X_18514_ _02673_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__xnor2_1
X_15726_ _08819_ _08820_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__xor2_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ net3984 _06113_ _06093_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__or3b_1
X_19494_ net1879 _02472_ _03344_ _03141_ net3520 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o32a_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18445_ _02617_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _02625_
+ sky130_fd_sc_hd__xor2_1
X_15657_ _08726_ _08750_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _06038_ _06042_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ _07609_ _07693_ _07776_ _07778_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__a22o_1
X_18376_ net4554 rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _02561_
+ sky130_fd_sc_hd__nand2_1
X_15588_ _08679_ _08682_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17327_ _09976_ vssd1 vssd1 vccd1 vccd1 _10346_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14539_ _07701_ _07709_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17258_ _10206_ _10183_ vssd1 vssd1 vccd1 vccd1 _10277_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16209_ _09299_ _09301_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17189_ _10098_ _10099_ vssd1 vssd1 vccd1 vccd1 _10209_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3205 _02345_ vssd1 vssd1 vccd1 vccd1 net3732 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3216 net5843 vssd1 vssd1 vccd1 vccd1 net3743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3227 net5857 vssd1 vssd1 vccd1 vccd1 net3754 sky130_fd_sc_hd__dlygate4sd3_1
X_20608__339 clknet_1_0__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__inv_2
Xhold3238 net4910 vssd1 vssd1 vccd1 vccd1 net3765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2504 _01356_ vssd1 vssd1 vccd1 vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3249 net8366 vssd1 vssd1 vccd1 vccd1 net3776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _03116_ vssd1 vssd1 vccd1 vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2526 _03575_ vssd1 vssd1 vccd1 vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2537 _03536_ vssd1 vssd1 vccd1 vccd1 net3064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 _01119_ vssd1 vssd1 vccd1 vccd1 net3075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1803 net3259 vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1814 _01486_ vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 _03374_ vssd1 vssd1 vccd1 vccd1 net3086 sky130_fd_sc_hd__buf_4
Xhold1825 net5681 vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1836 rbzero.pov.ready_buffer\[19\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1847 net5638 vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 _04115_ vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 net7566 vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21723_ clknet_leaf_103_i_clk net3506 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21654_ clknet_leaf_121_i_clk net3123 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20605_ clknet_1_1__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__buf_1
XFILLER_0_191_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21585_ net219 net2541 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
X_20353__109 clknet_1_0__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__inv_2
XFILLER_0_90_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_99 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_99/HI o_rgb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5130 net900 vssd1 vssd1 vccd1 vccd1 net5657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5141 net2380 vssd1 vssd1 vccd1 vccd1 net5668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5152 net3241 vssd1 vssd1 vccd1 vccd1 net5679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5163 net1125 vssd1 vssd1 vccd1 vccd1 net5690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5174 _04245_ vssd1 vssd1 vccd1 vccd1 net5701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4440 rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 net4967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5185 net2194 vssd1 vssd1 vccd1 vccd1 net5712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5196 _00526_ vssd1 vssd1 vccd1 vccd1 net5723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4451 net706 vssd1 vssd1 vccd1 vccd1 net4978 sky130_fd_sc_hd__dlygate4sd3_1
X_22137_ clknet_leaf_85_i_clk net3977 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4462 _00875_ vssd1 vssd1 vccd1 vccd1 net4989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4473 rbzero.spi_registers.texadd3\[13\] vssd1 vssd1 vccd1 vccd1 net5000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4484 net728 vssd1 vssd1 vccd1 vccd1 net5011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20548__286 clknet_1_0__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__inv_2
Xhold3750 rbzero.wall_tracer.visualWallDist\[-7\] vssd1 vssd1 vccd1 vccd1 net4277
+ sky130_fd_sc_hd__buf_2
Xhold4495 _00865_ vssd1 vssd1 vccd1 vccd1 net5022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3761 net7933 vssd1 vssd1 vccd1 vccd1 net4288 sky130_fd_sc_hd__dlygate4sd3_1
X_22068_ net510 net1993 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold3772 rbzero.wall_tracer.visualWallDist\[1\] vssd1 vssd1 vccd1 vccd1 net4299 sky130_fd_sc_hd__buf_1
Xhold3783 _00757_ vssd1 vssd1 vccd1 vccd1 net4310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3794 net8148 vssd1 vssd1 vccd1 vccd1 net4321 sky130_fd_sc_hd__clkbuf_2
X_21019_ clknet_leaf_57_i_clk net4282 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13910_ _07079_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__and2_1
X_14890_ rbzero.wall_tracer.visualWallDist\[-11\] _08037_ _08038_ vssd1 vssd1 vccd1
+ vccd1 _08039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13841_ _06719_ _06702_ _06705_ net79 vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__or4_1
XFILLER_0_187_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _09530_ _09635_ _09649_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__a21o_1
X_13772_ _06940_ _06941_ _06942_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a21oi_1
X_10984_ net6635 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _08564_ _08605_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__nor2_2
XFILLER_0_168_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ net38 net39 vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__or2_1
X_16491_ _09453_ _09455_ _09452_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18230_ _02444_ _02445_ _09845_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a21o_1
X_15442_ _08532_ _08536_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ _05831_ _05832_ net25 vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11605_ _04783_ _04786_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__xnor2_1
X_18161_ _02386_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15373_ _08456_ _08467_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__nand2_1
X_12585_ net50 _05747_ _05749_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__and3_1
XFILLER_0_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17112_ _08103_ _10132_ vssd1 vssd1 vccd1 vccd1 _10133_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__03850_ _03850_ vssd1 vssd1 vccd1 vccd1 clknet_0__03850_ sky130_fd_sc_hd__clkbuf_16
X_14324_ _07488_ _07494_ _07493_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_68_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _04708_ _04715_ net4153 _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or4_1
X_18092_ _06058_ net3701 _09801_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17043_ _09935_ _10063_ vssd1 vssd1 vccd1 vccd1 _10064_ sky130_fd_sc_hd__xor2_1
X_14255_ _07411_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11467_ net4176 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ net8051 _05992_ _05994_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__o31a_1
X_14186_ _07352_ _07356_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or2_1
X_11398_ _04503_ _04561_ _04586_ _04589_ _04584_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__o311a_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _06264_ _06267_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a21oi_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ net5812 net4490 _03058_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _02165_ _02180_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__nor2_1
X_13068_ net5531 _06028_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__xor2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _05206_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17876_ _02016_ _02017_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19615_ net1378 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__clkbuf_1
X_16827_ _09851_ _09852_ vssd1 vssd1 vccd1 vccd1 _09853_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19546_ net2098 net1426 _03388_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__mux2_1
X_16758_ _08979_ _08934_ vssd1 vssd1 vccd1 vccd1 _09791_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15709_ _08797_ _08802_ _08803_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__a21bo_1
X_19477_ _04459_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16689_ net8138 _09743_ _09744_ net4236 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18428_ _02607_ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18359_ _02541_ _02544_ _04489_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21370_ clknet_leaf_10_i_clk net5195 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20321_ net6317 net3866 _03825_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold900 _03378_ vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 net5705 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold922 _00591_ vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 _03819_ vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_20252_ net4092 _03792_ net4071 _03788_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__or4b_1
Xhold944 net3158 vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 _00911_ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold966 _02481_ vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__buf_4
Xhold3002 rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 net3529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _01267_ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3013 _03770_ vssd1 vssd1 vccd1 vccd1 net3540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3024 net8380 vssd1 vssd1 vccd1 vccd1 net3551 sky130_fd_sc_hd__dlygate4sd3_1
X_20183_ net4004 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
Xhold988 net6364 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 net6547 vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3035 net1655 vssd1 vssd1 vccd1 vccd1 net3562 sky130_fd_sc_hd__buf_2
Xhold2301 _01402_ vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3046 net8391 vssd1 vssd1 vccd1 vccd1 net3573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3057 net7598 vssd1 vssd1 vccd1 vccd1 net3584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 _03043_ vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2323 _01416_ vssd1 vssd1 vccd1 vccd1 net2850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3068 rbzero.spi_registers.spi_buffer\[12\] vssd1 vssd1 vccd1 vccd1 net3595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3079 _00603_ vssd1 vssd1 vccd1 vccd1 net3606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2334 _03581_ vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1600 _00663_ vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2345 net3949 vssd1 vssd1 vccd1 vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2356 net2977 vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 net6133 vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2367 _01032_ vssd1 vssd1 vccd1 vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1622 net6955 vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1633 _01527_ vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 _01146_ vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2389 _01530_ vssd1 vssd1 vccd1 vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 _04443_ vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1655 net7495 vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1666 net5709 vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1677 net7750 vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1688 net5590 vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1699 net6817 vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21706_ clknet_leaf_118_i_clk net4438 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21637_ clknet_leaf_125_i_clk net2936 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _05517_ _05552_ _05554_ _05465_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__o211a_1
X_20554__290 clknet_1_0__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__inv_2
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21568_ net202 net1714 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _04511_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21499_ clknet_leaf_3_i_clk net1333 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _07105_ _07106_ _07157_ _07158_ _06694_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__a32o_1
X_11252_ net6971 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ net2382 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__clkbuf_1
Xhold4270 _02857_ vssd1 vssd1 vccd1 vccd1 net4797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4281 _02884_ vssd1 vssd1 vccd1 vccd1 net4808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15991_ _09084_ net7769 vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17730_ _01871_ _01886_ _01884_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a21o_1
Xhold3580 _05068_ vssd1 vssd1 vccd1 vccd1 net4107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3591 net7563 vssd1 vssd1 vccd1 vccd1 net4118 sky130_fd_sc_hd__dlymetal6s2s_1
X_14942_ _08067_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__buf_4
X_17661_ _01898_ _01899_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__or2_1
Xhold2890 net5928 vssd1 vssd1 vccd1 vccd1 net3417 sky130_fd_sc_hd__buf_2
X_14873_ net4537 _08025_ _07976_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__mux2_1
X_19400_ net1643 _03303_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16612_ _09498_ _09568_ _09567_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__a21oi_1
X_19795__73 clknet_1_0__leaf__03511_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
X_13824_ _06926_ net533 _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a21bo_1
X_17592_ _10428_ _01708_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ net1505 _03237_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__or2_1
X_16543_ _09597_ _09632_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10967_ net1873 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
X_13755_ _06707_ _06922_ _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19262_ net5320 _03216_ _03224_ _03219_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ net51 net41 net40 _05203_ _05850_ _05851_ vssd1 vssd1 vccd1 vccd1 _05884_
+ sky130_fd_sc_hd__mux4_1
X_16474_ _09522_ _09564_ vssd1 vssd1 vccd1 vccd1 _09565_ sky130_fd_sc_hd__xnor2_1
X_10898_ net6926 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13686_ _06813_ _06698_ _06856_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__or3_1
X_18213_ _09809_ _02431_ _01844_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__o21ai_1
X_15425_ _08507_ _08518_ _08519_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__a21boi_2
X_19193_ net5212 _03182_ _03184_ _03176_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__o211a_1
X_12637_ _05811_ _05815_ _05797_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18144_ _02371_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__clkbuf_1
X_15356_ _08181_ _08446_ _08450_ vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__and3_1
X_12568_ net21 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14307_ _07471_ _07477_ _07469_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__o21a_1
X_11519_ net4176 net4324 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__or2_1
X_18075_ _02309_ _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15287_ net4461 _08117_ _08136_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12499_ net4128 _05043_ net4 vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold207 net5098 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 net4336 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ _09936_ _09938_ _10045_ vssd1 vssd1 vccd1 vccd1 _10047_ sky130_fd_sc_hd__and3_1
Xhold229 net8191 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _07395_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14169_ _07335_ _07338_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__nand2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ net3060 net5733 net2874 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _02004_ _02065_ _02073_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__o21ai_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17859_ _01981_ _01995_ _01993_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_191_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20870_ _02515_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ net3402 net7558 net3086 vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7802 net4482 vssd1 vssd1 vccd1 vccd1 net8329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7813 rbzero.texu_hot\[0\] vssd1 vssd1 vccd1 vccd1 net8340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7824 net4629 vssd1 vssd1 vccd1 vccd1 net8351 sky130_fd_sc_hd__dlygate4sd3_1
X_21422_ clknet_leaf_41_i_clk net2062 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7835 net7763 vssd1 vssd1 vccd1 vccd1 net8362 sky130_fd_sc_hd__clkbuf_2
Xhold7846 rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 net8373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7868 net4495 vssd1 vssd1 vccd1 vccd1 net8395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21353_ clknet_leaf_12_i_clk net5139 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20304_ _03813_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__buf_4
Xhold730 net6477 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21284_ clknet_leaf_23_i_clk net5507 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold741 _00989_ vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 _03439_ vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
X_20235_ _02866_ _03710_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__or2_1
Xhold763 _03148_ vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 net6304 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _00991_ vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 net6310 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ net3882 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2120 rbzero.tex_b0\[61\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2131 net7064 vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2142 _01327_ vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2153 net7126 vssd1 vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2164 net7185 vssd1 vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20097_ net4748 _03662_ net617 _03688_ _03689_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a221o_1
Xhold1430 _01311_ vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2175 _01461_ vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _04388_ vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2186 _03587_ vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2197 _01368_ vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1452 net5763 vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1463 _01305_ vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1474 _04339_ vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 net7162 vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 net7110 vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ net4057 _04665_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nand2_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ net2783 net6478 _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ clknet_leaf_81_i_clk _00486_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20359__115 clknet_1_0__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__inv_2
XFILLER_0_184_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ net2008 net6466 _04182_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__mux2_1
X_13540_ _06709_ _06710_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13471_ _06505_ _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10683_ net6488 net2450 _04149_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12422_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _05258_ vssd1 vssd1 vccd1 vccd1 _05607_
+ sky130_fd_sc_hd__mux2_1
X_15210_ _08181_ _08298_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__o21ai_2
X_16190_ _09156_ _09273_ _09282_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _04909_ _05535_ _05538_ _05017_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15141_ net5768 net3419 _08196_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__buf_4
X_15072_ _08166_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__buf_4
X_12284_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04916_ vssd1 vssd1 vccd1 vccd1 _05470_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18900_ net3056 net5476 _03014_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
X_14023_ _07193_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__clkbuf_4
X_11235_ net6870 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
X_19880_ net3343 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
X_18831_ _02969_ _02973_ net3910 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__and3_1
X_11166_ net6462 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18762_ _02865_ net4560 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__or2_1
X_15974_ _09067_ _09068_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__nand2_1
X_11097_ net5675 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
X_17713_ _01949_ _01951_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14925_ net4651 _08050_ _08052_ net3669 net4758 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__o221a_1
X_18693_ net4560 net3619 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__or2_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 _03686_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _01882_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__nor2_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _08011_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _06955_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__xnor2_1
X_17575_ _10102_ _10103_ _01695_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__or3_1
X_14787_ _07843_ _07950_ _07941_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__a21oi_1
X_11999_ _04658_ _05183_ net4177 _04460_ _04600_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__o2111a_1
X_19314_ net1677 _03251_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__or2_1
X_16526_ _09505_ _09506_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _06906_ _06907_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20570__305 clknet_1_1__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__inv_2
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19245_ net5077 _03201_ _03214_ _03206_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__o211a_1
X_16457_ net3724 _09413_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__nand2_1
X_13669_ _06816_ _06817_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7109 _02721_ vssd1 vssd1 vccd1 vccd1 net7636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15408_ _08389_ _08417_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19176_ net5005 _03168_ _03174_ _03160_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__o211a_1
X_16388_ _08542_ _09115_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__nor2_1
Xhold6408 rbzero.tex_g0\[20\] vssd1 vssd1 vccd1 vccd1 net6935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6419 net2082 vssd1 vssd1 vccd1 vccd1 net6946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18127_ _02356_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__clkbuf_1
X_15339_ _08430_ _08433_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__nand2_1
Xhold5707 rbzero.tex_g0\[38\] vssd1 vssd1 vccd1 vccd1 net6234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5718 net1192 vssd1 vssd1 vccd1 vccd1 net6245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5729 rbzero.spi_registers.new_texadd\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net6256
+ sky130_fd_sc_hd__dlygate4sd3_1
X_18058_ _02279_ _02293_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17009_ _08226_ _09345_ vssd1 vssd1 vccd1 vccd1 _10030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20020_ net3461 _03607_ net4492 _03628_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_193_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19759__40 clknet_1_0__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
X_21971_ net413 net3001 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer11 _06944_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 _06945_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20922_ clknet_leaf_70_i_clk _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer33 _07091_ vssd1 vssd1 vccd1 vccd1 net3498 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer44 _06815_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_6
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer55 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19774__54 clknet_1_0__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
X_20853_ net4202 _04001_ _04002_ _09084_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a22o_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20784_ net1038 net5581 vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7610 rbzero.traced_texa\[-5\] vssd1 vssd1 vccd1 vccd1 net8137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7621 rbzero.row_render.texu\[0\] vssd1 vssd1 vccd1 vccd1 net8148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7632 rbzero.spi_registers.vshift\[0\] vssd1 vssd1 vccd1 vccd1 net8159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7643 rbzero.map_overlay.i_otherx\[3\] vssd1 vssd1 vccd1 vccd1 net8170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7654 _03933_ vssd1 vssd1 vccd1 vccd1 net8181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21405_ clknet_leaf_35_i_clk net4962 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6920 net2804 vssd1 vssd1 vccd1 vccd1 net7447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7665 rbzero.debug_overlay.playerX\[-1\] vssd1 vssd1 vccd1 vccd1 net8192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6931 rbzero.tex_b0\[27\] vssd1 vssd1 vccd1 vccd1 net7458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7676 rbzero.traced_texa\[-2\] vssd1 vssd1 vccd1 vccd1 net8203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6942 net2610 vssd1 vssd1 vccd1 vccd1 net7469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7687 net3457 vssd1 vssd1 vccd1 vccd1 net8214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6953 rbzero.pov.ready_buffer\[38\] vssd1 vssd1 vccd1 vccd1 net7480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7698 net3445 vssd1 vssd1 vccd1 vccd1 net8225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6964 rbzero.tex_g1\[12\] vssd1 vssd1 vccd1 vccd1 net7491 sky130_fd_sc_hd__dlygate4sd3_1
X_21336_ clknet_leaf_6_i_clk net5286 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6975 net3220 vssd1 vssd1 vccd1 vccd1 net7502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6986 rbzero.tex_g1\[13\] vssd1 vssd1 vccd1 vccd1 net7513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6997 net889 vssd1 vssd1 vccd1 vccd1 net7524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21267_ clknet_leaf_123_i_clk net2184 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold560 net5435 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
X_20684__5 clknet_1_0__leaf__03506_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
Xhold571 net6110 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net6251 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
Xhold582 net5477 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 net8137 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_1
X_20218_ _04459_ net3539 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__or2_1
X_21198_ clknet_leaf_127_i_clk net1104 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ net4446 _03711_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__or2_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ net2185 net4049 vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__xnor2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1260 _01265_ vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 net6658 vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ net7813 _07876_ _07879_ net8354 vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__a31o_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 _03599_ vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net3990 _05109_ _05110_ net3389 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a22o_1
Xhold1293 net6805 vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ _08783_ _08784_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__xnor2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _07800_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__nand2_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ net4177 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__clkbuf_4
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _08103_ _10378_ vssd1 vssd1 vccd1 vccd1 _10379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10804_ net6643 net7153 _04216_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__mux2_1
X_11784_ _04972_ _04973_ _04921_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__mux2_1
X_14572_ _07489_ _07327_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16311_ _09292_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13523_ _06683_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__nor2_8
X_17291_ _10308_ _10309_ vssd1 vssd1 vccd1 vccd1 _10310_ sky130_fd_sc_hd__nand2_1
X_10735_ _04030_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19030_ net3878 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
X_20678__23 clknet_1_0__leaf__03872_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XFILLER_0_153_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ net4640 _08115_ _09333_ _09334_ _01633_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__o221a_1
X_10666_ net6840 net2625 _04138_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13454_ _06394_ _06528_ _06609_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ _05465_ _05585_ _05589_ _04967_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a211o_1
X_16173_ _09264_ _09265_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__nor2_1
X_13385_ _06547_ _06552_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__o21ai_2
X_10597_ net7103 net6983 _04105_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15124_ _08156_ _08218_ _08148_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__o21a_1
X_12336_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _05369_ vssd1 vssd1 vccd1 vccd1 _05522_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20413__164 clknet_1_1__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__inv_2
XFILLER_0_142_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12267_ _05203_ _05450_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__o21ba_1
X_19932_ net6201 net3121 _03572_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__mux2_1
X_15055_ _06374_ _06375_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11218_ net6802 net6030 _04434_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
X_14006_ _07151_ _07128_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__a21o_1
XFILLER_0_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19863_ net3186 net3056 _03539_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__mux2_1
X_12198_ _05276_ _05382_ _05384_ _04928_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ net2988 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
X_18814_ net1547 net3851 net4814 _02958_ net3909 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__o311a_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18745_ _02856_ net3678 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or2_1
X_15957_ _08486_ _08520_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14908_ net4293 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__o21a_1
X_18676_ _02809_ _02810_ net3619 _02789_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__o2bb2a_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _08855_ _08892_ _08980_ _08982_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__o22ai_4
X_17627_ _01865_ _01866_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__nor2_1
X_14839_ net8362 _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17558_ _01796_ _01797_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _08543_ _09345_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17489_ _01730_ net4651 _10260_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19228_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6205 _03034_ vssd1 vssd1 vccd1 vccd1 net6732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6216 rbzero.pov.spi_buffer\[47\] vssd1 vssd1 vccd1 vccd1 net6743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6227 net1991 vssd1 vssd1 vccd1 vccd1 net6754 sky130_fd_sc_hd__dlygate4sd3_1
X_19159_ net5416 _03144_ _03163_ _03160_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__o211a_1
Xhold6238 rbzero.tex_b1\[34\] vssd1 vssd1 vccd1 vccd1 net6765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5504 _04437_ vssd1 vssd1 vccd1 vccd1 net6031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6249 net1920 vssd1 vssd1 vccd1 vccd1 net6776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5515 _04017_ vssd1 vssd1 vccd1 vccd1 net6042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5526 _04382_ vssd1 vssd1 vccd1 vccd1 net6053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22170_ clknet_leaf_87_i_clk net4950 vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5537 rbzero.spi_registers.got_new_mapd vssd1 vssd1 vccd1 vccd1 net6064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4803 net833 vssd1 vssd1 vccd1 vccd1 net5330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5548 rbzero.spi_registers.new_texadd\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net6075
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4814 _01607_ vssd1 vssd1 vccd1 vccd1 net5341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5559 net767 vssd1 vssd1 vccd1 vccd1 net6086 sky130_fd_sc_hd__dlygate4sd3_1
X_21121_ clknet_leaf_107_i_clk net4871 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4825 net978 vssd1 vssd1 vccd1 vccd1 net5352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4836 rbzero.spi_registers.texadd0\[6\] vssd1 vssd1 vccd1 vccd1 net5363 sky130_fd_sc_hd__dlygate4sd3_1
X_20388__141 clknet_1_1__leaf__03844_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__inv_2
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_124_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold4847 net981 vssd1 vssd1 vccd1 vccd1 net5374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4858 _01602_ vssd1 vssd1 vccd1 vccd1 net5385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21052_ clknet_leaf_74_i_clk _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4869 net995 vssd1 vssd1 vccd1 vccd1 net5396 sky130_fd_sc_hd__dlygate4sd3_1
X_20003_ _03609_ net5836 vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ net396 net2571 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20905_ clknet_leaf_65_i_clk _00392_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ net327 net3109 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20836_ _03320_ clknet_1_0__leaf__05688_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__and2_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20767_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10520_ net2797 net7457 _04064_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20698_ _03879_ _03880_ _03876_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7440 rbzero.wall_tracer.trackDistY\[5\] vssd1 vssd1 vccd1 vccd1 net7967 sky130_fd_sc_hd__dlygate4sd3_1
X_10451_ net3067 net49 _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7451 net4668 vssd1 vssd1 vccd1 vccd1 net7978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7462 rbzero.wall_tracer.trackDistY\[3\] vssd1 vssd1 vccd1 vccd1 net7989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7473 _00512_ vssd1 vssd1 vccd1 vccd1 net8000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7484 net4263 vssd1 vssd1 vccd1 vccd1 net8011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7495 _00509_ vssd1 vssd1 vccd1 vccd1 net8022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6750 net2435 vssd1 vssd1 vccd1 vccd1 net7277 sky130_fd_sc_hd__dlygate4sd3_1
X_13170_ rbzero.wall_tracer.rcp_sel\[0\] _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__and2_1
Xhold6761 _04108_ vssd1 vssd1 vccd1 vccd1 net7288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6772 net2155 vssd1 vssd1 vccd1 vccd1 net7299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12121_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _04951_ vssd1 vssd1 vccd1 vccd1 _05309_
+ sky130_fd_sc_hd__mux2_1
Xhold6783 net1682 vssd1 vssd1 vccd1 vccd1 net7310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6794 rbzero.tex_b1\[22\] vssd1 vssd1 vccd1 vccd1 net7321 sky130_fd_sc_hd__dlygate4sd3_1
X_21319_ clknet_leaf_14_i_clk net5446 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12052_ _04938_ _05240_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold390 net4882 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net5576 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
X_16860_ _09882_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15811_ _08318_ _08905_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ _09817_ _09819_ _09820_ vssd1 vssd1 vccd1 vccd1 _09821_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_204_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18530_ _02702_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__xnor2_1
X_15742_ _08226_ _08474_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__nor2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12954_ net3999 _06039_ _06035_ _06048_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__and4_1
XFILLER_0_198_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1090 net5582 vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _02617_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02640_
+ sky130_fd_sc_hd__nand2_1
X_11905_ _04465_ net3919 _05071_ net4108 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__or4_2
X_15673_ _08661_ _08473_ _08494_ _08185_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__or4b_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ net5974 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__inv_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ _10343_ _10338_ vssd1 vssd1 vccd1 vccd1 _10430_ sky130_fd_sc_hd__or2b_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14624_ _07441_ _07445_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__and3_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11836_ net4321 _04848_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__nor2_1
X_18392_ net4603 rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _02576_
+ sky130_fd_sc_hd__nand2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19753__35 clknet_1_0__leaf__03507_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _10218_ _10231_ vssd1 vssd1 vccd1 vccd1 _10362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14555_ _07723_ _07725_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__or2b_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11767_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _04933_ vssd1 vssd1 vccd1 vccd1 _04957_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13506_ _06647_ _06653_ _06557_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__mux2_1
X_17274_ _10190_ _08614_ _09062_ _08383_ vssd1 vssd1 vccd1 vccd1 _10293_ sky130_fd_sc_hd__o22a_1
X_10718_ net5632 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__clkbuf_1
X_14486_ _07306_ _07197_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11698_ net3423 net3365 net3014 vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nand3_1
X_19013_ net3396 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16225_ _09218_ _09317_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13437_ _06401_ _06403_ _06549_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ net6735 net2094 _04127_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer2 _07028_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16156_ _08204_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__buf_2
X_13368_ _06399_ _06466_ _06469_ _06477_ _06511_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_i_clk clknet_4_9__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15107_ _07947_ net8397 _08113_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__mux2_1
X_12319_ _04915_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or2_1
X_16087_ _09180_ _09035_ _08128_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__a21o_2
X_13299_ _06365_ _06405_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__xnor2_1
Xhold3409 _02981_ vssd1 vssd1 vccd1 vccd1 net3936 sky130_fd_sc_hd__dlygate4sd3_1
X_15038_ _08124_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__buf_4
X_19915_ net3138 net7453 _03561_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__mux2_1
Xhold2708 _01117_ vssd1 vssd1 vccd1 vccd1 net3235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2719 net7531 vssd1 vssd1 vccd1 vccd1 net3246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_i_clk clknet_4_11__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19846_ net2771 net6231 _03528_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19777_ clknet_1_1__leaf__03506_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__buf_1
X_16989_ _09788_ net8375 net8383 _10010_ vssd1 vssd1 vccd1 vccd1 _10011_ sky130_fd_sc_hd__a31o_1
X_18728_ _02856_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02879_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18659_ net4709 rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02815_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21670_ clknet_leaf_125_i_clk net2314 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6002 _02502_ vssd1 vssd1 vccd1 vccd1 net6529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6013 net1713 vssd1 vssd1 vccd1 vccd1 net6540 sky130_fd_sc_hd__dlygate4sd3_1
X_20483_ clknet_1_1__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__buf_1
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6024 rbzero.spi_registers.new_texadd\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net6551
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6035 net1665 vssd1 vssd1 vccd1 vccd1 net6562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6046 rbzero.spi_registers.new_mapd\[15\] vssd1 vssd1 vccd1 vccd1 net6573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5301 _01175_ vssd1 vssd1 vccd1 vccd1 net5828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5312 net3349 vssd1 vssd1 vccd1 vccd1 net5839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6057 rbzero.spi_registers.new_texadd\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net6584
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6068 net1806 vssd1 vssd1 vccd1 vccd1 net6595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5323 _03626_ vssd1 vssd1 vccd1 vccd1 net5850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6079 rbzero.tex_r1\[7\] vssd1 vssd1 vccd1 vccd1 net6606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5334 net3316 vssd1 vssd1 vccd1 vccd1 net5861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4600 net753 vssd1 vssd1 vccd1 vccd1 net5127 sky130_fd_sc_hd__dlygate4sd3_1
X_22153_ clknet_leaf_54_i_clk _01640_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5356 _02580_ vssd1 vssd1 vccd1 vccd1 net5883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4611 _00840_ vssd1 vssd1 vccd1 vccd1 net5138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4622 net764 vssd1 vssd1 vccd1 vccd1 net5149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5367 rbzero.spi_registers.spi_cmd\[3\] vssd1 vssd1 vccd1 vccd1 net5894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4633 rbzero.spi_registers.texadd2\[2\] vssd1 vssd1 vccd1 vccd1 net5160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5378 _01171_ vssd1 vssd1 vccd1 vccd1 net5905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21104_ clknet_leaf_1_i_clk net1449 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4644 net813 vssd1 vssd1 vccd1 vccd1 net5171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5389 _04686_ vssd1 vssd1 vccd1 vccd1 net5916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4655 _00847_ vssd1 vssd1 vccd1 vccd1 net5182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3910 _01193_ vssd1 vssd1 vccd1 vccd1 net4437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22084_ net526 net2042 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
Xhold3921 _01207_ vssd1 vssd1 vccd1 vccd1 net4448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4666 net750 vssd1 vssd1 vccd1 vccd1 net5193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4677 gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 net5204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3932 net3574 vssd1 vssd1 vccd1 vccd1 net4459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3943 net8390 vssd1 vssd1 vccd1 vccd1 net4470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4688 rbzero.spi_registers.texadd2\[5\] vssd1 vssd1 vccd1 vccd1 net5215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3954 net3599 vssd1 vssd1 vccd1 vccd1 net4481 sky130_fd_sc_hd__buf_1
Xhold4699 net821 vssd1 vssd1 vccd1 vccd1 net5226 sky130_fd_sc_hd__dlygate4sd3_1
X_21035_ clknet_leaf_34_i_clk net3650 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3965 _03630_ vssd1 vssd1 vccd1 vccd1 net4492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3976 _01222_ vssd1 vssd1 vccd1 vccd1 net4503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3987 _03726_ vssd1 vssd1 vccd1 vccd1 net4514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3998 net7953 vssd1 vssd1 vccd1 vccd1 net4525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21937_ net379 net2640 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _05848_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21868_ net310 net2493 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11621_ _04757_ _04760_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a21o_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20819_ _09727_ net8200 _03983_ _03689_ net5480 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__a32o_1
X_21799_ net241 net1829 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ _07510_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__inv_2
X_11552_ net4431 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net5677 net3240 _04053_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ _06699_ _07305_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__or2_1
X_11483_ net4095 net3326 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7270 net4412 vssd1 vssd1 vccd1 vccd1 net7797 sky130_fd_sc_hd__dlygate4sd3_1
X_16010_ net7778 vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__buf_1
XFILLER_0_123_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7281 rbzero.wall_tracer.stepDistX\[7\] vssd1 vssd1 vccd1 vccd1 net7808 sky130_fd_sc_hd__dlygate4sd3_1
X_13222_ _06382_ _06383_ _06355_ _06366_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6580 net2527 vssd1 vssd1 vccd1 vccd1 net7107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6591 rbzero.tex_b0\[14\] vssd1 vssd1 vccd1 vccd1 net7118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13153_ _06278_ _06291_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ net4140 _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nand2_1
X_13084_ _06254_ _06255_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__or2_1
X_17961_ _02196_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__xnor2_1
Xhold5890 net1489 vssd1 vssd1 vccd1 vccd1 net6417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16912_ _08338_ _08374_ _08383_ _08142_ vssd1 vssd1 vccd1 vccd1 _09934_ sky130_fd_sc_hd__o22ai_1
X_12035_ _04967_ _05209_ _05214_ _04818_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__o311a_1
X_19700_ net6629 net3866 _03468_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17892_ _02031_ _02098_ _02129_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a21oi_1
X_16843_ net4665 net4471 vssd1 vssd1 vccd1 vccd1 _09867_ sky130_fd_sc_hd__or2_1
X_19631_ net6568 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__clkbuf_1
X_20525__265 clknet_1_1__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__inv_2
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ _04102_ net1778 vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16774_ net3945 net4353 vssd1 vssd1 vccd1 vccd1 _09805_ sky130_fd_sc_hd__nor2_1
X_13986_ _07153_ _07156_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18513_ _02687_ _02688_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__nand2_1
X_15725_ _08782_ _08785_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__xnor2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19493_ net3519 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__inv_2
X_12937_ net4420 _06062_ _06060_ net3983 _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a221o_1
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ net8109 _02537_ _02616_ net4793 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__o211ai_1
X_15656_ _08726_ _08750_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__xor2_4
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ _06043_ _06028_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14607_ _07609_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__xnor2_4
X_11819_ _04825_ _04996_ _05000_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__o31a_1
X_18375_ net3494 rbzero.wall_tracer.rayAddendX\[-2\] _02551_ vssd1 vssd1 vccd1 vccd1
+ _02560_ sky130_fd_sc_hd__o21a_1
X_15587_ _08266_ _08317_ _08679_ _08681_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__or4bb_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _05948_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17326_ _10337_ _10344_ vssd1 vssd1 vccd1 vccd1 _10345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ _07284_ _07457_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _10161_ _10177_ _10175_ vssd1 vssd1 vccd1 vccd1 _10276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14469_ _07634_ _07635_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__a21o_1
X_16208_ _09036_ _09177_ _09300_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__o21a_1
X_17188_ _10088_ _10089_ _10086_ vssd1 vssd1 vccd1 vccd1 _10208_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16139_ _08529_ _09062_ _09230_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3206 _02347_ vssd1 vssd1 vccd1 vccd1 net3733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3217 rbzero.spi_registers.spi_buffer\[11\] vssd1 vssd1 vccd1 vccd1 net3744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3228 net7956 vssd1 vssd1 vccd1 vccd1 net3755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3239 net3424 vssd1 vssd1 vccd1 vccd1 net3766 sky130_fd_sc_hd__clkbuf_2
Xhold2505 net4061 vssd1 vssd1 vccd1 vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 _00755_ vssd1 vssd1 vccd1 vccd1 net3043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2527 _01138_ vssd1 vssd1 vccd1 vccd1 net3054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2538 _01103_ vssd1 vssd1 vccd1 vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 _03040_ vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 rbzero.pov.spi_buffer\[15\] vssd1 vssd1 vccd1 vccd1 net3076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 net7225 vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1826 _01279_ vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
X_19829_ net6413 net1579 _03517_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__mux2_1
Xhold1837 net810 vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1848 _01565_ vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 _01524_ vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21722_ clknet_leaf_102_i_clk net4411 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21653_ clknet_leaf_121_i_clk net1112 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21584_ net218 net940 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5120 net2251 vssd1 vssd1 vccd1 vccd1 net5647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5131 _01632_ vssd1 vssd1 vccd1 vccd1 net5658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5142 rbzero.tex_b1\[48\] vssd1 vssd1 vccd1 vccd1 net5669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5153 rbzero.tex_b1\[2\] vssd1 vssd1 vccd1 vccd1 net5680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5164 rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 net5691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5175 net3105 vssd1 vssd1 vccd1 vccd1 net5702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4430 _00896_ vssd1 vssd1 vccd1 vccd1 net4957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5186 rbzero.tex_g0\[0\] vssd1 vssd1 vccd1 vccd1 net5713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4441 net640 vssd1 vssd1 vccd1 vccd1 net4968 sky130_fd_sc_hd__dlygate4sd3_1
X_22136_ clknet_leaf_85_i_clk net3629 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4452 rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 net4979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5197 net2969 vssd1 vssd1 vccd1 vccd1 net5724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4463 net716 vssd1 vssd1 vccd1 vccd1 net4990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4474 net729 vssd1 vssd1 vccd1 vccd1 net5001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3740 net1029 vssd1 vssd1 vccd1 vccd1 net4267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4485 rbzero.spi_registers.texadd2\[20\] vssd1 vssd1 vccd1 vccd1 net5012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22067_ net509 net1914 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold3751 net8127 vssd1 vssd1 vccd1 vccd1 net4278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4496 net749 vssd1 vssd1 vccd1 vccd1 net5023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3762 net778 vssd1 vssd1 vccd1 vccd1 net4289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3773 net8121 vssd1 vssd1 vccd1 vccd1 net4300 sky130_fd_sc_hd__dlygate4sd3_1
X_21018_ clknet_leaf_59_i_clk net4238 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3784 net3037 vssd1 vssd1 vccd1 vccd1 net4311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3795 net8149 vssd1 vssd1 vccd1 vccd1 net4322 sky130_fd_sc_hd__dlygate4sd3_1
X_13840_ _06768_ _06931_ _06795_ _06758_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__a22o_1
X_13771_ _06939_ _06927_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__and2b_1
X_10983_ net6633 net2116 _04309_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15510_ _08595_ _08603_ _08604_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__a21oi_2
X_12722_ _05899_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _09579_ _09580_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _08139_ _08535_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ _04020_ _04495_ _04494_ _04500_ net22 _05797_ vssd1 vssd1 vccd1 vccd1 _05832_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_194_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11604_ _04789_ _04792_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or3_2
X_18160_ _02385_ net4567 _02320_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ _08456_ _08459_ _08466_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__nand3_2
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ net16 _05747_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17111_ _10130_ _10131_ vssd1 vssd1 vccd1 vccd1 _10132_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_167_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14323_ _07419_ _07490_ _07493_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__o21a_4
X_18091_ net3700 _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__xnor2_1
X_11535_ _04720_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17042_ _10062_ _08413_ vssd1 vssd1 vccd1 vccd1 _10063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14254_ _07412_ _07423_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11466_ net3452 net3628 net2 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ net4917 net8051 _04491_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14185_ _07350_ _07351_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__and2_1
X_11397_ _04503_ _04587_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _06303_ _06304_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a21oi_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ net3267 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _02165_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and2_1
X_13067_ _06053_ _06054_ _06241_ _06242_ net5605 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a32o_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20449__196 clknet_1_0__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__inv_2
X_12018_ rbzero.tex_r1\[7\] rbzero.tex_r1\[6\] _04968_ vssd1 vssd1 vccd1 vccd1 _05207_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17875_ _01985_ _01986_ _02112_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19614_ net6285 net1396 _03430_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
X_16826_ net4500 net4789 vssd1 vssd1 vccd1 vccd1 _09852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16757_ net4667 net3822 vssd1 vssd1 vccd1 vccd1 _09790_ sky130_fd_sc_hd__or2_1
X_19545_ net1403 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
X_13969_ _07138_ _07139_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nor2_1
X_15708_ _08765_ _08796_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16688_ net8132 _09743_ _09744_ net4268 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
X_19476_ net2061 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15639_ _08243_ _08433_ _08732_ _08733_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__a31o_1
X_18427_ net4554 net3661 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _02541_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ _10327_ _09170_ _10193_ _10197_ vssd1 vssd1 vccd1 vccd1 _10328_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18289_ net6365 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20320_ net6679 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold901 _00928_ vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 net5707 vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 net6465 vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_20251_ _05730_ _05044_ net3996 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__or3b_1
Xhold934 _01258_ vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 _03063_ vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 net6433 vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _03377_ vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3003 net4829 vssd1 vssd1 vccd1 vccd1 net3530 sky130_fd_sc_hd__dlygate4sd3_1
X_20182_ _03728_ net4003 vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2_1
Xhold978 net6147 vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3014 _01233_ vssd1 vssd1 vccd1 vccd1 net3541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _00581_ vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3025 rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1 net3552 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3036 _03094_ vssd1 vssd1 vccd1 vccd1 net3563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2302 net7559 vssd1 vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3047 net7880 vssd1 vssd1 vccd1 vccd1 net3574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3058 _00743_ vssd1 vssd1 vccd1 vccd1 net3585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2313 _00692_ vssd1 vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 net7235 vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3069 net1541 vssd1 vssd1 vccd1 vccd1 net3596 sky130_fd_sc_hd__buf_2
XFILLER_0_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2335 _01144_ vssd1 vssd1 vccd1 vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1601 net6879 vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2346 _02991_ vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2357 net5587 vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 _01012_ vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1623 net6957 vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2368 net7374 vssd1 vssd1 vccd1 vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2379 rbzero.tex_g1\[63\] vssd1 vssd1 vccd1 vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 net7020 vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1645 _01035_ vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
X_20662__8 clknet_1_1__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1656 net6793 vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1667 net5711 vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1678 _02487_ vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__clkbuf_4
Xhold1689 _01309_ vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21705_ clknet_leaf_118_i_clk net4750 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21636_ clknet_leaf_125_i_clk net3127 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21567_ net201 net1775 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ rbzero.spi_registers.texadd3\[12\] rbzero.spi_registers.texadd1\[12\] rbzero.spi_registers.texadd0\[12\]
+ rbzero.spi_registers.texadd2\[12\] _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04512_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21498_ clknet_leaf_3_i_clk net1572 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11251_ net6969 net2164 _04445_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11182_ net7248 net7059 _04412_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4260 net3515 vssd1 vssd1 vccd1 vccd1 net4787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4271 _02861_ vssd1 vssd1 vccd1 vccd1 net4798 sky130_fd_sc_hd__dlygate4sd3_1
X_22119_ clknet_leaf_57_i_clk net5254 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
Xhold4282 net8063 vssd1 vssd1 vccd1 vccd1 net4809 sky130_fd_sc_hd__dlygate4sd3_1
X_15990_ net7768 net5887 _08111_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__mux2_1
Xhold4293 _02644_ vssd1 vssd1 vccd1 vccd1 net4820 sky130_fd_sc_hd__buf_1
Xhold3570 _03119_ vssd1 vssd1 vccd1 vccd1 net4097 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3581 _05082_ vssd1 vssd1 vccd1 vccd1 net4108 sky130_fd_sc_hd__clkbuf_2
X_14941_ _04489_ _08066_ vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__nor2_2
Xhold3592 _00479_ vssd1 vssd1 vccd1 vccd1 net4119 sky130_fd_sc_hd__dlygate4sd3_1
X_17660_ _01898_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__nand2_1
Xhold2880 net8171 vssd1 vssd1 vccd1 vccd1 net3407 sky130_fd_sc_hd__buf_1
X_14872_ _08024_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__inv_2
Xhold2891 _09095_ vssd1 vssd1 vccd1 vccd1 net3418 sky130_fd_sc_hd__dlygate4sd3_1
X_16611_ _09633_ _09700_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__xnor2_1
X_13823_ _06949_ _06950_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__nand2_1
X_17591_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16542_ _09630_ _09631_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__nand2_1
X_19330_ net5013 _03235_ _03263_ _03259_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__o211a_1
X_13754_ _06703_ _06695_ _06923_ _06924_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_70_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ net6705 net6197 _04298_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19261_ net6422 _03217_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__or2_1
X_12705_ net4066 _05852_ _05865_ net71 _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a221o_1
X_16473_ _09562_ _09563_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__and2b_1
X_20637__366 clknet_1_0__leaf__03868_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__inv_2
X_13685_ _06715_ _06695_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10897_ net6924 net2589 _04265_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__mux2_1
X_18212_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15424_ _08483_ _08487_ _08506_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__or3_4
XFILLER_0_156_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19192_ net6315 _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__or2_1
X_12636_ _05812_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18143_ _02370_ net3768 _02320_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ net3574 _08133_ _08441_ _08449_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__a22o_4
X_12567_ net17 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__buf_2
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ _07472_ _07475_ _07476_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_151_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ net4095 net1817 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__xor2_1
X_18074_ _02258_ _02308_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15286_ _07968_ net3453 _08379_ _08380_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__a22o_2
X_12498_ net4127 vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__clkbuf_2
Xhold208 net6124 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _09936_ _09938_ _10045_ vssd1 vssd1 vccd1 vccd1 _10046_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold219 net6692 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ _07401_ _07407_ _07399_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__o21a_1
X_11449_ rbzero.spi_registers.texadd1\[0\] _04548_ _04640_ vssd1 vssd1 vccd1 vccd1
+ _04641_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14168_ _07335_ _07338_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__or2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nor2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__inv_2
X_18976_ net3039 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _02085_ _02087_ _02163_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__o21a_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20382__136 clknet_1_0__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__inv_2
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17858_ _02094_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__xor2_1
X_16809_ _09818_ _09084_ vssd1 vssd1 vccd1 vccd1 _09837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17789_ _01794_ _09664_ _01905_ _02027_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19528_ net3334 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19459_ net2223 _03335_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7803 rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 net8330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7814 net4558 vssd1 vssd1 vccd1 vccd1 net8341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_146_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7825 rbzero.texu_hot\[4\] vssd1 vssd1 vccd1 vccd1 net8352 sky130_fd_sc_hd__dlygate4sd3_1
X_21421_ clknet_leaf_41_i_clk net2443 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7847 net4372 vssd1 vssd1 vccd1 vccd1 net8374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21352_ clknet_leaf_47_i_clk net5075 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20303_ net6311 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21283_ clknet_leaf_24_i_clk net4433 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold720 net6262 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 net6479 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 net6505 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20234_ net7508 _03706_ net4710 _03765_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold753 _00974_ vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 net4355 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold775 _03431_ vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 net6455 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _01263_ vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
X_20165_ _03728_ net7624 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__or2_1
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2110 _01491_ vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2121 net2360 vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2132 _01575_ vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2143 net7253 vssd1 vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ _04458_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__buf_4
Xhold2154 _01040_ vssd1 vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 _04258_ vssd1 vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1420 _03016_ vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2176 net5683 vssd1 vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 net6927 vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1442 _01085_ vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2187 _01149_ vssd1 vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2198 net7088 vssd1 vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1453 net5765 vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 net6753 vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1475 _01322_ vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1486 _01576_ vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _04240_ vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _04193_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__clkbuf_4
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20998_ clknet_leaf_81_i_clk _00485_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10751_ net2519 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13470_ _06538_ _06551_ _06591_ _06640_ _06527_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10682_ net2620 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12421_ _04949_ _05603_ _05605_ _05465_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21619_ clknet_leaf_128_i_clk net737 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15140_ net3339 net8413 vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__nand2_1
X_12352_ _05035_ _05285_ _05536_ _05537_ net3781 vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ net7708 vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__clkbuf_8
X_15071_ _08118_ _08164_ _08165_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _04913_ vssd1 vssd1 vccd1 vccd1 _05469_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _07191_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nand2_2
X_11234_ net6868 net2911 _04434_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__mux2_1
X_18830_ net2198 _02947_ net3909 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a21o_1
X_11165_ net6460 net1982 _04401_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__mux2_1
Xhold4090 _03665_ vssd1 vssd1 vccd1 vccd1 net4617 sky130_fd_sc_hd__dlygate4sd3_1
X_15973_ _08618_ _09066_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__or2_1
X_11096_ net5586 net5673 _04364_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__mux2_1
X_18761_ net8242 _02905_ net4857 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__nand3_1
XFILLER_0_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17712_ _01949_ _01951_ _08103_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__o21ai_1
X_14924_ net8009 _08047_ _04482_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__o21a_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18692_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__inv_2
Xhold80 net4953 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold91 net4749 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _01759_ _01770_ _01768_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a21oi_1
X_14855_ net4459 _08010_ _07976_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__mux2_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13806_ _06956_ _06957_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__nand2_1
X_17574_ _10105_ _01695_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__nand2b_2
X_14786_ _07877_ _07878_ _07841_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__o21ai_1
X_11998_ _05183_ _05050_ net5948 _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16525_ _09479_ _09480_ _09482_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__a21bo_1
X_19313_ net5300 _03250_ _03254_ _03246_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__o211a_1
X_13737_ _06906_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10949_ net6711 net2265 _04287_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ net8041 _06123_ _09413_ _09546_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__or4_4
X_19244_ net1552 _03203_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__or2_1
X_13668_ net541 vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15407_ _08500_ _08501_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__xor2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ _05797_ net22 vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19175_ net6263 _03170_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or2_1
X_16387_ _09357_ _09358_ _09356_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__a21o_1
X_13599_ _06673_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__or2_1
Xhold6409 net2265 vssd1 vssd1 vccd1 vccd1 net6936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _02355_ net3847 _02320_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ net4168 _08137_ net8400 vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__o21a_4
XFILLER_0_152_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5708 net1139 vssd1 vssd1 vccd1 vccd1 net6235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5719 rbzero.pov.spi_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net6246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _02283_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__xnor2_1
X_15269_ _04511_ _06020_ _08114_ _08363_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__o211a_1
X_17008_ _09133_ net4914 _10028_ vssd1 vssd1 vccd1 vccd1 _10029_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18959_ net3227 net5743 net2874 vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21970_ net412 net2822 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer12 _06898_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_1
X_20921_ clknet_leaf_71_i_clk _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer23 _06951_ vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer34 _06996_ vssd1 vssd1 vccd1 vccd1 net3503 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_179_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer45 net571 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer56 _06744_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20852_ net4206 _04001_ _04002_ _09089_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a22o_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20783_ _03878_ _03952_ _03953_ _03883_ net5622 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7600 _00503_ vssd1 vssd1 vccd1 vccd1 net8127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7611 net1120 vssd1 vssd1 vccd1 vccd1 net8138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7622 _00494_ vssd1 vssd1 vccd1 vccd1 net8149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7633 rbzero.map_overlay.i_otherx\[1\] vssd1 vssd1 vccd1 vccd1 net8160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7644 rbzero.pov.ready_buffer\[33\] vssd1 vssd1 vccd1 vccd1 net8171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6910 net3176 vssd1 vssd1 vccd1 vccd1 net7437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7655 _01611_ vssd1 vssd1 vccd1 vccd1 net8182 sky130_fd_sc_hd__dlygate4sd3_1
X_21404_ clknet_leaf_36_i_clk net3659 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6921 rbzero.pov.spi_buffer\[62\] vssd1 vssd1 vccd1 vccd1 net7448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7666 net2898 vssd1 vssd1 vccd1 vccd1 net8193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6932 net2962 vssd1 vssd1 vccd1 vccd1 net7459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6943 rbzero.pov.ready_buffer\[46\] vssd1 vssd1 vccd1 vccd1 net7470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7688 rbzero.debug_overlay.playerY\[-5\] vssd1 vssd1 vccd1 vccd1 net8215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6954 net3690 vssd1 vssd1 vccd1 vccd1 net7481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7699 rbzero.debug_overlay.playerX\[-8\] vssd1 vssd1 vccd1 vccd1 net8226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6965 net3152 vssd1 vssd1 vccd1 vccd1 net7492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21335_ clknet_leaf_6_i_clk net5322 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6976 rbzero.tex_b0\[47\] vssd1 vssd1 vccd1 vccd1 net7503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6987 net3249 vssd1 vssd1 vccd1 vccd1 net7514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6998 _03383_ vssd1 vssd1 vccd1 vccd1 net7525 sky130_fd_sc_hd__dlygate4sd3_1
X_21266_ clknet_leaf_123_i_clk net2057 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold550 _03136_ vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 net5437 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 net6112 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold583 net6200 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
X_20217_ net4528 net1862 _03709_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold594 net4237 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
X_21197_ clknet_leaf_126_i_clk net1620 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20365__120 clknet_1_0__leaf__03842_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__inv_2
X_20148_ net7093 _03707_ net4514 _03679_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20079_ net4327 _03485_ _03662_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__a211o_1
X_12970_ net4009 net5975 vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nand2_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 _03387_ vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__buf_2
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1261 net3226 vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _05079_ _05101_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_1
Xhold1272 _01302_ vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _01161_ vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 _01078_ vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _07805_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__xor2_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net4126 net4160 vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__nand2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ net6786 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _07072_ _07198_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__or2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _04837_ vssd1 vssd1 vccd1 vccd1 _04973_
+ sky130_fd_sc_hd__mux2_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16310_ _08417_ _09165_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13522_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__buf_2
X_17290_ _10204_ _10277_ _10307_ vssd1 vssd1 vccd1 vccd1 _10309_ sky130_fd_sc_hd__nand3_1
X_10734_ net1995 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16241_ net7779 _09332_ net3454 vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__a21o_1
X_13453_ _06564_ _06620_ _06623_ _06540_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__o211a_1
X_10665_ net2141 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _05517_ _05586_ _05588_ _05306_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__o211a_1
X_16172_ _08207_ _09262_ _09142_ _09140_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13384_ _06547_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__nand2_1
X_10596_ net2915 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ net3419 _08196_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__xnor2_2
X_12335_ _05517_ _05518_ _05520_ _05233_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19931_ net2543 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
X_15054_ rbzero.wall_tracer.visualWallDist\[-8\] _08117_ _08148_ vssd1 vssd1 vccd1
+ vccd1 _08149_ sky130_fd_sc_hd__a21o_1
X_12266_ net3781 _05015_ _05285_ _05452_ net42 vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__o311a_1
X_14005_ _07163_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__xnor2_1
X_11217_ net2480 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__clkbuf_1
X_19862_ net736 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__clkbuf_4
X_12197_ _04910_ _05383_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18813_ net3084 _02955_ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a21oi_1
X_11148_ net7405 net6995 _04390_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__mux2_1
X_18744_ _02879_ _02885_ _02892_ _04478_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a31o_1
X_15956_ _09015_ _09050_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__xnor2_1
X_11079_ net3092 net6948 _04353_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
X_14907_ net4500 _08034_ _08036_ net3768 net4683 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__o221a_1
X_15887_ _08855_ _08981_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__xor2_2
X_18675_ _02828_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__or2_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17626_ _01750_ _01751_ _01749_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14838_ _07952_ _07993_ _07994_ _07995_ _07913_ net7785 vssd1 vssd1 vccd1 vccd1 _07996_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17557_ _01796_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14769_ _07882_ _07886_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _09521_ _09500_ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17488_ _06058_ _10387_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19227_ _08092_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__clkbuf_4
X_16439_ _09524_ _09529_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6206 net1619 vssd1 vssd1 vccd1 vccd1 net6733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6217 net1885 vssd1 vssd1 vccd1 vccd1 net6744 sky130_fd_sc_hd__dlygate4sd3_1
X_19158_ net3002 _03146_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or2_1
Xhold6228 rbzero.tex_g0\[53\] vssd1 vssd1 vccd1 vccd1 net6755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6239 net1955 vssd1 vssd1 vccd1 vccd1 net6766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5505 net634 vssd1 vssd1 vccd1 vccd1 net6032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18109_ _02339_ _02340_ _09820_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5516 gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 net6043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5527 net661 vssd1 vssd1 vccd1 vccd1 net6054 sky130_fd_sc_hd__dlygate4sd3_1
X_19089_ net4095 net3970 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__nand2_1
Xhold5538 net886 vssd1 vssd1 vccd1 vccd1 net6065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5549 net2414 vssd1 vssd1 vccd1 vccd1 net6076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4804 rbzero.spi_registers.texadd1\[1\] vssd1 vssd1 vccd1 vccd1 net5331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4815 net916 vssd1 vssd1 vccd1 vccd1 net5342 sky130_fd_sc_hd__dlygate4sd3_1
X_21120_ clknet_leaf_92_i_clk net3892 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4826 _00810_ vssd1 vssd1 vccd1 vccd1 net5353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4837 net929 vssd1 vssd1 vccd1 vccd1 net5364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4848 rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 net5375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4859 net849 vssd1 vssd1 vccd1 vccd1 net5386 sky130_fd_sc_hd__dlygate4sd3_1
X_21051_ clknet_leaf_75_i_clk _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20002_ net5835 _08171_ _03615_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21953_ net395 net2473 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ clknet_leaf_65_i_clk _00391_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21884_ net326 net3248 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20835_ _09413_ net5923 net3872 _01633_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__o31a_1
XFILLER_0_210_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20766_ _03936_ _03937_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20697_ _03876_ _03879_ _03880_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7430 rbzero.wall_tracer.trackDistX\[-8\] vssd1 vssd1 vccd1 vccd1 net7957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__clkbuf_4
Xhold7441 net3802 vssd1 vssd1 vccd1 vccd1 net7968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7452 rbzero.wall_tracer.trackDistX\[5\] vssd1 vssd1 vccd1 vccd1 net7979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7463 net3810 vssd1 vssd1 vccd1 vccd1 net7990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7474 net4221 vssd1 vssd1 vccd1 vccd1 net8001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6740 rbzero.tex_r1\[47\] vssd1 vssd1 vccd1 vccd1 net7267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7485 net8007 vssd1 vssd1 vccd1 vccd1 net8012 sky130_fd_sc_hd__buf_2
XFILLER_0_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6751 rbzero.tex_g0\[45\] vssd1 vssd1 vccd1 vccd1 net7278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7496 net4257 vssd1 vssd1 vccd1 vccd1 net8023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6762 net2787 vssd1 vssd1 vccd1 vccd1 net7289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6773 rbzero.tex_b0\[23\] vssd1 vssd1 vccd1 vccd1 net7300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12120_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _04951_ vssd1 vssd1 vccd1 vccd1 _05308_
+ sky130_fd_sc_hd__mux2_1
Xhold6784 rbzero.pov.mosi vssd1 vssd1 vccd1 vccd1 net7311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6795 net3092 vssd1 vssd1 vccd1 vccd1 net7322 sky130_fd_sc_hd__dlygate4sd3_1
X_21318_ clknet_leaf_21_i_clk net5438 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12051_ rbzero.tex_r1\[27\] rbzero.tex_r1\[26\] _05239_ vssd1 vssd1 vccd1 vccd1 _05240_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold380 net5164 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
X_21249_ clknet_leaf_2_i_clk net3740 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold391 net4884 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net2285 net5574 _04320_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__mux2_1
X_15810_ _08458_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16790_ _09809_ _09091_ vssd1 vssd1 vccd1 vccd1 _09820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15741_ _08834_ _08835_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__xnor2_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ net3960 _06062_ _06061_ _06043_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__and4_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6__f_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold1080 _01593_ vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 net6730 vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _05079_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__nor2_2
XFILLER_0_198_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15672_ _08206_ _08457_ _08733_ _08732_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__or4b_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ net5874 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__clkbuf_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ net4048 vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__buf_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _10326_ _10328_ _10330_ vssd1 vssd1 vccd1 vccd1 _10429_ sky130_fd_sc_hd__o21ai_2
X_14623_ _07439_ _07792_ _07791_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__nand3_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ net87 _04977_ _04848_ net4321 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__or4b_1
X_18391_ net4603 rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _02575_
+ sky130_fd_sc_hd__or2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _10218_ _10231_ vssd1 vssd1 vccd1 vccd1 _10361_ sky130_fd_sc_hd__and2_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _07668_ _07724_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__xor2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _04949_ _04952_ _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _06540_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__buf_1
X_17273_ _10167_ _10168_ _10166_ vssd1 vssd1 vccd1 vccd1 _10292_ sky130_fd_sc_hd__a21bo_1
X_10717_ net5630 net5601 _04171_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14485_ _07610_ _07651_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__xor2_2
XFILLER_0_183_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ net3388 _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16224_ _09315_ _09316_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19012_ _02972_ net3395 _02969_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__or3b_1
X_13436_ _06596_ _06603_ _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__a21oi_2
X_10648_ net2756 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer3 net7786 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_1
X_16155_ _09155_ _09160_ _09247_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13367_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__clkbuf_4
X_10579_ net1529 net6928 _04097_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15106_ _06002_ _06324_ net4180 vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12318_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _04912_ vssd1 vssd1 vccd1 vccd1 _05504_
+ sky130_fd_sc_hd__mux2_1
X_16086_ net3551 _08491_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ _06467_ _06433_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__and3_2
X_15037_ _08127_ _08131_ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__nor2_1
X_19914_ net2070 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
X_12249_ rbzero.tex_g1\[55\] rbzero.tex_g1\[54\] _04837_ vssd1 vssd1 vccd1 vccd1 _05436_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03514_ _03514_ vssd1 vssd1 vccd1 vccd1 clknet_0__03514_ sky130_fd_sc_hd__clkbuf_16
Xhold2709 rbzero.pov.spi_buffer\[69\] vssd1 vssd1 vccd1 vccd1 net3236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19845_ net2870 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16988_ _08103_ _10009_ vssd1 vssd1 vccd1 vccd1 _10010_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18727_ net5777 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
X_15939_ _08010_ _08017_ _08439_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__or3_1
XFILLER_0_211_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20502__244 clknet_1_1__leaf__03855_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__inv_2
X_18658_ net4709 rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02814_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ _01847_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__or2b_1
XFILLER_0_176_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18589_ net7633 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6003 net1603 vssd1 vssd1 vccd1 vccd1 net6530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6014 rbzero.spi_registers.new_texadd\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 net6541
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6025 net1555 vssd1 vssd1 vccd1 vccd1 net6552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6036 _03478_ vssd1 vssd1 vccd1 vccd1 net6563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6047 net1637 vssd1 vssd1 vccd1 vccd1 net6574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5302 net2899 vssd1 vssd1 vccd1 vccd1 net5829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6058 net1677 vssd1 vssd1 vccd1 vccd1 net6585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6069 rbzero.spi_registers.new_mapd\[12\] vssd1 vssd1 vccd1 vccd1 net6596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5324 _03627_ vssd1 vssd1 vccd1 vccd1 net5851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5335 rbzero.spi_registers.sclk_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net5862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4601 rbzero.spi_registers.texadd2\[0\] vssd1 vssd1 vccd1 vccd1 net5128 sky130_fd_sc_hd__dlygate4sd3_1
X_22152_ clknet_leaf_53_i_clk _01639_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5346 _02639_ vssd1 vssd1 vccd1 vccd1 net5873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5357 net3828 vssd1 vssd1 vccd1 vccd1 net5884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4612 net788 vssd1 vssd1 vccd1 vccd1 net5139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4623 _00800_ vssd1 vssd1 vccd1 vccd1 net5150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5368 net4814 vssd1 vssd1 vccd1 vccd1 net5895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5379 rbzero.pov.ready_buffer\[69\] vssd1 vssd1 vccd1 vccd1 net5906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4634 net793 vssd1 vssd1 vccd1 vccd1 net5161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3900 net7847 vssd1 vssd1 vccd1 vccd1 net4427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21103_ clknet_leaf_0_i_clk net1604 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4645 rbzero.spi_registers.texadd3\[17\] vssd1 vssd1 vccd1 vccd1 net5172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4656 net829 vssd1 vssd1 vccd1 vccd1 net5183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3911 net665 vssd1 vssd1 vccd1 vccd1 net4438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22083_ net525 net2792 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3922 net776 vssd1 vssd1 vccd1 vccd1 net4449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4667 _00857_ vssd1 vssd1 vccd1 vccd1 net5194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3933 net8348 vssd1 vssd1 vccd1 vccd1 net4460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4678 net3516 vssd1 vssd1 vccd1 vccd1 net5205 sky130_fd_sc_hd__buf_2
XFILLER_0_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3944 net3573 vssd1 vssd1 vccd1 vccd1 net4471 sky130_fd_sc_hd__clkbuf_2
Xhold4689 net858 vssd1 vssd1 vccd1 vccd1 net5216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3955 net8328 vssd1 vssd1 vccd1 vccd1 net4482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21034_ clknet_leaf_34_i_clk net3783 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3966 _01174_ vssd1 vssd1 vccd1 vccd1 net4493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3977 net629 vssd1 vssd1 vccd1 vccd1 net4504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3988 _01206_ vssd1 vssd1 vccd1 vccd1 net4515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3999 net1663 vssd1 vssd1 vccd1 vccd1 net4526 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21936_ net378 net1259 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20477__221 clknet_1_1__leaf__03853_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__inv_2
XFILLER_0_171_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21867_ net309 net1874 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ _04805_ _04808_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a21oi_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818_ _03981_ _03980_ _03979_ _03976_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21798_ net240 net2580 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ net4354 _04464_ _04465_ net4369 _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20749_ net822 net4980 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ net5790 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__clkbuf_1
X_14270_ _07437_ _07440_ net8355 vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a21o_1
X_11482_ net4160 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7260 net530 vssd1 vssd1 vccd1 vccd1 net7787 sky130_fd_sc_hd__clkbuf_2
X_13221_ _06390_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__xor2_4
Xhold7271 net3507 vssd1 vssd1 vccd1 vccd1 net7798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7282 net4519 vssd1 vssd1 vccd1 vccd1 net7809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6570 net2601 vssd1 vssd1 vccd1 vccd1 net7097 sky130_fd_sc_hd__dlygate4sd3_1
X_13152_ _06265_ _06015_ _06322_ _04491_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a211oi_2
Xhold6581 _04428_ vssd1 vssd1 vccd1 vccd1 net7108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6592 net2170 vssd1 vssd1 vccd1 vccd1 net7119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _04707_ _05200_ _05291_ _04706_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5880 net1456 vssd1 vssd1 vccd1 vccd1 net6407 sky130_fd_sc_hd__dlygate4sd3_1
X_17960_ _10190_ _09612_ _02102_ _02100_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__o31a_1
X_13083_ _06254_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__nand2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5891 rbzero.spi_registers.new_texadd\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net6418
+ sky130_fd_sc_hd__dlygate4sd3_1
X_16911_ _09655_ _09662_ _09932_ vssd1 vssd1 vccd1 vccd1 _09933_ sky130_fd_sc_hd__a21bo_1
X_12034_ _05213_ _05217_ _05219_ _05222_ _04825_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a221o_1
X_17891_ _02111_ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19630_ net6566 net2953 _03430_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
X_16842_ _09866_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__clkbuf_1
X_19561_ _03363_ net1777 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16773_ net3805 _09798_ _09797_ vssd1 vssd1 vccd1 vccd1 _09804_ sky130_fd_sc_hd__o21a_1
X_13985_ _07154_ _07155_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ _02627_ net4603 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__nand2_1
X_15724_ _08814_ _08817_ _08818_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__a21boi_1
X_12936_ net4369 _06068_ _06105_ _06106_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__a221o_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ net1562 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18443_ _09747_ net4792 _02623_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _08745_ _08749_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__and2_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ net3848 vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__inv_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _05002_ _05004_ _05007_ _04988_ net85 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_123_i_clk clknet_4_4__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14606_ _07652_ _07693_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__nor2_2
X_15586_ _08244_ _08252_ _08254_ _08680_ _08246_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__a32o_1
X_18374_ _09738_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__buf_4
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ net4416 net3761 vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__or2_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _10338_ _10343_ vssd1 vssd1 vccd1 vccd1 _10344_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14537_ _07672_ _07707_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__xnor2_1
X_11749_ _04936_ _04937_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17256_ _10273_ _10274_ vssd1 vssd1 vccd1 vccd1 _10275_ sky130_fd_sc_hd__nor2_1
X_14468_ _07636_ _07637_ _07638_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16207_ _09171_ _09178_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__nand2_1
X_13419_ _06435_ _06545_ _06536_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__or3b_4
X_17187_ _10183_ _10206_ vssd1 vssd1 vccd1 vccd1 _10207_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14399_ _07568_ _07569_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16138_ _08529_ _09062_ _09230_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _08417_ _08411_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__nor2_1
Xhold3207 rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 net3734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3218 net1392 vssd1 vssd1 vccd1 vccd1 net3745 sky130_fd_sc_hd__buf_2
Xhold3229 net4915 vssd1 vssd1 vccd1 vccd1 net3756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2506 _03113_ vssd1 vssd1 vccd1 vccd1 net3033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2517 net7527 vssd1 vssd1 vccd1 vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2528 rbzero.pov.spi_buffer\[21\] vssd1 vssd1 vccd1 vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2539 rbzero.tex_r1\[63\] vssd1 vssd1 vccd1 vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 _00689_ vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 net5660 vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
X_19828_ net3046 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1827 net7012 vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1838 _03015_ vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 rbzero.tex_g1\[44\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21721_ clknet_leaf_100_i_clk net3689 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21652_ clknet_leaf_118_i_clk net2544 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21583_ net217 net2574 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5110 rbzero.tex_r1\[32\] vssd1 vssd1 vccd1 vccd1 net5637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5121 rbzero.tex_b1\[29\] vssd1 vssd1 vccd1 vccd1 net5648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5132 rbzero.tex_r1\[15\] vssd1 vssd1 vccd1 vccd1 net5659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5143 _04336_ vssd1 vssd1 vccd1 vccd1 net5670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5154 _04386_ vssd1 vssd1 vccd1 vccd1 net5681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4420 gpout2.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5165 net2494 vssd1 vssd1 vccd1 vccd1 net5692 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_203_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4431 net613 vssd1 vssd1 vccd1 vccd1 net4958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5176 rbzero.pov.ready_buffer\[45\] vssd1 vssd1 vccd1 vccd1 net5703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22135_ clknet_leaf_85_i_clk net4087 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5187 net2697 vssd1 vssd1 vccd1 vccd1 net5714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4442 _01600_ vssd1 vssd1 vccd1 vccd1 net4969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4453 net650 vssd1 vssd1 vccd1 vccd1 net4980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5198 rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 net5725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4464 rbzero.spi_registers.texadd3\[3\] vssd1 vssd1 vccd1 vccd1 net4991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3730 net8022 vssd1 vssd1 vccd1 vccd1 net4257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4475 _00868_ vssd1 vssd1 vccd1 vccd1 net5002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3741 rbzero.wall_tracer.visualWallDist\[-6\] vssd1 vssd1 vccd1 vccd1 net4268
+ sky130_fd_sc_hd__buf_2
XFILLER_0_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22066_ net508 net935 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold4486 net687 vssd1 vssd1 vccd1 vccd1 net5013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3752 net961 vssd1 vssd1 vccd1 vccd1 net4279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4497 rbzero.spi_registers.texadd3\[12\] vssd1 vssd1 vccd1 vccd1 net5024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3763 rbzero.wall_tracer.visualWallDist\[8\] vssd1 vssd1 vccd1 vccd1 net4290 sky130_fd_sc_hd__buf_1
Xhold3774 net949 vssd1 vssd1 vccd1 vccd1 net4301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3785 net8159 vssd1 vssd1 vccd1 vccd1 net4312 sky130_fd_sc_hd__dlymetal6s2s_1
X_21017_ clknet_leaf_57_i_clk net4270 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3796 net673 vssd1 vssd1 vccd1 vccd1 net4323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13770_ _06920_ _06913_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__xnor2_1
X_10982_ net1974 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_40_i_clk clknet_4_9__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12721_ reg_gpout\[4\] clknet_1_1__leaf__05898_ net45 vssd1 vssd1 vccd1 vccd1 _05899_
+ sky130_fd_sc_hd__mux2_2
X_21919_ net361 net1598 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15440_ _08534_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__buf_2
Xclkbuf_2_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_12652_ net4133 net4089 _05802_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ net950 net1217 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15371_ _08461_ net8033 _08464_ _08465_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_26_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_55_i_clk clknet_4_14__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17110_ _10006_ _10008_ _10004_ vssd1 vssd1 vccd1 vccd1 _10131_ sky130_fd_sc_hd__o21ai_2
X_14322_ _07491_ _07492_ _07418_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18090_ _02322_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__nand2_1
X_11534_ _04682_ net4306 net4315 _04684_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ net4918 vssd1 vssd1 vccd1 vccd1 _10062_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14253_ _07415_ _07422_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__nor2_1
X_11465_ net4083 net4862 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20531__270 clknet_1_1__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__inv_2
Xhold7090 net3675 vssd1 vssd1 vccd1 vccd1 net7617 sky130_fd_sc_hd__dlygate4sd3_1
X_13204_ _06269_ _06300_ _06373_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ _07237_ _07354_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__xnor2_1
X_11396_ _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__or2_1
X_13135_ _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__clkbuf_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ net7175 net5849 _03058_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _02172_ _02179_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__xor2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13066_ _06240_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__clkbuf_4
X_12017_ _04832_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__buf_4
X_17874_ _01760_ _08612_ _01982_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19613_ net1302 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__clkbuf_1
X_16825_ net4500 net4789 vssd1 vssd1 vccd1 vccd1 _09851_ sky130_fd_sc_hd__nor2_1
X_19544_ net5562 net1493 _03388_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__mux2_1
Xmax_cap1 _06465_ vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__clkbuf_1
X_16756_ net4667 net3822 vssd1 vssd1 vccd1 vccd1 _09789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13968_ _06911_ _07095_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__nor2_1
X_15707_ _08798_ _08801_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__xnor2_1
X_12919_ _04731_ net3893 _06048_ net4357 _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__o221a_1
X_19475_ net2205 net6007 _03345_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16687_ net8126 _09743_ _09744_ net4277 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a22o_1
X_13899_ _07032_ _07067_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18426_ net4554 net3661 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15638_ _08166_ _08185_ _08463_ _08572_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _02542_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__or2b_1
XFILLER_0_185_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _08186_ _08433_ _08662_ _08663_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20614__345 clknet_1_1__leaf__03866_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__inv_2
X_17308_ _08326_ vssd1 vssd1 vccd1 vccd1 _10327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18288_ net6363 net2953 _02477_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17239_ _09788_ _10139_ _10140_ _10258_ vssd1 vssd1 vccd1 vccd1 _10259_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold902 net6410 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _01518_ vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20250_ _04500_ net3642 _03789_ net5208 _08093_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__o311a_1
Xhold924 net6467 vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 net6483 vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _00710_ vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _03444_ vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
X_20181_ net7746 net3080 _03723_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__mux2_1
Xhold968 _00927_ vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3004 net7919 vssd1 vssd1 vccd1 vccd1 net3531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3015 net7848 vssd1 vssd1 vccd1 vccd1 net3542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold979 net6149 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3026 _04685_ vssd1 vssd1 vccd1 vccd1 net3553 sky130_fd_sc_hd__buf_1
Xhold3037 _00735_ vssd1 vssd1 vccd1 vccd1 net3564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3048 net7739 vssd1 vssd1 vccd1 vccd1 net3575 sky130_fd_sc_hd__clkbuf_4
Xhold2303 net7466 vssd1 vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 net7146 vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3059 net8349 vssd1 vssd1 vccd1 vccd1 net3586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2325 _04040_ vssd1 vssd1 vccd1 vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2336 net2926 vssd1 vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1602 net6881 vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2347 _03047_ vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__clkbuf_4
Xhold2358 _01291_ vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 net6859 vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 _04455_ vssd1 vssd1 vccd1 vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _01282_ vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 _03010_ vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 net6984 vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1657 _00754_ vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 _00697_ vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 net7304 vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21704_ clknet_leaf_118_i_clk net4904 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21635_ clknet_leaf_125_i_clk net3097 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21566_ net200 net2746 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20589__322 clknet_1_1__leaf__03864_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__inv_2
XFILLER_0_160_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21497_ clknet_leaf_1_i_clk net1905 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11250_ net2316 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11181_ net7027 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4250 net4660 vssd1 vssd1 vccd1 vccd1 net4777 sky130_fd_sc_hd__clkbuf_2
X_22118_ clknet_leaf_57_i_clk net5406 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4261 net7928 vssd1 vssd1 vccd1 vccd1 net4788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4272 _02863_ vssd1 vssd1 vccd1 vccd1 net4799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4283 net3760 vssd1 vssd1 vccd1 vccd1 net4810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4294 _02645_ vssd1 vssd1 vccd1 vccd1 net4821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3560 _01622_ vssd1 vssd1 vccd1 vccd1 net4087 sky130_fd_sc_hd__dlygate4sd3_1
X_22049_ net491 net1960 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold3571 _03803_ vssd1 vssd1 vccd1 vccd1 net4098 sky130_fd_sc_hd__clkdlybuf4s25_1
X_14940_ net3871 net3976 net3774 _04485_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__or4_1
Xhold3582 _00477_ vssd1 vssd1 vccd1 vccd1 net4109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3593 net4131 vssd1 vssd1 vccd1 vccd1 net4120 sky130_fd_sc_hd__clkbuf_1
Xhold2870 _03077_ vssd1 vssd1 vccd1 vccd1 net3397 sky130_fd_sc_hd__buf_2
Xhold2881 net4627 vssd1 vssd1 vccd1 vccd1 net3408 sky130_fd_sc_hd__dlygate4sd3_1
X_14871_ net7794 _07973_ _08023_ _08020_ _07869_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__a221oi_4
Xhold2892 net5903 vssd1 vssd1 vccd1 vccd1 net3419 sky130_fd_sc_hd__buf_2
XFILLER_0_173_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16610_ _09698_ _09699_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _06882_ _06908_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__xnor2_2
X_17590_ _01780_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16541_ _09519_ _09598_ _09629_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__nand3_1
X_13753_ _06706_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ net2492 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12704_ net49 _05864_ _05881_ _05862_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__a211o_1
XFILLER_0_211_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19260_ net8135 _03216_ net987 _03219_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__o211a_1
X_16472_ _09559_ _09561_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__nand2_1
X_13684_ _06715_ _06698_ _06714_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ net3203 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18211_ _02422_ _02423_ _02420_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15423_ _08512_ _08517_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__xor2_2
X_12635_ net24 vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19191_ _03169_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15354_ _08008_ _08009_ _08447_ _08448_ _08114_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__a311o_1
X_18142_ _09809_ _02369_ _09855_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__o21ai_1
X_12566_ _05744_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14305_ _07242_ _07198_ _07473_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__or3_1
X_11517_ _04691_ _04694_ _04700_ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a31o_1
X_15285_ _04510_ _06025_ _08112_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__o21a_1
X_18073_ _02258_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ net4103 net4024 net5965 net6044 net4 net7 vssd1 vssd1 vccd1 vccd1 _05679_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17024_ _10043_ _10044_ vssd1 vssd1 vccd1 vccd1 _10045_ sky130_fd_sc_hd__xnor2_1
Xhold209 net6126 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ _07402_ _07405_ _07406_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _04554_ _04555_ rbzero.spi_registers.texadd3\[0\] vssd1 vssd1 vccd1 vccd1
+ _04640_ sky130_fd_sc_hd__or3b_1
XFILLER_0_180_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _07336_ _07337_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ _04503_ _04569_ _04570_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _07210_ _07218_ _07216_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__o21a_1
X_18975_ net3283 net6061 net2874 vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17926_ _02080_ _02088_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__or2b_1
X_13049_ _06180_ _06181_ _06224_ _06171_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o31a_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17857_ _02012_ _02034_ _02010_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a21oi_1
X_16808_ net4632 _09835_ vssd1 vssd1 vccd1 vccd1 _09836_ sky130_fd_sc_hd__xnor2_1
X_17788_ _01903_ _01904_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19527_ net3816 net3333 net3086 vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__mux2_1
X_16739_ _09750_ _09751_ _09774_ _09770_ vssd1 vssd1 vccd1 vccd1 _09775_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19458_ net5464 _03334_ _03341_ _03339_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18409_ _02570_ _02571_ net3661 _02549_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19389_ net5248 _03268_ _03297_ _03288_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7804 net4497 vssd1 vssd1 vccd1 vccd1 net8331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21420_ clknet_leaf_41_i_clk net1726 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7815 rbzero.wall_tracer.stepDistY\[9\] vssd1 vssd1 vccd1 vccd1 net8342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7826 net4768 vssd1 vssd1 vccd1 vccd1 net8353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7837 _08134_ vssd1 vssd1 vccd1 vccd1 net8364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7848 _09885_ vssd1 vssd1 vccd1 vccd1 net8375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21351_ clknet_leaf_47_i_clk net5298 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20302_ net6309 net2953 _03814_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold710 _01568_ vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21282_ clknet_leaf_24_i_clk net4422 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold721 _03434_ vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 _01423_ vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold743 net6507 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
X_20233_ net4709 _03710_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 net6290 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 net6286 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 _00966_ vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 net6457 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 net6346 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
X_20164_ rbzero.debug_overlay.facingY\[-5\] net1915 _03723_ vssd1 vssd1 vccd1 vccd1
+ _03737_ sky130_fd_sc_hd__mux2_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2100 _01495_ vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2111 net7292 vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2122 _04392_ vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 rbzero.tex_r0\[7\] vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2144 net7255 vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ net4748 _03682_ _03687_ _03659_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__a22o_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _01446_ vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2155 net2844 vssd1 vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2166 _01395_ vssd1 vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1421 _00667_ vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2177 net5685 vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 net6929 vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2188 net7313 vssd1 vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1443 net7002 vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2199 _04420_ vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1454 _00717_ vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1465 _04078_ vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1476 net3401 vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 net6883 vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1498 _01412_ vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20997_ clknet_4_15__leaf_i_clk _00484_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ net6466 net7275 _04182_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ net6989 net6488 _04149_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12420_ _04943_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21618_ clknet_leaf_98_i_clk net3157 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ net4080 _05021_ _05372_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_129_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21549_ net183 net1723 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ net7678 vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__buf_6
X_15070_ net4390 _08123_ _08148_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__a21o_2
X_12282_ _05466_ _05467_ _05206_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _07148_ _07190_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__nand2_1
X_11233_ net2171 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ net3118 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4080 net8342 vssd1 vssd1 vccd1 vccd1 net4607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4091 _03666_ vssd1 vssd1 vccd1 vccd1 net4618 sky130_fd_sc_hd__dlygate4sd3_1
X_18760_ _02904_ _02905_ net4857 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a21o_1
X_15972_ _08618_ _09066_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__nand2_1
X_11095_ net1070 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17711_ _01723_ _01726_ _01841_ _01950_ _01840_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__o311a_4
X_20643__371 clknet_1_1__leaf__03869_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__inv_2
Xhold3390 net5945 vssd1 vssd1 vccd1 vccd1 net3917 sky130_fd_sc_hd__dlygate4sd3_1
X_14923_ net4610 _08050_ _08052_ net3811 net4738 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__o221a_1
X_18691_ net5856 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 net6392 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 net4947 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _01872_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__xnor2_1
Xhold92 net4959 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _08008_ _08009_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__nand2_2
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ _06961_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17573_ _01806_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__xnor2_1
X_14785_ _07905_ _07906_ _07843_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__a21o_1
X_11997_ net4095 _04462_ _05179_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor3_1
XFILLER_0_203_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19312_ net1456 _03251_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__or2_1
X_16524_ _09611_ _09613_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__xor2_1
X_10948_ net6109 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
X_13736_ _06823_ _06825_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19243_ net5029 _03201_ _03213_ _03206_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16455_ _08421_ _09544_ _09545_ _08442_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__a31o_2
X_10879_ net7186 net6756 _04253_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__mux2_1
X_13667_ _06836_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _08161_ _08418_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12618_ net23 vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__clkbuf_4
X_19174_ net5236 _03168_ _03173_ _03160_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__o211a_1
X_16386_ _09475_ _09476_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__and2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _06768_ _06720_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18125_ _09809_ _02354_ _09837_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__o21ai_1
X_15337_ _06119_ net8399 vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ net5965 vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5709 _04277_ vssd1 vssd1 vccd1 vccd1 net6236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_152_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18056_ _02288_ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _04597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15268_ net4181 _06361_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17007_ _08226_ _09225_ vssd1 vssd1 vccd1 vccd1 _10028_ sky130_fd_sc_hd__nor2_1
X_14219_ _07146_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15199_ _08290_ _08291_ _08293_ _06121_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__a22o_4
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18958_ net2873 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17909_ _01855_ _02045_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a21oi_2
X_18889_ net3063 net7045 _03003_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
X_20920_ clknet_leaf_73_i_clk _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer13 _06808_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
Xrebuffer24 _06878_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 _06526_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_1
XFILLER_0_156_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer46 net571 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_1
X_20851_ _09738_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__clkbuf_4
Xrebuffer57 _06960_ vssd1 vssd1 vccd1 vccd1 net3526 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20782_ _03948_ _03949_ _03950_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20471__216 clknet_1_1__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__inv_2
XFILLER_0_135_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7601 rbzero.wall_tracer.rayAddendY\[-5\] vssd1 vssd1 vccd1 vccd1 net8128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7612 _00505_ vssd1 vssd1 vccd1 vccd1 net8139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7623 rbzero.map_overlay.i_mapdy\[0\] vssd1 vssd1 vccd1 vccd1 net8150 sky130_fd_sc_hd__dlygate4sd3_1
X_21403_ clknet_leaf_41_i_clk net3654 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7634 rbzero.map_overlay.i_othery\[1\] vssd1 vssd1 vccd1 vccd1 net8161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6900 net2999 vssd1 vssd1 vccd1 vccd1 net7427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7645 _01197_ vssd1 vssd1 vccd1 vccd1 net8172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6911 rbzero.tex_r1\[27\] vssd1 vssd1 vccd1 vccd1 net7438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6922 net2712 vssd1 vssd1 vccd1 vccd1 net7449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7667 rbzero.spi_registers.got_new_texadd\[1\] vssd1 vssd1 vccd1 vccd1 net8194
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7678 _08042_ vssd1 vssd1 vccd1 vccd1 net8205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6933 rbzero.pov.ready_buffer\[41\] vssd1 vssd1 vccd1 vccd1 net7460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6944 net3252 vssd1 vssd1 vccd1 vccd1 net7471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7689 net4344 vssd1 vssd1 vccd1 vccd1 net8216 sky130_fd_sc_hd__clkdlybuf4s25_1
X_21334_ clknet_leaf_9_i_clk net4209 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6955 _03035_ vssd1 vssd1 vccd1 vccd1 net7482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6966 _04234_ vssd1 vssd1 vccd1 vccd1 net7493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6977 net3117 vssd1 vssd1 vccd1 vccd1 net7504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6988 rbzero.pov.spi_buffer\[31\] vssd1 vssd1 vccd1 vccd1 net7515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6999 net2954 vssd1 vssd1 vccd1 vccd1 net7526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21265_ clknet_leaf_122_i_clk net3034 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold540 net5443 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold551 net4307 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 net6151 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
X_20216_ net7419 _03706_ net4636 _03765_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__o211a_1
Xhold573 _01662_ vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _03577_ vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold595 net5451 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
X_21196_ clknet_leaf_125_i_clk net3364 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20147_ net4513 _03711_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or2_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _08258_ _03610_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nor2_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1240 net6676 vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 _03401_ vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1262 _03048_ vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ _05079_ _05085_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1273 net6531 vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1284 net6519 vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 net5595 vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__buf_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11851_ _04707_ net4155 _05039_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o22a_1
XFILLER_0_197_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10802_ net2515 net6784 _04216_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14570_ _07413_ _07391_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__nor2_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _04968_ vssd1 vssd1 vccd1 vccd1 _04972_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ net6227 net6796 _04097_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
X_13521_ _06436_ _06684_ _06686_ _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a31o_4
X_19780__59 clknet_1_0__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16240_ net7779 _09332_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__nor2_1
X_13452_ _06538_ _06621_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__or3b_1
X_10664_ net6860 net6840 _04138_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12403_ _04922_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16171_ _09261_ _09263_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ _06438_ _06447_ _06450_ _06441_ _06551_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_
+ sky130_fd_sc_hd__mux4_1
X_10595_ net7415 net7103 _04105_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _05276_ _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15122_ net3419 _08156_ vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19930_ net3052 net6201 _03572_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__mux2_1
X_15053_ _06118_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12265_ net4335 _05306_ _05451_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _07164_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__xnor2_1
X_11216_ net7297 net6802 _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_1
X_19861_ net6125 net3186 _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12196_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _04912_ vssd1 vssd1 vccd1 vccd1 _05383_
+ sky130_fd_sc_hd__mux2_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 o_gpout[4] sky130_fd_sc_hd__buf_1
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18812_ net3851 net4814 net1547 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__o21a_1
X_11147_ net6536 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _02879_ _02885_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a21oi_1
X_15955_ _09047_ _09049_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__xor2_1
X_11078_ net6701 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
X_14906_ net4280 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08048_ sky130_fd_sc_hd__o21a_1
X_18674_ net3575 _05164_ _02826_ _02827_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o22a_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _08808_ _08813_ _08853_ _08893_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__a31o_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__nand2_1
X_14837_ _07877_ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__inv_2
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17556_ _10327_ _09664_ _01664_ _01668_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__o31a_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ net7785 vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__clkbuf_4
X_16507_ _09477_ _09495_ _09493_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ _06887_ _06888_ _06889_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a21bo_1
X_17487_ net90 _01727_ _01728_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__or3_4
XFILLER_0_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14699_ net7833 _07848_ _07867_ _07869_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__a31o_2
X_19226_ net6474 _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__or2_1
X_16438_ _09527_ _09528_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6207 rbzero.tex_r0\[35\] vssd1 vssd1 vccd1 vccd1 net6734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19157_ net5157 _03144_ _03162_ _03160_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__o211a_1
X_16369_ _09323_ _09325_ _09449_ _09459_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__o31a_4
Xhold6218 rbzero.tex_b0\[58\] vssd1 vssd1 vccd1 vccd1 net6745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6229 net2052 vssd1 vssd1 vccd1 vccd1 net6756 sky130_fd_sc_hd__dlygate4sd3_1
X_18108_ net3731 _02338_ _09845_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__a21o_1
Xhold5506 rbzero.tex_g1\[8\] vssd1 vssd1 vccd1 vccd1 net6033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19088_ net7681 net5981 net4102 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__and3_1
Xhold5517 net3995 vssd1 vssd1 vccd1 vccd1 net6044 sky130_fd_sc_hd__buf_2
Xhold5528 rbzero.spi_registers.new_floor\[3\] vssd1 vssd1 vccd1 vccd1 net6055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5539 _03420_ vssd1 vssd1 vccd1 vccd1 net6066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4805 net868 vssd1 vssd1 vccd1 vccd1 net5332 sky130_fd_sc_hd__dlygate4sd3_1
X_18039_ _09181_ _09060_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__nor2_1
Xhold4816 rbzero.spi_registers.texadd2\[23\] vssd1 vssd1 vccd1 vccd1 net5343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4827 net979 vssd1 vssd1 vccd1 vccd1 net5354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4838 _00789_ vssd1 vssd1 vccd1 vccd1 net5365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4849 net884 vssd1 vssd1 vccd1 vccd1 net5376 sky130_fd_sc_hd__dlygate4sd3_1
X_21050_ clknet_leaf_65_i_clk _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20001_ net3536 _03607_ net5818 _03339_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21952_ net394 net2461 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ clknet_leaf_37_i_clk net5410 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21883_ net325 net3091 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20834_ _04474_ net4083 net3871 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20395__147 clknet_1_1__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__inv_2
X_20765_ _03931_ _03935_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20696_ net756 net4984 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7420 rbzero.wall_tracer.trackDistX\[-4\] vssd1 vssd1 vccd1 vccd1 net7947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7431 net4568 vssd1 vssd1 vccd1 vccd1 net7958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7442 rbzero.wall_tracer.trackDistX\[4\] vssd1 vssd1 vccd1 vccd1 net7969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7453 net4658 vssd1 vssd1 vccd1 vccd1 net7980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7464 rbzero.wall_tracer.trackDistY\[7\] vssd1 vssd1 vccd1 vccd1 net7991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6730 rbzero.tex_b0\[8\] vssd1 vssd1 vccd1 vccd1 net7257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7475 net8264 vssd1 vssd1 vccd1 vccd1 net8002 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6741 net2984 vssd1 vssd1 vccd1 vccd1 net7268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7486 _00513_ vssd1 vssd1 vccd1 vccd1 net8013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6752 net2589 vssd1 vssd1 vccd1 vccd1 net7279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6763 rbzero.tex_g0\[51\] vssd1 vssd1 vccd1 vccd1 net7290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6774 net2854 vssd1 vssd1 vccd1 vccd1 net7301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21317_ clknet_leaf_4_i_clk net5350 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6785 net1814 vssd1 vssd1 vccd1 vccd1 net7312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6796 rbzero.tex_r1\[9\] vssd1 vssd1 vccd1 vccd1 net7323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ _04835_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__buf_4
Xhold370 net4294 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
X_21248_ clknet_leaf_2_i_clk net3564 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold381 net5166 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net5655 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
Xhold392 net6057 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
X_21179_ clknet_leaf_99_i_clk net2366 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15740_ _08771_ _08770_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__and2b_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ net4034 net3893 _06039_ net3999 _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__o221a_1
Xhold1070 net6294 vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _06503_ vssd1 vssd1 vccd1 vccd1 net3638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 net6732 vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net4108 _05091_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__or2b_2
X_15671_ _08735_ _08738_ _08737_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__a21o_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ net3682 vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__inv_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17410_ _10393_ _10427_ vssd1 vssd1 vccd1 vccd1 _10428_ sky130_fd_sc_hd__xnor2_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _07439_ _07791_ _07792_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net4080 _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__xnor2_1
X_18390_ net4784 _02564_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__nand2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _10336_ _10359_ vssd1 vssd1 vccd1 vccd1 _10360_ sky130_fd_sc_hd__xnor2_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _04850_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ _07685_ _07684_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__and2b_1
XFILLER_0_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20454__200 clknet_1_1__leaf__03851_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__inv_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ net591 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__clkbuf_1
X_13504_ _06644_ _06674_ _06547_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17272_ _10287_ _10290_ vssd1 vssd1 vccd1 vccd1 _10291_ sky130_fd_sc_hd__xor2_1
X_14484_ _07608_ _07654_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__xnor2_2
X_11696_ net3365 net3014 net3423 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19011_ net3695 net1250 _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__nor3_1
X_16223_ _09219_ _09220_ _09314_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10647_ net7238 net6735 _04127_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_125_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer4 net7787 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_1
XFILLER_0_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ _09161_ _09154_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__or2b_1
X_13366_ _06503_ _06511_ _06515_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or3_1
X_10578_ net6556 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15105_ _08192_ net8425 _08195_ _08199_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__a2bb2o_4
X_12317_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _05249_ vssd1 vssd1 vccd1 vccd1 _05503_
+ sky130_fd_sc_hd__mux2_1
X_16085_ _09171_ _09178_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13297_ _06389_ _06401_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _05433_ _05434_ _04915_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__mux2_1
X_15036_ _08128_ net4918 vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__or2_2
X_19913_ net7178 net3138 _03561_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03513_ _03513_ vssd1 vssd1 vccd1 vccd1 clknet_0__03513_ sky130_fd_sc_hd__clkbuf_16
X_19844_ net7542 net2771 _03528_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
X_12179_ _04825_ _05354_ _05358_ _05366_ _04844_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16987_ _10006_ _10008_ vssd1 vssd1 vccd1 vccd1 _10009_ sky130_fd_sc_hd__xor2_4
XFILLER_0_208_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18726_ rbzero.wall_tracer.rayAddendY\[4\] _02877_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15938_ _08010_ net553 _08017_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18657_ net8025 _02803_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15869_ _08907_ _08942_ _08944_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17608_ net3875 net4624 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18588_ _02749_ net7631 net4648 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17539_ _01744_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20550_ clknet_1_0__leaf__03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__buf_1
XFILLER_0_11_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19209_ net6727 _03183_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__05847_ clknet_0__05847_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05847_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6004 rbzero.spi_registers.new_texadd\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net6531
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6015 net1668 vssd1 vssd1 vccd1 vccd1 net6542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6026 rbzero.tex_r1\[4\] vssd1 vssd1 vccd1 vccd1 net6553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6037 net1666 vssd1 vssd1 vccd1 vccd1 net6564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6048 _03419_ vssd1 vssd1 vccd1 vccd1 net6575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6059 rbzero.tex_g0\[62\] vssd1 vssd1 vccd1 vccd1 net6586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5314 _02903_ vssd1 vssd1 vccd1 vccd1 net5841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5325 _01173_ vssd1 vssd1 vccd1 vccd1 net5852 sky130_fd_sc_hd__dlygate4sd3_1
X_22151_ clknet_leaf_51_i_clk _01638_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5336 net3041 vssd1 vssd1 vccd1 vccd1 net5863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5347 net3813 vssd1 vssd1 vccd1 vccd1 net5874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4602 net721 vssd1 vssd1 vccd1 vccd1 net5129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5358 _00601_ vssd1 vssd1 vccd1 vccd1 net5885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4613 rbzero.spi_registers.texadd1\[5\] vssd1 vssd1 vccd1 vccd1 net5140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4624 net765 vssd1 vssd1 vccd1 vccd1 net5151 sky130_fd_sc_hd__dlygate4sd3_1
X_21102_ clknet_leaf_0_i_clk net1720 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5369 _03108_ vssd1 vssd1 vccd1 vccd1 net5896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4635 _00833_ vssd1 vssd1 vccd1 vccd1 net5162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22082_ net524 net2562 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold3901 net3542 vssd1 vssd1 vccd1 vccd1 net4428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4646 net808 vssd1 vssd1 vccd1 vccd1 net5173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3912 net8379 vssd1 vssd1 vccd1 vccd1 net4439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4657 rbzero.spi_registers.texadd0\[5\] vssd1 vssd1 vccd1 vccd1 net5184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4668 net751 vssd1 vssd1 vccd1 vccd1 net5195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3923 net7568 vssd1 vssd1 vccd1 vccd1 net4450 sky130_fd_sc_hd__clkbuf_4
Xhold3934 net3586 vssd1 vssd1 vccd1 vccd1 net4461 sky130_fd_sc_hd__buf_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21033_ clknet_leaf_55_i_clk net4252 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4679 _04501_ vssd1 vssd1 vccd1 vccd1 net5206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3956 net3600 vssd1 vssd1 vccd1 vccd1 net4483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3967 net3462 vssd1 vssd1 vccd1 vccd1 net4494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3978 net7930 vssd1 vssd1 vccd1 vccd1 net4505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3989 net780 vssd1 vssd1 vccd1 vccd1 net4516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21935_ net377 net2785 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ net308 net1132 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20817_ _03976_ _03979_ _03980_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__o211ai_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21797_ net239 net2538 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
X_11550_ net4420 _04460_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__xor2_1
X_20748_ _03878_ _03922_ _03923_ _03883_ net4972 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10501_ net3240 net5788 _04053_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ net4177 net4436 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _06382_ _06383_ _06365_ _06355_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__o2bb2a_4
Xhold7250 _06033_ vssd1 vssd1 vccd1 vccd1 net7777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7261 rbzero.wall_tracer.stepDistY\[1\] vssd1 vssd1 vccd1 vccd1 net7788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7272 net4751 vssd1 vssd1 vccd1 vccd1 net7799 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7283 _06493_ vssd1 vssd1 vccd1 vccd1 net7810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7294 net4777 vssd1 vssd1 vccd1 vccd1 net7821 sky130_fd_sc_hd__buf_1
Xhold6560 net2981 vssd1 vssd1 vccd1 vccd1 net7087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ net4280 _06265_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
Xhold6571 rbzero.tex_b1\[37\] vssd1 vssd1 vccd1 vccd1 net7098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6582 net2528 vssd1 vssd1 vccd1 vccd1 net7109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6593 rbzero.tex_r1\[62\] vssd1 vssd1 vccd1 vccd1 net7120 sky130_fd_sc_hd__dlygate4sd3_1
X_12102_ _05202_ _05290_ net7570 vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13082_ _06249_ _06252_ _06247_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a21oi_1
Xhold5870 net1320 vssd1 vssd1 vccd1 vccd1 net6397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5881 rbzero.spi_registers.new_texadd\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net6408
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5892 net1416 vssd1 vssd1 vccd1 vccd1 net6419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16910_ _09656_ _09661_ vssd1 vssd1 vccd1 vccd1 _09932_ sky130_fd_sc_hd__nand2_1
X_12033_ _04977_ _05221_ _04988_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__o21a_1
X_17890_ _02126_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _09865_ net3888 net4649 vssd1 vssd1 vccd1 vccd1 _09866_ sky130_fd_sc_hd__mux2_1
X_19560_ _03352_ net3376 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__nor2_1
X_16772_ _09803_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__clkbuf_1
X_13984_ _06576_ net3533 net571 _06693_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__o22a_1
X_18511_ _02627_ net4603 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__or2_1
X_15723_ _08815_ _08816_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ _04738_ net4034 net3965 _06108_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a221o_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ net2205 net6021 _03354_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18442_ net4791 _02619_ _02621_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__and3_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ _08745_ _08746_ _08748_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__nand3_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ net3893 _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _07695_ _07732_ _07774_ _07775_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__o31ai_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11817_ _05005_ _05006_ _04832_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__mux2_1
X_18373_ net5832 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__clkbuf_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15585_ _08277_ _08278_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12797_ _05964_ _05970_ _05972_ _05961_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _10341_ _10342_ vssd1 vssd1 vccd1 vccd1 _10343_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _07682_ _07681_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__and2b_1
X_11748_ _04832_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17255_ _10179_ _10271_ _10272_ vssd1 vssd1 vccd1 vccd1 _10274_ sky130_fd_sc_hd__and3_1
X_14467_ _07072_ _06754_ _07233_ _07280_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ net2910 _04856_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16206_ _09293_ _09298_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__xor2_2
XFILLER_0_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ _06540_ _06582_ _06587_ _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__a31o_4
X_17186_ _10204_ _10205_ vssd1 vssd1 vccd1 vccd1 _10206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14398_ _07562_ _07566_ _07567_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _08277_ _08614_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__or2_1
X_13349_ _06481_ _06398_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16068_ _09154_ _09161_ vssd1 vssd1 vccd1 vccd1 _09162_ sky130_fd_sc_hd__xnor2_1
Xhold3208 net6016 vssd1 vssd1 vccd1 vccd1 net3735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3219 _03091_ vssd1 vssd1 vccd1 vccd1 net3746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _08113_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__buf_4
Xhold2507 _00752_ vssd1 vssd1 vccd1 vccd1 net3034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2518 net2506 vssd1 vssd1 vccd1 vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2529 net2920 vssd1 vssd1 vccd1 vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1806 net7400 vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_19827_ net3045 net6413 _03517_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__mux2_1
Xhold1817 _01548_ vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 _04311_ vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 _00666_ vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20426__176 clknet_1_0__leaf__03847_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__inv_2
X_18709_ net4797 _02858_ _02860_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19689_ net1454 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21720_ clknet_leaf_109_i_clk net4449 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21651_ clknet_leaf_118_i_clk net3054 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21582_ net216 net2490 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20335__93 clknet_1_0__leaf__03514_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__inv_2
XFILLER_0_145_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5100 _04456_ vssd1 vssd1 vccd1 vccd1 net5627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5111 _04067_ vssd1 vssd1 vccd1 vccd1 net5638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5122 net2823 vssd1 vssd1 vccd1 vccd1 net5649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5133 _04085_ vssd1 vssd1 vccd1 vccd1 net5660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5144 net2623 vssd1 vssd1 vccd1 vccd1 net5671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5155 net2352 vssd1 vssd1 vccd1 vccd1 net5682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4410 _01661_ vssd1 vssd1 vccd1 vccd1 net4937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5166 _01616_ vssd1 vssd1 vccd1 vccd1 net5693 sky130_fd_sc_hd__dlygate4sd3_1
X_22134_ clknet_leaf_56_i_clk net5611 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold4421 net608 vssd1 vssd1 vccd1 vccd1 net4948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5177 net4616 vssd1 vssd1 vccd1 vccd1 net5704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4432 rbzero.color_floor\[1\] vssd1 vssd1 vccd1 vccd1 net4959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4443 net641 vssd1 vssd1 vccd1 vccd1 net4970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5188 _04317_ vssd1 vssd1 vccd1 vccd1 net5715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4454 net8198 vssd1 vssd1 vccd1 vccd1 net4981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5199 net2753 vssd1 vssd1 vccd1 vccd1 net5726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3720 rbzero.wall_tracer.visualWallDist\[5\] vssd1 vssd1 vccd1 vccd1 net4247 sky130_fd_sc_hd__buf_1
Xhold4465 net668 vssd1 vssd1 vccd1 vccd1 net4992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3731 net823 vssd1 vssd1 vccd1 vccd1 net4258 sky130_fd_sc_hd__dlygate4sd3_1
X_22065_ net507 net1841 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold4476 net730 vssd1 vssd1 vccd1 vccd1 net5003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3742 net8133 vssd1 vssd1 vccd1 vccd1 net4269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4487 _00851_ vssd1 vssd1 vccd1 vccd1 net5014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3753 rbzero.wall_tracer.visualWallDist\[-4\] vssd1 vssd1 vccd1 vccd1 net4280
+ sky130_fd_sc_hd__buf_2
Xhold4498 net717 vssd1 vssd1 vccd1 vccd1 net5025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3764 net8089 vssd1 vssd1 vccd1 vccd1 net4291 sky130_fd_sc_hd__dlygate4sd3_1
X_21016_ clknet_leaf_59_i_clk net4279 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3775 net8309 vssd1 vssd1 vccd1 vccd1 net4302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3786 _00897_ vssd1 vssd1 vccd1 vccd1 net4313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3797 net8163 vssd1 vssd1 vccd1 vccd1 net4324 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10981_ net6655 net6633 _04309_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ net4164 _05855_ _05861_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__o22a_2
X_21918_ net360 net2505 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12651_ net24 _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__or2_1
X_21849_ net291 net2868 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11602_ _04790_ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15370_ _08421_ _08424_ _08426_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__a21o_1
X_12582_ _05757_ _05761_ _05747_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14321_ _06924_ _06755_ _07303_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__or3_4
X_11533_ net4091 _04721_ _04722_ _04460_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_191_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ _09954_ _09962_ vssd1 vssd1 vccd1 vccd1 _10061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14252_ _07415_ _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__nand2_1
X_11464_ net3871 net3975 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7080 net3684 vssd1 vssd1 vccd1 vccd1 net7607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13203_ _06269_ _06300_ _06373_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nand3_1
Xhold7091 gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 net7618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14183_ _07341_ _07353_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__xor2_1
X_11395_ _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__nand2_1
X_20566__301 clknet_1_0__leaf__03862_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__inv_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6390 rbzero.tex_r0\[32\] vssd1 vssd1 vccd1 vccd1 net6917 sky130_fd_sc_hd__dlygate4sd3_1
X_13134_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__inv_2
X_18991_ net2864 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17942_ _02173_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__xor2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _06058_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__nor2_2
XFILLER_0_178_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12016_ rbzero.tex_r1\[5\] rbzero.tex_r1\[4\] _04838_ vssd1 vssd1 vccd1 vccd1 _05205_
+ sky130_fd_sc_hd__mux2_1
X_17873_ _02109_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19612_ net6305 net3897 _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__mux2_1
X_16824_ net4633 _09841_ _09842_ vssd1 vssd1 vccd1 vccd1 _09850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19543_ net1583 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16755_ net91 vssd1 vssd1 vccd1 vccd1 _09788_ sky130_fd_sc_hd__clkbuf_8
X_13967_ _06910_ _06865_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__and2b_1
X_15706_ _08692_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__nand2_1
X_19474_ net2442 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
X_12918_ net4384 net4044 vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__xnor2_1
X_16686_ net754 _09743_ _09744_ rbzero.wall_tracer.visualWallDist\[-8\] vssd1 vssd1
+ vccd1 vccd1 _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13898_ _07004_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__xnor2_1
X_18425_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15637_ _08185_ _08463_ _08572_ _08166_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__a22o_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12849_ _06022_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_158_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18356_ net4698 rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _02543_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15568_ _08630_ _08167_ _08464_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__and3b_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17307_ _10324_ _10325_ vssd1 vssd1 vccd1 vccd1 _10326_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14519_ _07627_ _07646_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__xnor2_1
X_18287_ net1509 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__clkbuf_1
X_15499_ _08586_ _08592_ _08593_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17238_ _08103_ _10257_ vssd1 vssd1 vccd1 vccd1 _10258_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold903 _03404_ vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ _10185_ _10188_ vssd1 vssd1 vccd1 vccd1 _10189_ sky130_fd_sc_hd__and2_1
Xhold914 net6377 vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold925 _01455_ vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold936 _03472_ vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 net6445 vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
X_20180_ net3929 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
Xhold958 _00978_ vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold969 net6421 vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3005 net7789 vssd1 vssd1 vccd1 vccd1 net3532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3016 net7586 vssd1 vssd1 vccd1 vccd1 net3543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3027 net6062 vssd1 vssd1 vccd1 vccd1 net3554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3038 net7737 vssd1 vssd1 vccd1 vccd1 net3565 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3049 _03773_ vssd1 vssd1 vccd1 vccd1 net3576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2304 _00702_ vssd1 vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2315 _04419_ vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 _01589_ vssd1 vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2337 _03064_ vssd1 vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1603 _01579_ vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 _03051_ vssd1 vssd1 vccd1 vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1614 _04145_ vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 rbzero.tex_g0\[56\] vssd1 vssd1 vccd1 vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1625 net7438 vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1636 _00662_ vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1647 _04077_ vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 net8157 vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1669 net7984 vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21703_ clknet_leaf_119_i_clk net4286 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21634_ clknet_leaf_125_i_clk net3300 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21565_ net199 net2458 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20516_ clknet_1_1__leaf__03849_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__buf_1
XFILLER_0_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21496_ clknet_leaf_0_i_clk net2270 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ net7025 net2381 _04412_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4240 net3916 vssd1 vssd1 vccd1 vccd1 net4767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22117_ clknet_leaf_57_i_clk net5382 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4251 _06091_ vssd1 vssd1 vccd1 vccd1 net4778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4262 net3637 vssd1 vssd1 vccd1 vccd1 net4789 sky130_fd_sc_hd__buf_1
Xhold4273 net8114 vssd1 vssd1 vccd1 vccd1 net4800 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_122_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold4284 net3972 vssd1 vssd1 vccd1 vccd1 net4811 sky130_fd_sc_hd__clkbuf_1
Xhold4295 net8087 vssd1 vssd1 vccd1 vccd1 net4822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3550 _03082_ vssd1 vssd1 vccd1 vccd1 net4077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22048_ net490 net1531 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold3561 net4144 vssd1 vssd1 vccd1 vccd1 net4088 sky130_fd_sc_hd__clkbuf_1
Xhold3572 _03808_ vssd1 vssd1 vccd1 vccd1 net4099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3583 net7680 vssd1 vssd1 vccd1 vccd1 net4110 sky130_fd_sc_hd__clkbuf_2
Xhold3594 net4146 vssd1 vssd1 vccd1 vccd1 net4121 sky130_fd_sc_hd__clkbuf_2
Xhold2860 net5747 vssd1 vssd1 vccd1 vccd1 net3387 sky130_fd_sc_hd__dlygate4sd3_1
X_20409__160 clknet_1_1__leaf__03846_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__inv_2
Xhold2871 _03089_ vssd1 vssd1 vccd1 vccd1 net3398 sky130_fd_sc_hd__buf_4
X_14870_ _08001_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__inv_2
Xhold2882 net4916 vssd1 vssd1 vccd1 vccd1 net3409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 _09210_ vssd1 vssd1 vccd1 vccd1 net3420 sky130_fd_sc_hd__buf_1
X_13821_ _06991_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _09519_ _09598_ _09629_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _06577_ net579 vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__xnor2_1
X_10964_ net7194 net6705 _04298_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12703_ net50 _05850_ _05851_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__and3_1
X_16471_ _09559_ _09561_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _06812_ _06819_ _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__a21o_1
X_10895_ net7500 net6924 _04265_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ _02427_ _02428_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__or2b_1
X_15422_ _08514_ _08516_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19190_ _03167_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__buf_4
X_12634_ net4128 _05043_ net22 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ _02365_ _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__xnor2_1
X_15353_ _07991_ _07998_ _08004_ _08404_ _08010_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__o41a_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12565_ net19 net18 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ _07473_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__xnor2_2
X_11516_ net4132 _04703_ _04704_ net5965 _04705_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a221o_2
X_18072_ _02259_ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15284_ net4181 _06314_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__nand2_1
X_12496_ net5981 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ _09249_ _09600_ vssd1 vssd1 vccd1 vccd1 _10044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14235_ _07242_ _07194_ _07403_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ rbzero.spi_registers.texadd2\[0\] _04566_ _04567_ vssd1 vssd1 vccd1 vccd1
+ _04639_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14166_ _06696_ _07233_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__nor2_1
X_11378_ _04564_ _04568_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _06286_ _06287_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__nor2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _07266_ _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__nor2_1
X_18974_ net3224 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _02160_ _02161_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__nor2_1
X_13048_ _06221_ _06223_ _06184_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a21oi_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ _02092_ _02093_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16807_ _09833_ _09834_ vssd1 vssd1 vccd1 vccd1 _09835_ sky130_fd_sc_hd__or2b_1
X_19786__65 clknet_1_1__leaf__03510_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
X_17787_ _02024_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__xor2_1
X_20620__350 clknet_1_0__leaf__03867_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__inv_2
X_14999_ _08093_ net7727 vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19526_ net3368 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
X_16738_ _09752_ _09762_ vssd1 vssd1 vccd1 vccd1 _09774_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19457_ net1742 _03335_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16669_ net4512 _09737_ _09740_ _07968_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18408_ _02589_ _02590_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19388_ net6080 _03270_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7805 rbzero.wall_tracer.stepDistY\[7\] vssd1 vssd1 vccd1 vccd1 net8332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18339_ _05155_ net3565 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__nand2_1
Xhold7816 net4607 vssd1 vssd1 vccd1 vccd1 net8343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7827 _06676_ vssd1 vssd1 vccd1 vccd1 net8354 sky130_fd_sc_hd__buf_2
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7838 net4893 vssd1 vssd1 vccd1 vccd1 net8365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21350_ clknet_leaf_47_i_clk net5119 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20301_ net1215 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold700 _01289_ vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21281_ clknet_leaf_24_i_clk net4371 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03859_ clknet_0__03859_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03859_
+ sky130_fd_sc_hd__clkbuf_16
Xhold711 net6741 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold722 _00969_ vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
X_20232_ net7490 _03706_ net4561 _03765_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__o211a_1
Xhold733 net6326 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _01359_ vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold755 _02484_ vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold766 net6288 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 net6408 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold788 _01438_ vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
X_20163_ net3581 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
Xhold799 net6348 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2101 net3366 vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2112 _04226_ vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2123 _01082_ vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
X_20094_ net4748 _03682_ _03615_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__o21ai_1
Xhold2134 net2318 vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2145 _01350_ vssd1 vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1400 _04163_ vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2156 _04319_ vssd1 vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1411 net2718 vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_54_i_clk clknet_4_14__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold1422 net5633 vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2167 net7305 vssd1 vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _01536_ vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2178 _01280_ vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2189 _04310_ vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1444 _02999_ vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 net6787 vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1466 _01555_ vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1477 _03412_ vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1488 net6885 vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1499 net6939 vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20996_ clknet_leaf_81_i_clk _00483_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_i_clk clknet_4_13__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10680_ net2033 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21617_ clknet_leaf_98_i_clk net1708 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12350_ _05306_ _05517_ _04848_ _05033_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21548_ net182 net2172 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ net71 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__inv_2
X_12281_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _05237_ vssd1 vssd1 vccd1 vccd1 _05467_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21479_ clknet_leaf_15_i_clk net1303 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11232_ net7119 net6868 _04434_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14020_ _07148_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__or2_4
XFILLER_0_205_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ net7504 net6460 _04401_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4070 net817 vssd1 vssd1 vccd1 vccd1 net4597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4081 net3587 vssd1 vssd1 vccd1 vccd1 net4608 sky130_fd_sc_hd__dlygate4sd3_1
X_15971_ _09059_ _09065_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__xor2_1
XFILLER_0_179_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11094_ net5673 net6184 _04364_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__mux2_1
Xhold4092 _01183_ vssd1 vssd1 vccd1 vccd1 net4619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17710_ _01737_ _01738_ _01838_ _01720_ _01718_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a311o_1
Xhold3380 _03343_ vssd1 vssd1 vccd1 vccd1 net3907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3391 _05064_ vssd1 vssd1 vccd1 vccd1 net3918 sky130_fd_sc_hd__dlygate4sd3_1
X_14922_ net8012 _08047_ _04482_ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__o21a_1
X_18690_ rbzero.wall_tracer.rayAddendY\[2\] _02843_ _02664_ vssd1 vssd1 vccd1 vccd1
+ _02844_ sky130_fd_sc_hd__mux2_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 net5987 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 _03240_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__nor2_1
Xhold82 net4949 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2690 net5977 vssd1 vssd1 vccd1 vccd1 net3217 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ net7794 _07956_ net4704 vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__a21oi_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 net4961 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _06968_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__nand2_1
X_17572_ _01807_ _01812_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__xnor2_1
X_14784_ _07948_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__clkbuf_1
X_11996_ net5947 _04600_ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__and3_1
X_19311_ net5085 _03250_ _03253_ _03246_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__o211a_1
X_16523_ _08127_ _09612_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13735_ net545 _06901_ _06905_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__o21a_1
X_10947_ net6107 net2110 _04287_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19242_ net6532 _03203_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__or2_1
X_16454_ _08025_ _08028_ _08030_ net75 vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__or4b_1
XFILLER_0_156_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13666_ _06834_ _06835_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10878_ net2924 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15405_ net8414 _08384_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ net27 net26 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19173_ net6253 _03170_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
X_16385_ _09348_ _09474_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__or2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ _06662_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18124_ _02350_ _02353_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__xnor2_1
X_15336_ net3417 rbzero.wall_tracer.visualWallDist\[-9\] _08117_ vssd1 vssd1 vccd1
+ vccd1 _08431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ _05727_ _05728_ net13 vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18055_ _02289_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__xnor2_1
X_15267_ _08360_ _08361_ _08114_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12479_ _05649_ _05657_ _05659_ _05660_ net9 vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__o2111a_1
XANTENNA_2 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17006_ _06124_ net4913 vssd1 vssd1 vccd1 vccd1 _10027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14218_ _07144_ _07145_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__and2_1
X_15198_ _08292_ _04695_ _08194_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__mux2_2
XFILLER_0_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14149_ _07312_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__xor2_2
X_18957_ net1146 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17908_ _02043_ _02044_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__nor2_1
X_18888_ net2162 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
X_17839_ _01784_ _09410_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor2_1
Xrebuffer14 net540 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer25 _06952_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 net562 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_1
X_20850_ _09736_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__clkbuf_4
Xrebuffer47 _06953_ vssd1 vssd1 vccd1 vccd1 net3523 sky130_fd_sc_hd__dlymetal6s4s_1
Xrebuffer58 _06734_ vssd1 vssd1 vccd1 vccd1 net3533 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19509_ net2205 net6739 _03365_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__mux2_1
X_20781_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7602 net1002 vssd1 vssd1 vccd1 vccd1 net8129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7613 rbzero.traced_texa\[-4\] vssd1 vssd1 vccd1 vccd1 net8140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7624 rbzero.traced_texa\[-11\] vssd1 vssd1 vccd1 vccd1 net8151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7635 rbzero.map_overlay.i_othery\[0\] vssd1 vssd1 vccd1 vccd1 net8162 sky130_fd_sc_hd__dlygate4sd3_1
X_21402_ clknet_leaf_41_i_clk net5051 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6901 rbzero.tex_g1\[24\] vssd1 vssd1 vccd1 vccd1 net7428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7646 rbzero.map_overlay.i_mapdx\[2\] vssd1 vssd1 vccd1 vccd1 net8173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6912 net2152 vssd1 vssd1 vccd1 vccd1 net7439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7657 _03713_ vssd1 vssd1 vccd1 vccd1 net8184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6923 rbzero.tex_b1\[50\] vssd1 vssd1 vccd1 vccd1 net7450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7668 rbzero.traced_texa\[2\] vssd1 vssd1 vccd1 vccd1 net8195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6934 net3131 vssd1 vssd1 vccd1 vccd1 net7461 sky130_fd_sc_hd__dlygate4sd3_1
X_21333_ clknet_leaf_6_i_clk net5171 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7679 rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 net8206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6945 rbzero.tex_g0\[15\] vssd1 vssd1 vccd1 vccd1 net7472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6956 rbzero.tex_g0\[28\] vssd1 vssd1 vccd1 vccd1 net7483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6967 net3153 vssd1 vssd1 vccd1 vccd1 net7494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6978 rbzero.pov.ss_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net7505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6989 net3233 vssd1 vssd1 vccd1 vccd1 net7516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold530 rbzero.pov.ready_buffer\[23\] vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
X_21264_ clknet_leaf_123_i_clk net2437 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold541 net5445 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold552 net8302 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_1
Xhold563 net6153 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
X_20215_ net4635 _03710_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold574 net7900 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21195_ clknet_leaf_126_i_clk net1648 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold585 _01140_ vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold596 net5453 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20146_ net3721 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20077_ net3317 _03660_ net4363 _03628_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__o211a_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _01540_ vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 net6678 vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 _03402_ vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__buf_2
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1263 _00696_ vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1274 _03465_ vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 net6521 vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 net5597 vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _04706_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__inv_2
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19765__46 clknet_1_1__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
XFILLER_0_135_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ net6170 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _04969_ _04970_ _04847_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20979_ clknet_leaf_57_i_clk _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_138_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13520_ _06687_ _06688_ _06690_ _06632_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__o22ai_1
X_10732_ net6798 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13451_ _06490_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__or3_1
X_10663_ net6279 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12402_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _04924_ vssd1 vssd1 vccd1 vccd1 _05587_
+ sky130_fd_sc_hd__mux2_1
X_16170_ _08211_ _09262_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__nor2_1
X_10594_ net7289 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__clkbuf_1
X_13382_ _06549_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ net4236 _08215_ _08123_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__mux2_1
X_12333_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _04913_ vssd1 vssd1 vccd1 vccd1 _05519_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15052_ net3489 _06033_ _08123_ _08146_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12264_ net4335 _05306_ _05018_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14003_ _07172_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__nor2_1
X_11215_ _04264_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__clkbuf_4
X_12195_ rbzero.tex_g1\[15\] rbzero.tex_g1\[14\] _05249_ vssd1 vssd1 vccd1 vccd1 _05382_
+ sky130_fd_sc_hd__mux2_1
X_19860_ net2312 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__buf_1
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__clkbuf_4
X_18811_ net1547 net3909 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__nor2_1
X_11146_ net6534 net2987 _04390_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15954_ _08400_ _08485_ _09048_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__a21oi_1
X_11077_ net2274 net6699 _04353_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
X_18742_ _02856_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02892_
+ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14905_ _06237_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__clkbuf_4
X_18673_ net3575 _05164_ _02826_ _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nor4_2
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _08934_ _08978_ _08979_ vssd1 vssd1 vccd1 vccd1 _08980_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17624_ _01861_ _01862_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__or2_1
X_14836_ _07860_ _07830_ _07878_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__a21oi_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _01793_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _07843_ _07876_ _07879_ _07932_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__a31o_1
X_11979_ _04670_ net4127 _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and3_1
X_16506_ _09593_ _09595_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__xnor2_1
X_13718_ _06702_ _06692_ _06705_ net556 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__or4b_1
X_17486_ _01723_ _01726_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ net4704 vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__clkbuf_4
X_16437_ _08509_ _08411_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19225_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__buf_2
X_13649_ _06812_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20669__15 clknet_1_0__leaf__03871_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_0_211_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19156_ net1319 _03146_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__or2_1
X_16368_ _09336_ _09321_ _09448_ vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__a21o_1
Xhold6208 net1853 vssd1 vssd1 vccd1 vccd1 net6735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__05794_ clknet_0__05794_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05794_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6219 net1761 vssd1 vssd1 vccd1 vccd1 net6746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ net3731 _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__nor2_1
X_15319_ _08413_ _08367_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__nand2_2
XFILLER_0_125_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5507 net630 vssd1 vssd1 vccd1 vccd1 net6034 sky130_fd_sc_hd__dlygate4sd3_1
X_19087_ net3042 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__clkbuf_1
X_16299_ _08246_ _08414_ _09276_ _09279_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5518 _01253_ vssd1 vssd1 vccd1 vccd1 net6045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5529 net1625 vssd1 vssd1 vccd1 vccd1 net6056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _02272_ _02273_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__xnor2_1
Xhold4806 _00808_ vssd1 vssd1 vccd1 vccd1 net5333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4817 net1000 vssd1 vssd1 vccd1 vccd1 net5344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4828 rbzero.color_sky\[0\] vssd1 vssd1 vccd1 vccd1 net5355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4839 net930 vssd1 vssd1 vccd1 vccd1 net5366 sky130_fd_sc_hd__dlygate4sd3_1
X_20349__106 clknet_1_1__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__inv_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20000_ _03609_ net5817 vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__or2_1
XFILLER_0_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19989_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21951_ net393 net1315 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ clknet_leaf_37_i_clk net5620 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_21882_ net324 net3265 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ net3976 _03992_ _03993_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__o21a_1
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20764_ net948 net5492 vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20695_ net756 net4984 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7410 rbzero.wall_tracer.stepDistX\[-9\] vssd1 vssd1 vccd1 vccd1 net7937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7421 net4499 vssd1 vssd1 vccd1 vccd1 net7948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7432 rbzero.wall_tracer.trackDistY\[6\] vssd1 vssd1 vccd1 vccd1 net7959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7443 net4650 vssd1 vssd1 vccd1 vccd1 net7970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7454 rbzero.wall_tracer.trackDistX\[-5\] vssd1 vssd1 vccd1 vccd1 net7981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6720 rbzero.tex_b0\[38\] vssd1 vssd1 vccd1 vccd1 net7247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7465 net3819 vssd1 vssd1 vccd1 vccd1 net7992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6731 net2832 vssd1 vssd1 vccd1 vccd1 net7258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7476 _00516_ vssd1 vssd1 vccd1 vccd1 net8003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6742 rbzero.tex_b0\[32\] vssd1 vssd1 vccd1 vccd1 net7269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7487 net4254 vssd1 vssd1 vccd1 vccd1 net8014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6753 rbzero.tex_b0\[12\] vssd1 vssd1 vccd1 vccd1 net7280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7498 _02800_ vssd1 vssd1 vccd1 vccd1 net8025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6764 net2575 vssd1 vssd1 vccd1 vccd1 net7291 sky130_fd_sc_hd__dlygate4sd3_1
X_21316_ clknet_leaf_4_i_clk net5338 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6775 rbzero.spi_registers.new_mapd\[5\] vssd1 vssd1 vccd1 vccd1 net7302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6786 rbzero.tex_g0\[8\] vssd1 vssd1 vccd1 vccd1 net7313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6797 net2370 vssd1 vssd1 vccd1 vccd1 net7324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21247_ clknet_leaf_21_i_clk net3598 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold360 net6066 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 net5275 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold382 net5307 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net5574 net5653 _04320_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__mux2_1
Xhold393 net6059 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
X_21178_ clknet_leaf_98_i_clk net1877 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20129_ net7593 _03707_ net4473 _03679_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12951_ net3999 _06039_ net3848 _06104_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_172_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 net6586 vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 _01406_ vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _04666_ net4058 _05072_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a21boi_1
X_15670_ _08741_ _08743_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__xor2_2
Xhold1082 net8108 vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12882_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__buf_4
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _00684_ vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _07305_ _07339_ _07440_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__and3b_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ net3781 net3648 _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and3_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _10357_ _10358_ vssd1 vssd1 vccd1 vccd1 _10359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _07706_ _07721_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__a21oi_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _04910_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__or2_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _06445_ _06447_ _06450_ _06453_ _06493_ _06553_ vssd1 vssd1 vccd1 vccd1 _06674_
+ sky130_fd_sc_hd__mux4_1
X_17271_ _09133_ _10289_ vssd1 vssd1 vccd1 vccd1 _10290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ net5991 net5630 _04171_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__mux2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _07606_ _07653_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ _04882_ _04883_ _04884_ net4145 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19010_ net3485 net3935 net1547 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__or3_1
X_16222_ _09219_ _09220_ _09314_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _06568_ _06604_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__nand2_1
X_10646_ net2951 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16153_ _09139_ _09148_ _09146_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer5 net7787 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13365_ _06527_ _06529_ _06535_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__and3_1
X_10577_ net1958 net6554 _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__mux2_1
X_15104_ _08194_ _08198_ _06120_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__o21a_1
X_12316_ _05500_ _05501_ _04984_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16084_ _09175_ _09176_ _09036_ _09177_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13296_ _06413_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__buf_2
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ net4917 _08129_ vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19912_ net2975 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
X_12247_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _04933_ vssd1 vssd1 vccd1 vccd1 _05434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03512_ _03512_ vssd1 vssd1 vccd1 vccd1 clknet_0__03512_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19843_ net3102 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
X_12178_ _05360_ _05362_ _05365_ _04988_ net85 vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11129_ net6904 net6946 _04309_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ _09460_ _09587_ _09710_ _10007_ vssd1 vssd1 vccd1 vccd1 _10008_ sky130_fd_sc_hd__o31a_4
X_18725_ _02868_ _02876_ _02526_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
X_15937_ _08458_ _09031_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15868_ _08958_ _08960_ _08962_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__o21ai_1
X_18656_ _02809_ _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__xnor2_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17607_ net3875 net4624 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__nor2_1
X_14819_ _07935_ _07965_ _07966_ _07978_ _07913_ net7785 vssd1 vssd1 vccd1 vccd1 _07979_
+ sky130_fd_sc_hd__mux4_2
X_15799_ _08854_ _08857_ _08891_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18587_ net4019 _02748_ net89 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_140 vssd1 vssd1 vccd1 vccd1 ones[13] top_ew_algofoogle_140/LO sky130_fd_sc_hd__conb_1
XFILLER_0_176_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ _01777_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17469_ _01709_ _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__05946_ _05946_ vssd1 vssd1 vccd1 vccd1 clknet_0__05946_ sky130_fd_sc_hd__clkbuf_16
X_19208_ net5149 _03182_ _03192_ _03189_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6005 net1800 vssd1 vssd1 vccd1 vccd1 net6532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6016 rbzero.spi_registers.new_vshift\[4\] vssd1 vssd1 vccd1 vccd1 net6543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6027 net1383 vssd1 vssd1 vccd1 vccd1 net6554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19139_ net1133 _03147_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__or2_1
Xhold6038 rbzero.spi_registers.new_texadd\[0\]\[9\] vssd1 vssd1 vccd1 vccd1 net6565
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold5304 _02558_ vssd1 vssd1 vccd1 vccd1 net5831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6049 net1638 vssd1 vssd1 vccd1 vccd1 net6576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5315 net3742 vssd1 vssd1 vccd1 vccd1 net5842 sky130_fd_sc_hd__dlygate4sd3_1
X_22150_ clknet_leaf_51_i_clk _01637_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5326 net3458 vssd1 vssd1 vccd1 vccd1 net5853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5337 _02972_ vssd1 vssd1 vccd1 vccd1 net5864 sky130_fd_sc_hd__buf_1
XFILLER_0_160_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5348 _00605_ vssd1 vssd1 vccd1 vccd1 net5875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4603 _00831_ vssd1 vssd1 vccd1 vccd1 net5130 sky130_fd_sc_hd__dlygate4sd3_1
X_21101_ clknet_leaf_0_i_clk net1373 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5359 rbzero.debug_overlay.playerX\[-6\] vssd1 vssd1 vccd1 vccd1 net5886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4614 net738 vssd1 vssd1 vccd1 vccd1 net5141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4625 rbzero.spi_registers.texadd3\[16\] vssd1 vssd1 vccd1 vccd1 net5152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22081_ net523 net1237 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4636 net794 vssd1 vssd1 vccd1 vccd1 net5163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3902 net7918 vssd1 vssd1 vccd1 vccd1 net4429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4647 _00872_ vssd1 vssd1 vccd1 vccd1 net5174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3913 net3551 vssd1 vssd1 vccd1 vccd1 net4440 sky130_fd_sc_hd__buf_1
Xhold4658 net862 vssd1 vssd1 vccd1 vccd1 net5185 sky130_fd_sc_hd__dlygate4sd3_1
X_21032_ clknet_leaf_55_i_clk net4267 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4669 rbzero.spi_registers.texadd3\[19\] vssd1 vssd1 vccd1 vccd1 net5196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3924 _03142_ vssd1 vssd1 vccd1 vccd1 net4451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3935 rbzero.debug_overlay.facingX\[-6\] vssd1 vssd1 vccd1 vccd1 net4462 sky130_fd_sc_hd__buf_1
Xhold3946 net8179 vssd1 vssd1 vccd1 vccd1 net4473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3957 net8326 vssd1 vssd1 vccd1 vccd1 net4484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3968 net8394 vssd1 vssd1 vccd1 vccd1 net4495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3979 net3718 vssd1 vssd1 vccd1 vccd1 net4506 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21934_ net376 net2087 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20403__155 clknet_1_0__leaf__03845_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__inv_2
XFILLER_0_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21865_ net307 net1717 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ net1028 net5480 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21796_ net238 net662 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20747_ _03920_ _03921_ _03919_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ net2260 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11480_ net4176 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__buf_2
XFILLER_0_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7240 rbzero.debug_overlay.playerY\[-6\] vssd1 vssd1 vccd1 vccd1 net7767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7251 _09104_ vssd1 vssd1 vccd1 vccd1 net7778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7262 net4434 vssd1 vssd1 vccd1 vccd1 net7789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7284 _06494_ vssd1 vssd1 vccd1 vccd1 net7811 sky130_fd_sc_hd__buf_2
Xhold6550 net2665 vssd1 vssd1 vccd1 vccd1 net7077 sky130_fd_sc_hd__dlygate4sd3_1
X_13150_ _06288_ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__xnor2_2
Xhold6561 rbzero.tex_b0\[35\] vssd1 vssd1 vccd1 vccd1 net7088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6572 net2357 vssd1 vssd1 vccd1 vccd1 net7099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6583 rbzero.tex_g1\[7\] vssd1 vssd1 vccd1 vccd1 net7110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6594 net2548 vssd1 vssd1 vccd1 vccd1 net7121 sky130_fd_sc_hd__dlygate4sd3_1
X_12101_ _05203_ _05284_ _05286_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5860 rbzero.spi_registers.new_texadd\[0\]\[13\] vssd1 vssd1 vccd1 vccd1 net6387
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13081_ net5618 _06244_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__xnor2_1
Xhold5871 rbzero.spi_registers.new_texadd\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net6398
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5882 net1304 vssd1 vssd1 vccd1 vccd1 net6409 sky130_fd_sc_hd__dlygate4sd3_1
X_20484__227 clknet_1_1__leaf__03854_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__inv_2
Xhold5893 _03463_ vssd1 vssd1 vccd1 vccd1 net6420 sky130_fd_sc_hd__dlygate4sd3_1
X_12032_ rbzero.tex_r1\[13\] rbzero.tex_r1\[12\] _05220_ vssd1 vssd1 vccd1 vccd1 _05221_
+ sky130_fd_sc_hd__mux2_1
Xhold190 net5024 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _09862_ _09863_ _09864_ vssd1 vssd1 vccd1 vccd1 _09865_ sky130_fd_sc_hd__o21ai_1
X_16771_ _09802_ net4506 _09769_ vssd1 vssd1 vccd1 vccd1 _09803_ sky130_fd_sc_hd__mux2_1
X_13983_ _06693_ net573 _07109_ _06577_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_137_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15722_ _08815_ _08816_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__xor2_1
X_18510_ _02677_ _02678_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12934_ net4431 net3999 vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__xor2_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ net2233 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _08725_ _08747_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__nor2_1
X_18441_ net4791 _02619_ _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a21oi_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _06038_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__nor2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _07696_ _07731_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__nand2_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20378__132 clknet_1_1__leaf__03843_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__inv_2
XFILLER_0_157_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11816_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _04836_ vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18372_ rbzero.wall_tracer.rayAddendX\[-2\] _02557_ _02537_ vssd1 vssd1 vccd1 vccd1
+ _02558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _08220_ _08678_ _08271_ _08252_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__or4b_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ _05971_ _05962_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__or2b_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17323_ _09272_ _09664_ vssd1 vssd1 vccd1 vccd1 _10342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _07704_ _07705_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__and2_1
X_11747_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _04912_ vssd1 vssd1 vccd1 vccd1 _04937_
+ sky130_fd_sc_hd__mux2_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17254_ _10179_ _10271_ _10272_ vssd1 vssd1 vccd1 vccd1 _10273_ sky130_fd_sc_hd__a21oi_2
X_14466_ _07489_ _07233_ _07281_ _07072_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ net3488 _04857_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16205_ _09177_ _09297_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__xor2_2
X_13417_ _06568_ _06560_ _06562_ net559 vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__o31ai_1
X_10629_ net1895 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__clkbuf_1
X_17185_ _10184_ _10203_ vssd1 vssd1 vccd1 vccd1 _10205_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14397_ _07562_ _07566_ _07567_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16136_ _08542_ _08616_ _09137_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13348_ _06505_ _06506_ _06485_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _09155_ _09160_ vssd1 vssd1 vccd1 vccd1 _09161_ sky130_fd_sc_hd__xnor2_1
X_13279_ _06448_ _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__xnor2_4
Xhold3209 _00609_ vssd1 vssd1 vccd1 vccd1 net3736 sky130_fd_sc_hd__dlygate4sd3_1
X_15018_ _08112_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__buf_4
Xhold2508 net3332 vssd1 vssd1 vccd1 vccd1 net3035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 _03522_ vssd1 vssd1 vccd1 vccd1 net3046 sky130_fd_sc_hd__dlygate4sd3_1
X_19826_ net2507 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
Xhold1807 _04346_ vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1818 net7331 vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1829 _01348_ vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
X_16969_ _09953_ _09990_ vssd1 vssd1 vccd1 vccd1 _09991_ sky130_fd_sc_hd__xnor2_1
X_18708_ net4797 _02858_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19688_ net6370 net3596 _03468_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _02789_ _02790_ _02796_ _04481_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__a22o_1
X_21650_ clknet_leaf_117_i_clk net2413 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21581_ net215 net3119 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5101 net2836 vssd1 vssd1 vccd1 vccd1 net5628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5112 net2374 vssd1 vssd1 vccd1 vccd1 net5639 sky130_fd_sc_hd__dlygate4sd3_1
X_20394_ clknet_1_1__leaf__03513_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__buf_1
Xhold5123 _04357_ vssd1 vssd1 vccd1 vccd1 net5650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5134 net2343 vssd1 vssd1 vccd1 vccd1 net5661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5145 rbzero.tex_b1\[15\] vssd1 vssd1 vccd1 vccd1 net5672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4400 gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4411 net601 vssd1 vssd1 vccd1 vccd1 net4938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5156 rbzero.tex_b1\[3\] vssd1 vssd1 vccd1 vccd1 net5683 sky130_fd_sc_hd__dlygate4sd3_1
X_22133_ clknet_leaf_56_i_clk net5482 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5167 net2495 vssd1 vssd1 vccd1 vccd1 net5694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4422 _01657_ vssd1 vssd1 vccd1 vccd1 net4949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5178 rbzero.tex_r0\[49\] vssd1 vssd1 vccd1 vccd1 net5705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4433 net619 vssd1 vssd1 vccd1 vccd1 net4960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5189 net2698 vssd1 vssd1 vccd1 vccd1 net5716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4444 rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 net4971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4455 net651 vssd1 vssd1 vccd1 vccd1 net4982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3710 net8139 vssd1 vssd1 vccd1 vccd1 net4237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3721 net8016 vssd1 vssd1 vccd1 vccd1 net4248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4466 _00858_ vssd1 vssd1 vccd1 vccd1 net4993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3732 net8145 vssd1 vssd1 vccd1 vccd1 net4259 sky130_fd_sc_hd__clkbuf_2
X_22064_ net506 net2643 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4477 rbzero.spi_registers.texadd0\[3\] vssd1 vssd1 vccd1 vccd1 net5004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3743 net1049 vssd1 vssd1 vccd1 vccd1 net4270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4488 net688 vssd1 vssd1 vccd1 vccd1 net5015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3754 net8142 vssd1 vssd1 vccd1 vccd1 net4281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4499 _00867_ vssd1 vssd1 vccd1 vccd1 net5026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3765 net992 vssd1 vssd1 vccd1 vccd1 net4292 sky130_fd_sc_hd__dlygate4sd3_1
X_21015_ clknet_leaf_62_i_clk net4320 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3776 net8311 vssd1 vssd1 vccd1 vccd1 net4303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3787 net1035 vssd1 vssd1 vccd1 vccd1 net4314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3798 _00763_ vssd1 vssd1 vccd1 vccd1 net4325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ net2355 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
X_21917_ net359 net2478 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _04648_ _04461_ _04468_ _04023_ _05802_ _05797_ vssd1 vssd1 vccd1 vccd1 _05829_
+ sky130_fd_sc_hd__mux4_1
X_21848_ net290 net3165 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ net950 net1217 net1233 net1008 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _05758_ _05759_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__mux2_1
X_21779_ clknet_leaf_9_i_clk net1202 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _07072_ _06754_ _07303_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__or3_1
XFILLER_0_167_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11532_ net4315 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _07417_ _07421_ _07418_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__a21oi_1
X_11463_ net2 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7070 net3481 vssd1 vssd1 vccd1 vccd1 net7597 sky130_fd_sc_hd__dlygate4sd3_1
X_13202_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__inv_2
Xhold7081 rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 net7608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14182_ _07345_ _07349_ _07352_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__a21oi_1
Xhold7092 _03793_ vssd1 vssd1 vccd1 vccd1 net7619 sky130_fd_sc_hd__dlygate4sd3_1
X_11394_ _04558_ _04559_ _04560_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6380 _04112_ vssd1 vssd1 vccd1 vccd1 net6907 sky130_fd_sc_hd__dlygate4sd3_1
X_13133_ net4446 net5952 vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__nand2_2
Xhold6391 net2405 vssd1 vssd1 vccd1 vccd1 net6918 sky130_fd_sc_hd__dlygate4sd3_1
X_18990_ net2927 net5783 _03058_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5690 net1149 vssd1 vssd1 vccd1 vccd1 net6217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _02176_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__xnor2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ net4647 _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__nand2_2
XFILLER_0_178_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12015_ _04977_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17872_ _09915_ net4891 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19611_ _03429_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__buf_4
X_16823_ _09849_ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19542_ net5513 net1396 _03388_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__mux2_1
X_13966_ _07135_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__and2b_1
X_16754_ net3976 _04476_ net3871 vssd1 vssd1 vccd1 vccd1 _09787_ sky130_fd_sc_hd__nor3b_2
X_19801__78 clknet_1_1__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15705_ _08326_ _08329_ _08691_ _08799_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__o22ai_2
X_12917_ _06075_ _06087_ net4778 _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__o211a_1
X_16685_ _09738_ vssd1 vssd1 vccd1 vccd1 _09744_ sky130_fd_sc_hd__clkbuf_4
X_19473_ net4016 net6005 _03345_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13897_ _07023_ _07022_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18424_ net5972 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15636_ _08186_ _08433_ _08730_ _08662_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12848_ _06023_ _05996_ _05971_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o21a_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _08661_ _08474_ _08630_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__o21ai_1
X_18355_ net4698 rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _02542_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _05953_
+ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a31o_4
XFILLER_0_185_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17306_ _09262_ _09165_ vssd1 vssd1 vccd1 vccd1 _10325_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14518_ _07665_ _07687_ _07688_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15498_ _08568_ _08569_ _08585_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18286_ net6405 net3402 _02477_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17237_ _10253_ _10256_ vssd1 vssd1 vccd1 vccd1 _10257_ sky130_fd_sc_hd__xnor2_4
X_14449_ _07618_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ _10063_ _10187_ vssd1 vssd1 vccd1 vccd1 _10188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold904 _00945_ vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 _03822_ vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 net6369 vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
X_20432__181 clknet_1_0__leaf__03848_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__inv_2
Xclkbuf_0__05645_ _05645_ vssd1 vssd1 vccd1 vccd1 clknet_0__05645_ sky130_fd_sc_hd__clkbuf_16
X_16119_ _09086_ _09099_ _09211_ vssd1 vssd1 vccd1 vccd1 _09213_ sky130_fd_sc_hd__and3_1
Xhold937 _01003_ vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold948 _03826_ vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_17099_ _10058_ _10119_ vssd1 vssd1 vccd1 vccd1 _10120_ sky130_fd_sc_hd__xnor2_2
Xhold959 net6614 vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3017 _03622_ vssd1 vssd1 vccd1 vccd1 net3544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3028 _01195_ vssd1 vssd1 vccd1 vccd1 net3555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3039 _03750_ vssd1 vssd1 vccd1 vccd1 net3566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2305 net7257 vssd1 vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2316 _01057_ vssd1 vssd1 vccd1 vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2327 net7300 vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 _00711_ vssd1 vssd1 vccd1 vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1604 net6757 vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 _00699_ vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 _01497_ vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1626 net5548 vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1637 net7112 vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 _01556_ vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 net5572 vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21702_ clknet_leaf_118_i_clk net5774 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21633_ clknet_leaf_124_i_clk net1360 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21564_ net198 net906 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20515__256 clknet_1_0__leaf__03856_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__inv_2
XFILLER_0_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21495_ clknet_leaf_7_i_clk net1330 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4230 net4262 vssd1 vssd1 vccd1 vccd1 net4757 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22116_ clknet_leaf_55_i_clk net5402 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
Xhold4241 net8352 vssd1 vssd1 vccd1 vccd1 net4768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4252 _06093_ vssd1 vssd1 vccd1 vccd1 net4779 sky130_fd_sc_hd__buf_1
XFILLER_0_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4274 net1676 vssd1 vssd1 vccd1 vccd1 net4801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4285 net8052 vssd1 vssd1 vccd1 vccd1 net4812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3540 _05056_ vssd1 vssd1 vccd1 vccd1 net4067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3551 _00724_ vssd1 vssd1 vccd1 vccd1 net4078 sky130_fd_sc_hd__dlygate4sd3_1
X_22047_ net489 net1277 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold4296 net3948 vssd1 vssd1 vccd1 vccd1 net4823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3562 _04025_ vssd1 vssd1 vccd1 vccd1 net4089 sky130_fd_sc_hd__buf_4
Xhold3573 _01252_ vssd1 vssd1 vccd1 vccd1 net4100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3584 _05672_ vssd1 vssd1 vccd1 vccd1 net4111 sky130_fd_sc_hd__clkbuf_4
Xhold2850 _00944_ vssd1 vssd1 vccd1 vccd1 net3377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3595 _09718_ vssd1 vssd1 vccd1 vccd1 net4122 sky130_fd_sc_hd__clkbuf_4
Xhold2861 net8313 vssd1 vssd1 vccd1 vccd1 net3388 sky130_fd_sc_hd__clkbuf_2
Xhold2872 _03092_ vssd1 vssd1 vccd1 vccd1 net3399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2883 net4509 vssd1 vssd1 vccd1 vccd1 net3410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2894 net7992 vssd1 vssd1 vccd1 vccd1 net3421 sky130_fd_sc_hd__dlygate4sd3_1
X_13820_ net552 _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20596__328 clknet_1_0__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__inv_2
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ net547 _06912_ _06921_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__o21ai_1
X_10963_ net3030 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12702_ net30 _05872_ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__o21a_1
X_16470_ _09401_ _09429_ _09560_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__a21oi_1
X_13682_ _06820_ _06810_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ net7479 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _08358_ _08515_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__nand2_1
X_12633_ net4103 net4024 _05730_ net3996 net22 net25 vssd1 vssd1 vccd1 vccd1 _05812_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15352_ _08436_ _08422_ _08437_ _08360_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__and4_1
X_18140_ _02366_ _02367_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__or2b_1
X_12564_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14303_ _06914_ _07197_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__nor2_1
X_18071_ _02264_ _02306_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__xor2_1
X_11515_ net6044 net4145 net1 vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or3b_1
XFILLER_0_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15283_ _04476_ net3452 vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12495_ net4102 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__buf_1
X_17022_ _10040_ _10041_ _10042_ _09617_ vssd1 vssd1 vccd1 vccd1 _10043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14234_ _07403_ _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11446_ _04502_ _04633_ _04634_ _04635_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__o32a_1
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ _06699_ _07281_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11377_ _04564_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _07207_ _07248_ _07265_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__and3_1
X_18973_ net3312 net5737 net2874 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _01815_ _02066_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__and2b_1
X_13047_ _06166_ _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__or2_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17855_ _02070_ _02091_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ net4547 net4583 vssd1 vssd1 vccd1 vccd1 _09834_ sky130_fd_sc_hd__nand2_1
X_17786_ _01794_ _10096_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ net4165 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
X_19525_ net3863 net3367 net3086 vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__mux2_1
X_16737_ net5472 _09102_ vssd1 vssd1 vccd1 vccd1 _09773_ sky130_fd_sc_hd__xor2_1
X_13949_ _06846_ _07119_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19456_ net4230 _03334_ net1366 _03339_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__o211a_1
X_16668_ net4305 _09737_ _09740_ _07962_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18407_ net3509 _05155_ _02587_ _02588_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__o22a_1
X_15619_ _08266_ _08318_ _08679_ _08681_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19387_ net4988 _03268_ _03296_ _03288_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__o211a_1
X_16599_ _09684_ _09685_ _09687_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18338_ _04478_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__buf_4
Xhold7806 net4536 vssd1 vssd1 vccd1 vccd1 net8333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7817 rbzero.wall_tracer.trackDistX\[-11\] vssd1 vssd1 vccd1 vccd1 net8344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7828 _07104_ vssd1 vssd1 vccd1 vccd1 net8355 sky130_fd_sc_hd__buf_2
Xhold7839 rbzero.wall_tracer.stepDistY\[-1\] vssd1 vssd1 vccd1 vccd1 net8366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18269_ net1397 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20300_ net6265 net3402 _03814_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21280_ clknet_leaf_25_i_clk net4356 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03858_ clknet_0__03858_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03858_
+ sky130_fd_sc_hd__clkbuf_16
Xhold701 net5479 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold712 _03152_ vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 net5798 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20231_ net4560 _03710_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__or2_1
Xhold734 net6328 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 net6499 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold756 _00575_ vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold767 _00954_ vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
X_20162_ _03728_ net7643 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__or2_1
Xhold778 _03818_ vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold789 net6412 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2102 _03127_ vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2113 _01424_ vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20093_ net616 _03631_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__or2_1
Xhold2124 net7249 vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 _04167_ vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1401 _01481_ vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2146 net7390 vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2157 _01340_ vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1412 _04073_ vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 net5635 vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 net7307 vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2179 net7345 vssd1 vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 net6807 vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1445 _00652_ vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 net6789 vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1467 net6795 vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1478 _00953_ vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 _01391_ vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20995_ clknet_leaf_52_i_clk net4081 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21616_ clknet_leaf_97_i_clk net3065 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21547_ net181 net1911 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ net8217 _04486_ _04487_ _04483_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a31o_1
X_12280_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _05237_ vssd1 vssd1 vccd1 vccd1 _05466_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21478_ clknet_leaf_19_i_clk net4818 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11231_ net6782 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11162_ net7379 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4060 net1664 vssd1 vssd1 vccd1 vccd1 net4587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4071 net8248 vssd1 vssd1 vccd1 vccd1 net4598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4082 net7963 vssd1 vssd1 vccd1 vccd1 net4609 sky130_fd_sc_hd__dlygate4sd3_1
X_15970_ _08615_ _09063_ _09064_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__o21ba_1
X_11093_ net2368 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
Xhold4093 net3490 vssd1 vssd1 vccd1 vccd1 net4620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3370 net1621 vssd1 vssd1 vccd1 vccd1 net3897 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3381 _00903_ vssd1 vssd1 vccd1 vccd1 net3908 sky130_fd_sc_hd__dlygate4sd3_1
X_14921_ net4657 _08050_ _08052_ net3766 net4691 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__o221a_1
Xhold3392 _05065_ vssd1 vssd1 vccd1 vccd1 net3919 sky130_fd_sc_hd__buf_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2680 net3301 vssd1 vssd1 vccd1 vccd1 net3207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 net5989 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _01873_ _01788_ _01878_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__and3_1
Xhold72 net4199 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net5044 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2691 net5979 vssd1 vssd1 vccd1 vccd1 net3218 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _07934_ _08006_ _08007_ net7824 vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 net4963 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1990 _01431_ vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _06968_ _06969_ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__nand3_1
X_17571_ _01810_ _01811_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__xnor2_1
X_14783_ net4379 _07947_ _07872_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__mux2_1
X_11995_ _04022_ _04467_ _04460_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__and3_1
X_19310_ net1859 _03251_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__or2_1
X_16522_ _09472_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__buf_4
X_13734_ net558 _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__or2b_1
X_10946_ net2483 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19241_ net5228 _03201_ _03212_ _03206_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13665_ _06834_ _06835_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__nor2_1
X_16453_ _08024_ _09414_ net75 _09543_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__a31o_1
X_10877_ net7355 net7186 _04253_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12616_ _05795_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _08488_ _08490_ _08498_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16384_ _09348_ _09474_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19172_ net5053 _03168_ _03172_ _03160_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__o211a_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _06761_ _06766_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__xor2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15335_ _08427_ _08428_ _08429_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__a21o_2
X_18123_ _02351_ _02352_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12547_ net4111 _05673_ net4071 net4092 _05691_ net12 vssd1 vssd1 vccd1 vccd1 _05728_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20650__377 clknet_1_0__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__inv_2
XFILLER_0_124_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _08472_ _09612_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__nor2_1
X_15266_ _07968_ _07975_ _07981_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__or3_1
X_12478_ net7 net6 net8 vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a21o_1
XANTENNA_3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17005_ _09952_ _09931_ vssd1 vssd1 vccd1 vccd1 _10026_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14217_ _06699_ _07327_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ _04021_ _04531_ _04620_ _04584_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15197_ net3461 _08261_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14148_ _07317_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14079_ _07104_ _06576_ net541 _06914_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__or4_1
X_18956_ net2801 net7573 _03036_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
X_17907_ _01966_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18887_ net3077 net7021 _03003_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20544__282 clknet_1_1__leaf__03859_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__inv_2
X_17838_ _10062_ _09540_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer15 net541 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 _08439_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer37 _07832_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_1
X_17769_ _02006_ _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__nand2_1
Xrebuffer48 _06643_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_1
Xrebuffer59 net3533 vssd1 vssd1 vccd1 vccd1 net3579 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19508_ net1672 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20780_ _03948_ _03949_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19439_ net4952 _03323_ _03329_ _03316_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_121_i_clk clknet_4_1__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7603 _00624_ vssd1 vssd1 vccd1 vccd1 net8130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7614 net1106 vssd1 vssd1 vccd1 vccd1 net8141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21401_ clknet_leaf_41_i_clk net3673 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7625 rbzero.map_overlay.i_othery\[4\] vssd1 vssd1 vccd1 vccd1 net8152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7636 rbzero.map_overlay.i_othery\[2\] vssd1 vssd1 vccd1 vccd1 net8163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6902 net2996 vssd1 vssd1 vccd1 vccd1 net7429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7647 rbzero.spi_registers.got_new_texadd\[3\] vssd1 vssd1 vccd1 vccd1 net8174
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold6913 rbzero.tex_r0\[43\] vssd1 vssd1 vccd1 vccd1 net7440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6924 net2667 vssd1 vssd1 vccd1 vccd1 net7451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7669 rbzero.traced_texa\[-1\] vssd1 vssd1 vccd1 vccd1 net8196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6935 _03039_ vssd1 vssd1 vccd1 vccd1 net7462 sky130_fd_sc_hd__dlygate4sd3_1
X_21332_ clknet_leaf_8_i_clk net5147 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6946 net3029 vssd1 vssd1 vccd1 vccd1 net7473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6957 net3263 vssd1 vssd1 vccd1 vccd1 net7484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6968 rbzero.spi_registers.sclk_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net7495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6979 net2309 vssd1 vssd1 vccd1 vccd1 net7506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold520 net5449 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
X_21263_ clknet_leaf_122_i_clk net2048 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi
+ sky130_fd_sc_hd__dfxtp_1
Xhold531 net7946 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 net6183 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold553 net6163 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
X_20214_ net4825 _03743_ _03767_ _03765_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__o211a_1
Xhold564 _01483_ vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold575 net2933 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
X_21194_ clknet_leaf_126_i_clk net3275 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold586 net7592 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 net5687 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20145_ _03689_ net3720 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ net4362 _03485_ _03662_ _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a211o_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _01008_ vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 net6849 vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 _01271_ vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 _03418_ vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1264 net8331 vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1275 _00997_ vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _00981_ vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 net6801 vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ net1985 net6168 _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__mux2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _04837_ vssd1 vssd1 vccd1 vccd1 _04970_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20978_ clknet_leaf_81_i_clk net4184 vssd1 vssd1 vccd1 vccd1 rbzero.side_hot sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ net6796 net2049 _04097_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _06491_ _06600_ _06601_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__and3_1
X_10662_ net6277 net2140 _04138_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12401_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _05369_ vssd1 vssd1 vccd1 vccd1 _05586_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ _06522_ _06499_ _06461_ _06548_ _06549_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_
+ sky130_fd_sc_hd__mux4_2
X_10593_ net7287 net2914 _04105_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15120_ _08214_ net4344 _06027_ vssd1 vssd1 vccd1 vccd1 _08215_ sky130_fd_sc_hd__mux2_1
X_12332_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _05250_ vssd1 vssd1 vccd1 vccd1 _05518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15051_ _06033_ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__nand2_1
X_12263_ _04849_ _05398_ _05415_ _05432_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o32a_1
XFILLER_0_32_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _07165_ _07166_ _07171_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__nor3_1
X_11214_ net2855 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__clkbuf_1
X_12194_ net7733 net4952 _04845_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__mux2_1
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__clkbuf_4
X_18810_ net3940 _02954_ net4814 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11145_ net2513 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__clkbuf_1
Xoutput73 net143 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__buf_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18741_ _09739_ net4808 net8062 net3759 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__a31o_1
X_15953_ _08470_ _08484_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__and2b_1
X_11076_ net6659 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
X_14904_ net4508 _08034_ _08036_ net3757 net8240 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__o221a_1
XFILLER_0_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18672_ net4686 net4635 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__and2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _08858_ _08859_ _08895_ _08932_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__and4_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _01861_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ _07860_ _07804_ _07875_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__a21oi_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _01794_ _09403_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__nor2_1
X_11978_ rbzero.debug_overlay.vplaneY\[10\] _05135_ _05162_ _05166_ vssd1 vssd1 vccd1
+ vccd1 _05167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14766_ net7813 _07883_ _07885_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16505_ _08611_ net7818 vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10929_ net7488 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
X_13717_ _06702_ _06692_ _06758_ net555 vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__a2bb2o_1
X_17485_ _01723_ _01726_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__and2_1
X_14697_ net4703 vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_168_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19224_ net1030 _03123_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__nand2_2
X_16436_ _09525_ _09526_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__xnor2_1
X_13648_ _06814_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ net5468 _03144_ _03161_ _03160_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13579_ _06718_ _06741_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__or3_1
X_16367_ net3502 _08115_ _09457_ _09458_ _01633_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__o221a_1
Xhold6209 _04137_ vssd1 vssd1 vccd1 vccd1 net6736 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_53_i_clk clknet_4_11__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18106_ _02336_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__or2b_1
X_15318_ _08181_ _08366_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__nand2_2
XFILLER_0_83_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16298_ _09371_ _09389_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_4_11__f_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19086_ net7496 net5863 _03109_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5508 _04239_ vssd1 vssd1 vccd1 vccd1 net6035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5519 net3601 vssd1 vssd1 vccd1 vccd1 net6046 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18037_ _08366_ _10289_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__nor2_1
X_15249_ _08306_ _08328_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4807 net869 vssd1 vssd1 vccd1 vccd1 net5334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4818 _00854_ vssd1 vssd1 vccd1 vccd1 net5345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4829 net846 vssd1 vssd1 vccd1 vccd1 net5356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_i_clk clknet_4_13__leaf_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ net40 _03605_ _03122_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__o21a_2
XFILLER_0_158_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18939_ net1933 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21950_ net392 net2410 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20901_ clknet_leaf_37_i_clk net5430 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21881_ net323 net2724 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ net3976 _03992_ _04490_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20763_ net948 net5492 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19770__50 clknet_1_1__leaf__03509_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
X_20694_ _09727_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7400 net755 vssd1 vssd1 vccd1 vccd1 net7927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7411 net4352 vssd1 vssd1 vccd1 vccd1 net7938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7422 rbzero.wall_tracer.trackDistX\[-7\] vssd1 vssd1 vccd1 vccd1 net7949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7433 net4574 vssd1 vssd1 vccd1 vccd1 net7960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7444 rbzero.wall_tracer.trackDistY\[-6\] vssd1 vssd1 vccd1 vccd1 net7971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6710 rbzero.tex_r0\[36\] vssd1 vssd1 vccd1 vccd1 net7237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7455 net4507 vssd1 vssd1 vccd1 vccd1 net7982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6721 net2381 vssd1 vssd1 vccd1 vccd1 net7248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7466 rbzero.wall_tracer.trackDistY\[8\] vssd1 vssd1 vccd1 vccd1 net7993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6732 _04450_ vssd1 vssd1 vccd1 vccd1 net7259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7477 net4234 vssd1 vssd1 vccd1 vccd1 net8004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6743 net2744 vssd1 vssd1 vccd1 vccd1 net7270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7488 net8270 vssd1 vssd1 vccd1 vccd1 net8015 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6754 net2911 vssd1 vssd1 vccd1 vccd1 net7281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7499 _02802_ vssd1 vssd1 vccd1 vccd1 net8026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21315_ clknet_leaf_3_i_clk net5222 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6765 rbzero.tex_g1\[19\] vssd1 vssd1 vccd1 vccd1 net7292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6776 net957 vssd1 vssd1 vccd1 vccd1 net7303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6787 net2715 vssd1 vssd1 vccd1 vccd1 net7314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6798 rbzero.tex_r0\[37\] vssd1 vssd1 vccd1 vccd1 net7325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold350 net4418 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
X_21246_ clknet_leaf_8_i_clk net3400 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold361 _00961_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 net5277 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 net5309 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _01599_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
X_21177_ clknet_leaf_98_i_clk net1754 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_20128_ rbzero.debug_overlay.facingX\[-7\] _03711_ vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12950_ _06068_ _06061_ _06043_ net3960 _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__o221a_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__clkbuf_4
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 net6497 vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1061 net6588 vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11901_ _05085_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__nor2_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1072 net6159 vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 net4794 vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12881_ net4865 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__buf_8
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 net3896 vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _04852_ _05019_ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a21oi_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _07251_ _07342_ _07363_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__a21o_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _07708_ _07720_ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__nor2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _04933_ vssd1 vssd1 vccd1 vccd1 _04953_
+ sky130_fd_sc_hd__mux2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _04104_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__clkbuf_4
X_13502_ _06672_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17270_ _10288_ vssd1 vssd1 vccd1 vccd1 _10289_ sky130_fd_sc_hd__buf_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _07609_ _07652_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ net4132 _04863_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16221_ _09245_ _09313_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13433_ _06516_ _06539_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__or2_1
X_10645_ net7326 net7238 _04127_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16152_ _09243_ _09244_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ _06496_ _06528_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__a21oi_1
X_10576_ _04030_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__clkbuf_4
Xrebuffer6 net1674 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12315_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _05237_ vssd1 vssd1 vccd1 vccd1 _05501_
+ sky130_fd_sc_hd__mux2_1
X_15103_ _08196_ _08197_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__nand2_2
X_16083_ net8065 _08128_ _08491_ _09174_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__or4_4
X_13295_ _06403_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15034_ _08119_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__clkbuf_8
X_19911_ net2974 net7178 _03561_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_1
X_12246_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _04950_ vssd1 vssd1 vccd1 vccd1 _05433_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03511_ _03511_ vssd1 vssd1 vccd1 vccd1 clknet_0__03511_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19842_ net3111 net7542 _03528_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ _05363_ _05364_ _04938_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11128_ net1968 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
X_16985_ _09590_ _09588_ _09709_ vssd1 vssd1 vccd1 vccd1 _10007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ _02874_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__or2_1
X_11059_ net5636 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
X_15936_ net4405 _08128_ _08461_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18655_ net3619 _02789_ _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _08139_ net8042 _08959_ _08961_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__and4b_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _01846_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14818_ _07860_ _07830_ _07878_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _09751_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_130 vssd1 vssd1 vccd1 vccd1 ones[3] top_ew_algofoogle_130/LO sky130_fd_sc_hd__conb_1
X_15798_ _08854_ _08857_ _08891_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__and3_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_141 vssd1 vssd1 vccd1 vccd1 ones[14] top_ew_algofoogle_141/LO sky130_fd_sc_hd__conb_1
XFILLER_0_15_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17537_ _01677_ _01745_ _01776_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14749_ _07909_ _07911_ _07915_ net7824 net7806 vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__a221o_2
XFILLER_0_54_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20656__383 clknet_1_1__leaf__03870_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__inv_2
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17468_ _10311_ _10366_ _10364_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a21oi_1
X_20355__111 clknet_1_1__leaf__03841_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__inv_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19207_ net6862 _03183_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16419_ _08326_ _08403_ _09508_ vssd1 vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__o21ai_1
X_17399_ _10415_ _10414_ vssd1 vssd1 vccd1 vccd1 _10417_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6006 rbzero.tex_b0\[55\] vssd1 vssd1 vccd1 vccd1 net6533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6017 net1742 vssd1 vssd1 vccd1 vccd1 net6544 sky130_fd_sc_hd__dlygate4sd3_1
X_19138_ net4431 _03145_ net1239 _03149_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__o211a_1
Xhold6028 _04098_ vssd1 vssd1 vccd1 vccd1 net6555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6039 net1628 vssd1 vssd1 vccd1 vccd1 net6566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5305 net3716 vssd1 vssd1 vccd1 vccd1 net5832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5316 _00635_ vssd1 vssd1 vccd1 vccd1 net5843 sky130_fd_sc_hd__dlygate4sd3_1
X_19069_ net3940 _02472_ _03104_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5338 _00644_ vssd1 vssd1 vccd1 vccd1 net5865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5349 rbzero.spi_registers.spi_counter\[1\] vssd1 vssd1 vccd1 vccd1 net5876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4604 net722 vssd1 vssd1 vccd1 vccd1 net5131 sky130_fd_sc_hd__dlygate4sd3_1
X_21100_ clknet_leaf_7_i_clk net1446 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4615 _00812_ vssd1 vssd1 vccd1 vccd1 net5142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22080_ net522 net2776 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
Xhold4626 net785 vssd1 vssd1 vccd1 vccd1 net5153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4637 rbzero.spi_registers.texadd0\[18\] vssd1 vssd1 vccd1 vccd1 net5164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3903 net3531 vssd1 vssd1 vccd1 vccd1 net4430 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold4648 net809 vssd1 vssd1 vccd1 vccd1 net5175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3914 net5782 vssd1 vssd1 vccd1 vccd1 net4441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4659 _00788_ vssd1 vssd1 vccd1 vccd1 net5186 sky130_fd_sc_hd__dlygate4sd3_1
X_21031_ clknet_leaf_55_i_clk net4292 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3925 _00766_ vssd1 vssd1 vccd1 vccd1 net4452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3936 _03715_ vssd1 vssd1 vccd1 vccd1 net4463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3947 _01199_ vssd1 vssd1 vccd1 vccd1 net4474 sky130_fd_sc_hd__dlygate4sd3_1
X_19807__84 clknet_1_0__leaf__03512_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__inv_2
XFILLER_0_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3958 net3617 vssd1 vssd1 vccd1 vccd1 net4485 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3969 net3630 vssd1 vssd1 vccd1 vccd1 net4496 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21933_ net375 net2031 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21864_ net306 net1274 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20815_ net1028 net5480 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__nand2_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21795_ net237 net2151 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20746_ _03919_ _03920_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7241 net3372 vssd1 vssd1 vccd1 vccd1 net7768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7252 _09105_ vssd1 vssd1 vccd1 vccd1 net7779 sky130_fd_sc_hd__buf_2
XFILLER_0_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6540 net2327 vssd1 vssd1 vccd1 vccd1 net7067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7285 _06564_ vssd1 vssd1 vccd1 vccd1 net7812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6551 rbzero.tex_g1\[45\] vssd1 vssd1 vccd1 vccd1 net7078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7296 _06546_ vssd1 vssd1 vccd1 vccd1 net7823 sky130_fd_sc_hd__buf_1
Xhold6562 net2725 vssd1 vssd1 vccd1 vccd1 net7089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6573 rbzero.tex_b1\[57\] vssd1 vssd1 vccd1 vccd1 net7100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12100_ _05018_ _05287_ _05288_ _05203_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6584 net2023 vssd1 vssd1 vccd1 vccd1 net7111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6595 rbzero.tex_r1\[52\] vssd1 vssd1 vccd1 vccd1 net7122 sky130_fd_sc_hd__dlygate4sd3_1
X_13080_ net5428 _06242_ _06241_ _06253_ vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a22o_1
Xhold5850 rbzero.spi_registers.new_texadd\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net6377
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5861 net1405 vssd1 vssd1 vccd1 vccd1 net6388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5872 net1552 vssd1 vssd1 vccd1 vccd1 net6399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5883 rbzero.spi_registers.new_mapd\[0\] vssd1 vssd1 vccd1 vccd1 net6410 sky130_fd_sc_hd__dlygate4sd3_1
X_12031_ _04978_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__buf_4
Xhold5894 rbzero.spi_registers.new_texadd\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net6421
+ sky130_fd_sc_hd__dlygate4sd3_1
X_21229_ clknet_leaf_123_i_clk net3193 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold180 net5068 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold191 net5026 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_205_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _06058_ _09799_ _09801_ vssd1 vssd1 vccd1 vccd1 _09802_ sky130_fd_sc_hd__o21ai_1
X_13982_ _06729_ _06839_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__nand2_1
X_15721_ net8414 _08279_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__nor2_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ net3998 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__clkbuf_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _02585_ _02596_ _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a21o_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _08715_ _08723_ _08724_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__and3_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _06039_ _06028_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14603_ _07698_ _07730_ _07773_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__o21ai_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _04978_ vssd1 vssd1 vccd1 vccd1 _05005_
+ sky130_fd_sc_hd__mux2_1
X_18371_ _02549_ _02550_ _02556_ _04481_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _08240_ _08277_ _08278_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17322_ _10339_ _10340_ vssd1 vssd1 vccd1 vccd1 _10341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _04912_ vssd1 vssd1 vccd1 vccd1 _04936_
+ sky130_fd_sc_hd__mux2_1
X_14534_ _07033_ _07457_ _07703_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17253_ _10159_ _10160_ _10157_ vssd1 vssd1 vccd1 vccd1 _10272_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14465_ _07413_ _07194_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__nor2_1
X_11677_ _04858_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__nand2_1
X_16204_ net8041 _06122_ _08491_ _09296_ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__or4_2
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ net2817 net6172 _04116_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13416_ _06583_ _06586_ _06538_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__a21o_1
X_17184_ _10184_ _10203_ vssd1 vssd1 vccd1 vccd1 _10204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14396_ _07522_ _07525_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16135_ _09227_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13347_ _06389_ _06467_ _06433_ _06517_ _06424_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__a311o_1
XFILLER_0_109_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10559_ net2881 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16066_ _09158_ _09159_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__xnor2_1
X_13278_ _06353_ _06327_ _06404_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12229_ rbzero.tex_g1\[35\] rbzero.tex_g1\[34\] _04838_ vssd1 vssd1 vccd1 vccd1 _05416_
+ sky130_fd_sc_hd__mux2_1
X_15017_ _04476_ net3452 vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__nor2_1
Xhold2509 _03129_ vssd1 vssd1 vccd1 vccd1 net3036 sky130_fd_sc_hd__dlygate4sd3_1
X_19825_ net7554 net3045 _03517_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__mux2_1
Xhold1808 _01316_ vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 _04441_ vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16968_ _09988_ _09989_ vssd1 vssd1 vccd1 vccd1 _09990_ sky130_fd_sc_hd__xor2_2
X_18707_ _02824_ _02835_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a21o_1
X_15919_ _09012_ _09013_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__nand2_1
X_19687_ net1350 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__clkbuf_1
X_16899_ _09908_ _09920_ vssd1 vssd1 vccd1 vccd1 _09921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18638_ _02791_ _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ net3991 _09788_ _02734_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21580_ net214 net1199 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5102 rbzero.tex_r0\[3\] vssd1 vssd1 vccd1 vccd1 net5629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5113 rbzero.tex_g0\[1\] vssd1 vssd1 vccd1 vccd1 net5640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5124 net2824 vssd1 vssd1 vccd1 vccd1 net5651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5135 net5699 vssd1 vssd1 vccd1 vccd1 net5662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5146 net2306 vssd1 vssd1 vccd1 vccd1 net5673 sky130_fd_sc_hd__dlygate4sd3_1
X_22132_ clknet_leaf_52_i_clk net5741 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold4401 net593 vssd1 vssd1 vccd1 vccd1 net4928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5157 net2703 vssd1 vssd1 vccd1 vccd1 net5684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4412 gpout1.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5168 rbzero.tex_r1\[29\] vssd1 vssd1 vccd1 vccd1 net5695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4423 net609 vssd1 vssd1 vccd1 vccd1 net4950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4434 _00892_ vssd1 vssd1 vccd1 vccd1 net4961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5179 net1438 vssd1 vssd1 vccd1 vccd1 net5706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3700 net972 vssd1 vssd1 vccd1 vccd1 net4227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4445 net648 vssd1 vssd1 vccd1 vccd1 net4972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4456 rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 net4983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3711 net1121 vssd1 vssd1 vccd1 vccd1 net4238 sky130_fd_sc_hd__dlygate4sd3_1
X_22063_ net505 net2022 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold3722 net970 vssd1 vssd1 vccd1 vccd1 net4249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4467 net669 vssd1 vssd1 vccd1 vccd1 net4994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3733 _00495_ vssd1 vssd1 vccd1 vccd1 net4260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4478 net697 vssd1 vssd1 vccd1 vccd1 net5005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3744 net8146 vssd1 vssd1 vccd1 vccd1 net4271 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold4489 rbzero.spi_registers.texadd3\[0\] vssd1 vssd1 vccd1 vccd1 net5016 sky130_fd_sc_hd__dlygate4sd3_1
X_21014_ clknet_leaf_62_i_clk net4298 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3755 net1107 vssd1 vssd1 vccd1 vccd1 net4282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3766 rbzero.wall_tracer.visualWallDist\[-3\] vssd1 vssd1 vccd1 vccd1 net4293
+ sky130_fd_sc_hd__clkbuf_4
Xhold3777 rbzero.row_render.size\[5\] vssd1 vssd1 vccd1 vccd1 net4304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3788 net8158 vssd1 vssd1 vccd1 vccd1 net4315 sky130_fd_sc_hd__clkbuf_2
Xhold3799 net1063 vssd1 vssd1 vccd1 vccd1 net4326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21916_ net358 net1589 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21847_ net289 net2115 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11600_ net1008 net1233 net1046 net647 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ net18 vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21778_ clknet_leaf_8_i_clk net1787 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11531_ net1803 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20729_ _03904_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14250_ _07418_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ _06371_ _06301_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nor2_1
Xhold7060 net3543 vssd1 vssd1 vccd1 vccd1 net7587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7071 _03102_ vssd1 vssd1 vccd1 vccd1 net7598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _07350_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nor2_1
Xhold7082 net3648 vssd1 vssd1 vccd1 vccd1 net7609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11393_ _04576_ _04583_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__o21a_1
Xhold7093 rbzero.spi_registers.spi_buffer\[15\] vssd1 vssd1 vccd1 vccd1 net7620 sky130_fd_sc_hd__dlygate4sd3_1
X_20341__98 clknet_1_0__leaf__03840_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__inv_2
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6370 rbzero.tex_r1\[6\] vssd1 vssd1 vccd1 vccd1 net6897 sky130_fd_sc_hd__dlygate4sd3_1
X_13132_ _06268_ _06269_ _06300_ _06301_ _06302_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a311o_2
Xhold6381 net2159 vssd1 vssd1 vccd1 vccd1 net6908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6392 _04141_ vssd1 vssd1 vccd1 vccd1 net6919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17940_ _01794_ _10346_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5680 net1523 vssd1 vssd1 vccd1 vccd1 net6207 sky130_fd_sc_hd__dlygate4sd3_1
X_13063_ _06238_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__buf_2
Xhold5691 rbzero.tex_b1\[36\] vssd1 vssd1 vccd1 vccd1 net6218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12014_ net42 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__clkbuf_8
Xhold4990 rbzero.floor_leak\[4\] vssd1 vssd1 vccd1 vccd1 net5517 sky130_fd_sc_hd__dlygate4sd3_1
X_17871_ _02107_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19610_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__buf_2
XFILLER_0_206_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16822_ _09848_ net4508 net4649 vssd1 vssd1 vccd1 vccd1 _09849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19541_ net1623 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
X_16753_ _09768_ _09785_ _09786_ _09769_ net5328 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__a32o_1
X_13965_ _07132_ _07134_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__nand2_1
X_15704_ _08309_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__buf_4
X_12916_ net8034 vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__inv_4
X_19472_ net1725 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
X_16684_ _09736_ vssd1 vssd1 vccd1 vccd1 _09743_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13896_ _07040_ _07066_ _07064_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18423_ net3604 _02604_ _02537_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
X_15635_ _08661_ _08473_ _08630_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__or3_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__nor2_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20573__307 clknet_1_0__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__inv_2
XFILLER_0_69_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18354_ _02529_ _02530_ _02531_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__o21a_1
X_15566_ _08118_ _08164_ _08165_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__a21oi_4
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__and2_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17305_ _10322_ _10323_ vssd1 vssd1 vccd1 vccd1 _10324_ sky130_fd_sc_hd__xor2_2
XFILLER_0_138_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _07666_ _07686_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nor2_1
X_11729_ _04828_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18285_ net1632 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__clkbuf_1
X_15497_ _08587_ _08591_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ _10006_ _10008_ _10130_ _10255_ vssd1 vssd1 vccd1 vccd1 _10256_ sky130_fd_sc_hd__o31a_4
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _07242_ _07457_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__nor2_1
X_17167_ _08140_ _10186_ vssd1 vssd1 vccd1 vccd1 _10187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold905 net6429 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ _07535_ _07549_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__xor2_4
Xhold916 _01261_ vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold927 _03471_ vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ _09086_ _09099_ _09211_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__a21oi_2
Xhold938 net6449 vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _10117_ _10118_ vssd1 vssd1 vccd1 vccd1 _10119_ sky130_fd_sc_hd__and2b_1
Xhold949 _01264_ vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20467__212 clknet_1_1__leaf__03852_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__inv_2
Xhold3007 _02808_ vssd1 vssd1 vccd1 vccd1 net3534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16049_ _08207_ _08323_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3018 _03623_ vssd1 vssd1 vccd1 vccd1 net3545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3029 net7588 vssd1 vssd1 vccd1 vccd1 net3556 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_122_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2306 net7259 vssd1 vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2317 rbzero.tex_b1\[63\] vssd1 vssd1 vccd1 vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2328 _04433_ vssd1 vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 net3162 vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 net6759 vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1616 net7284 vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 _01561_ vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1638 net7114 vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 net7104 vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
X_19739_ net7656 net2310 net3824 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__and3b_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21701_ clknet_leaf_115_i_clk net4330 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21632_ clknet_leaf_129_i_clk net3075 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21563_ net197 net1899 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21494_ clknet_leaf_7_i_clk net1813 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_texadd\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4220 rbzero.debug_overlay.playerY\[1\] vssd1 vssd1 vccd1 vccd1 net4747 sky130_fd_sc_hd__dlygate4sd3_1
X_22115_ clknet_leaf_62_i_clk net5386 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
Xhold4231 net8266 vssd1 vssd1 vccd1 vccd1 net4758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4242 net3702 vssd1 vssd1 vccd1 vccd1 net4769 sky130_fd_sc_hd__clkbuf_2
Xhold4253 net5976 vssd1 vssd1 vccd1 vccd1 net4780 sky130_fd_sc_hd__buf_1
Xhold4264 _02618_ vssd1 vssd1 vccd1 vccd1 net4791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4275 rbzero.pov.ready_buffer\[12\] vssd1 vssd1 vccd1 vccd1 net4802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3530 net7561 vssd1 vssd1 vccd1 vccd1 net4057 sky130_fd_sc_hd__clkbuf_4
X_22046_ net488 net2949 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
Xhold3541 _05295_ vssd1 vssd1 vccd1 vccd1 net4068 sky130_fd_sc_hd__buf_4
Xhold4286 net3973 vssd1 vssd1 vccd1 vccd1 net4813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3552 net5967 vssd1 vssd1 vccd1 vccd1 net4079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4297 rbzero.pov.ready_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net4824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3563 net5950 vssd1 vssd1 vccd1 vccd1 net4090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3574 net5999 vssd1 vssd1 vccd1 vccd1 net4101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3585 _03799_ vssd1 vssd1 vccd1 vccd1 net4112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2840 net2628 vssd1 vssd1 vccd1 vccd1 net3367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2851 net7936 vssd1 vssd1 vccd1 vccd1 net3378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3596 _09719_ vssd1 vssd1 vccd1 vccd1 net4123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2862 net5914 vssd1 vssd1 vccd1 vccd1 net3389 sky130_fd_sc_hd__clkbuf_2
Xhold2873 _00733_ vssd1 vssd1 vccd1 vccd1 net3400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2884 net5834 vssd1 vssd1 vccd1 vccd1 net3411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2895 net4707 vssd1 vssd1 vccd1 vccd1 net3422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ net7473 net7194 _04298_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__mux2_1
X_13750_ net3513 _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__or2b_1
XFILLER_0_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12701_ _05862_ _05875_ _05877_ _05878_ net33 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ net7477 net3202 _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__mux2_1
X_13681_ _06713_ _06717_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__or2b_1
XFILLER_0_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ _08207_ _08509_ _08357_ vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ net4111 _05673_ net4071 net4092 _05802_ net24 vssd1 vssd1 vccd1 vccd1 _05811_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12563_ _05743_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
X_15351_ net8041 _08124_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14302_ _07033_ _07193_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__or2_1
X_11514_ net4091 net4138 _04661_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__or3_1
X_18070_ _02225_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ _08161_ net8414 _08368_ _08376_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__or4_2
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ net4111 _05673_ net4071 net4092 _05633_ net6 vssd1 vssd1 vccd1 vccd1 _05676_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17021_ _08661_ _09062_ vssd1 vssd1 vccd1 vccd1 _10042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14233_ _06914_ _07193_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11445_ rbzero.spi_registers.texadd1\[3\] _04548_ _04636_ vssd1 vssd1 vccd1 vccd1
+ _04637_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14164_ _07234_ _07235_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ rbzero.spi_registers.texadd3\[21\] rbzero.spi_registers.texadd1\[21\] rbzero.spi_registers.texadd0\[21\]
+ rbzero.spi_registers.texadd2\[21\] _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__inv_2
X_14095_ _07207_ _07248_ _07265_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__a21oi_1
X_18972_ net7467 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _01816_ _02066_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__nor2_1
X_13046_ _06187_ _06176_ _06165_ net3729 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__o2bb2a_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17854_ _02070_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16805_ net4547 net4583 vssd1 vssd1 vccd1 vccd1 _09833_ sky130_fd_sc_hd__nor2_1
X_17785_ _02022_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14997_ _08093_ net4164 vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19524_ net1701 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
X_16736_ net5666 _09769_ _09768_ _09772_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__a22o_1
X_13948_ _06841_ _06848_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__and2b_1
XFILLER_0_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19455_ net2098 _03335_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16667_ net4407 _09737_ _09740_ net7825 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a22o_1
X_13879_ _06703_ _06832_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__nor2_1
X_18406_ net3509 _05155_ _02587_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__nor4_2
X_15618_ _08666_ _08253_ _08254_ _08711_ _08712_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__a41o_1
XFILLER_0_201_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19386_ net6136 _03270_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__or2_1
X_16598_ _09684_ _09685_ _09687_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__nand3_1
X_18337_ net4883 _02508_ _09739_ net8255 _02525_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a221o_1
X_15549_ _08628_ _08641_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7807 rbzero.wall_tracer.stepDistY\[8\] vssd1 vssd1 vccd1 vccd1 net8334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7818 net4666 vssd1 vssd1 vccd1 vccd1 net8345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7829 rbzero.wall_tracer.trackDistX\[10\] vssd1 vssd1 vccd1 vccd1 net8356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18268_ net6393 net1396 _02477_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17219_ _10082_ _10113_ _10238_ vssd1 vssd1 vccd1 vccd1 _10239_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03857_ clknet_0__03857_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03857_
+ sky130_fd_sc_hd__clkbuf_16
X_18199_ _02419_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold702 net5481 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
X_20230_ net3680 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
Xhold713 net4432 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold724 _02987_ vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold735 _01158_ vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 net6501 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 net5521 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20161_ rbzero.debug_overlay.facingY\[-6\] net2485 _03723_ vssd1 vssd1 vccd1 vccd1
+ _03735_ sky130_fd_sc_hd__mux2_1
Xhold768 net6296 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold779 _01257_ vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2103 net5756 vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 net7054 vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_20092_ net3326 _03660_ net4902 _03679_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__o211a_1
Xhold2125 _04222_ vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2136 _01477_ vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2147 _04414_ vssd1 vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1402 net7024 vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2158 net7215 vssd1 vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _01559_ vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1424 _01310_ vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2169 _01296_ vssd1 vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 net6809 vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 net6654 vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1457 _01066_ vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1468 _04181_ vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 net5553 vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20994_ clknet_leaf_112_i_clk net5951 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20521__261 clknet_1_0__leaf__03857_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__inv_2
XFILLER_0_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21615_ clknet_leaf_97_i_clk net3079 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21546_ net180 net2913 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21477_ clknet_leaf_18_i_clk net4846 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_texadd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11230_ net6780 net2170 _04434_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ net7377 net3117 _04401_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4050 _08053_ vssd1 vssd1 vccd1 vccd1 net4577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4061 net7961 vssd1 vssd1 vccd1 vccd1 net4588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4072 _02755_ vssd1 vssd1 vccd1 vccd1 net4599 sky130_fd_sc_hd__dlygate4sd3_1
X_11092_ net6184 net7407 _04364_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__mux2_1
Xhold4083 net3831 vssd1 vssd1 vccd1 vccd1 net4610 sky130_fd_sc_hd__clkbuf_2
Xhold4094 net8336 vssd1 vssd1 vccd1 vccd1 net4621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3360 net4919 vssd1 vssd1 vccd1 vccd1 net3887 sky130_fd_sc_hd__dlygate4sd3_1
X_22029_ net471 net2612 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3371 _02470_ vssd1 vssd1 vccd1 vccd1 net3898 sky130_fd_sc_hd__dlygate4sd3_1
X_14920_ net8071 _08047_ _08043_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__o21a_1
Xhold3382 net5876 vssd1 vssd1 vccd1 vccd1 net3909 sky130_fd_sc_hd__clkbuf_2
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3393 _00475_ vssd1 vssd1 vccd1 vccd1 net3920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20604__336 clknet_1_1__leaf__03865_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__inv_2
XFILLER_0_199_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2670 _00674_ vssd1 vssd1 vccd1 vccd1 net3197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _01155_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2681 _03027_ vssd1 vssd1 vccd1 vccd1 net3208 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net7811 _07995_ _07934_ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__o21ai_1
Xhold73 net4935 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2692 _00924_ vssd1 vssd1 vccd1 vccd1 net3219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 net5046 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 net4965 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ net568 _06708_ _06970_ _06971_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__a41o_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _09272_ _10220_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nor2_1
Xhold1980 _03521_ vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1991 net7274 vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_14782_ _07940_ _07942_ _07946_ net7824 net4704 vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__a221o_2
X_11994_ net4161 vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_9__f_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16521_ _09609_ _09610_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__nor2_1
X_13733_ _06882_ _06903_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__and2_1
X_10945_ net7361 net6107 _04287_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19240_ net6599 _03203_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__or2_1
X_16452_ _08030_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__inv_2
X_13664_ _06759_ _06800_ _06756_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__a21boi_1
X_10876_ net7357 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15403_ _08496_ _08497_ _08495_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12615_ reg_gpout\[2\] clknet_1_1__leaf__05794_ net45 vssd1 vssd1 vccd1 vccd1 _05795_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19171_ net6285 _03170_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__or2_1
X_16383_ _09470_ _09473_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__xnor2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _06762_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__nand2_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18122_ net3847 net4415 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__nand2_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ net4401 _06121_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ _04648_ net4133 _04461_ net4089 net12 _05691_ vssd1 vssd1 vccd1 vccd1 _05727_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18053_ _02192_ _02195_ _02193_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15265_ _07968_ _07975_ _07981_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12477_ net8 _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17004_ _09951_ _09933_ vssd1 vssd1 vccd1 vccd1 _10025_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _07328_ _07386_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__and2_1
X_11428_ _04530_ _04523_ _04528_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__nand3_1
X_15196_ net8263 _08119_ _06120_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ _07313_ _07316_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__nor2_1
X_11359_ rbzero.spi_registers.texadd2\[14\] _04506_ _04507_ _04550_ vssd1 vssd1 vccd1
+ vccd1 _04551_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14078_ net580 _07206_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__nand2_1
X_18955_ net1907 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13029_ net3785 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__inv_2
X_17906_ _02141_ _02143_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__xor2_1
X_18886_ net2080 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17837_ _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nand2_1
X_20579__313 clknet_1_1__leaf__03863_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__inv_2
XFILLER_0_179_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer16 net542 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_1
Xrebuffer27 _06502_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_1
X_17768_ _01818_ _02005_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__or2_1
Xrebuffer38 _08439_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__dlygate4sd3_1
Xrebuffer49 _06643_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19507_ net4016 net6578 _03365_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__mux2_1
X_16719_ net3965 _08194_ vssd1 vssd1 vccd1 vccd1 _09757_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ _01937_ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__and2b_1
XFILLER_0_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19438_ net1625 net3519 _03141_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ net6257 _03284_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7604 rbzero.traced_texa\[-6\] vssd1 vssd1 vccd1 vccd1 net8131 sky130_fd_sc_hd__dlygate4sd3_1
X_21400_ clknet_leaf_41_i_clk net4966 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7615 _00506_ vssd1 vssd1 vccd1 vccd1 net8142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7626 rbzero.row_render.texu\[2\] vssd1 vssd1 vccd1 vccd1 net8153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7637 rbzero.map_overlay.i_mapdx\[1\] vssd1 vssd1 vccd1 vccd1 net8164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6903 rbzero.tex_g0\[61\] vssd1 vssd1 vccd1 vccd1 net7430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7648 rbzero.map_overlay.i_mapdx\[3\] vssd1 vssd1 vccd1 vccd1 net8175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6914 net2993 vssd1 vssd1 vccd1 vccd1 net7441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7659 _03740_ vssd1 vssd1 vccd1 vccd1 net8186 sky130_fd_sc_hd__dlygate4sd3_1
X_21331_ clknet_leaf_8_i_clk net5426 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6925 rbzero.pov.spi_buffer\[46\] vssd1 vssd1 vccd1 vccd1 net7452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6936 net3132 vssd1 vssd1 vccd1 vccd1 net7463 sky130_fd_sc_hd__dlygate4sd3_1
X_20551__287 clknet_1_1__leaf__03861_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__inv_2
XFILLER_0_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6947 rbzero.spi_registers.new_mapd\[7\] vssd1 vssd1 vccd1 vccd1 net7474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6958 rbzero.tex_g0\[31\] vssd1 vssd1 vccd1 vccd1 net7485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6969 net2182 vssd1 vssd1 vccd1 vccd1 net7496 sky130_fd_sc_hd__dlygate4sd3_1
X_21262_ clknet_leaf_122_i_clk net1729 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold510 net5425 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold521 net8131 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold532 net7551 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold543 net6185 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
X_20213_ _05164_ _03744_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__or2_1
Xhold554 net6165 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
X_21193_ clknet_leaf_124_i_clk net1246 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold565 net6121 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold576 net7482 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 net4474 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 net5689 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
X_20144_ net3719 net3131 _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ _08232_ _03610_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__nor2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _03376_ vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 net5629 vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1232 net6851 vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1243 net6696 vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1254 _00959_ vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
X_20445__192 clknet_1_1__leaf__03850_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__inv_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1265 _08064_ vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1276 net8152 vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 net7311 vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _04436_ vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ clknet_leaf_42_i_clk net4014 vssd1 vssd1 vccd1 vccd1 rbzero.wall_hot\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ net6820 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ net2391 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12400_ _05583_ _05584_ _05204_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13380_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__buf_6
X_10592_ net2304 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12331_ _04943_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__buf_4
X_21529_ clknet_leaf_124_i_clk net3706 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12262_ _04991_ _05440_ _05448_ _04821_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a31o_1
X_15050_ net3489 net3417 vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ net7301 net7297 _04423_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14001_ _07165_ _07166_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__o21a_1
X_12193_ _05380_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
XFILLER_0_43_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11144_ net7242 net6534 _04390_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__mux2_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 o_reset sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20528__267 clknet_1_0__leaf__03858_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__inv_2
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18740_ _02889_ _02890_ rbzero.wall_tracer.rayAddendY\[5\] _09735_ vssd1 vssd1 vccd1
+ vccd1 _02891_ sky130_fd_sc_hd__a2bb2o_1
X_11075_ net1660 net6657 _04353_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__mux2_1
X_15952_ _09024_ _09046_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3190 net5833 vssd1 vssd1 vccd1 vccd1 net3717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14903_ net4236 _08037_ _08043_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__o21a_1
X_18671_ net4686 net4635 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__nor2_2
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08859_ _08936_ _08977_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__and3_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _08661_ _09612_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _07992_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19756__37 clknet_1_0__leaf__03508_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _09262_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__buf_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _06505_ net7839 vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__nor2_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ rbzero.debug_overlay.vplaneY\[-7\] _05090_ _05163_ _05165_ vssd1 vssd1 vccd1
+ vccd1 _05166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ net8034 _08181_ _08129_ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__and3_1
X_13716_ _06673_ _06755_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__nor2_1
X_17484_ _10267_ _10256_ _10377_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__o31a_4
X_10928_ net7486 net3246 _04276_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ _07843_ _07858_ _07866_ net7839 vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__a211o_1
X_19223_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16435_ _08880_ _09165_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _06816_ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__xor2_2
X_10859_ net2504 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ net1292 _03146_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ net7779 _09456_ net3454 vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__a21o_1
X_13578_ _06747_ _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18105_ net3787 net4539 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15317_ _08401_ _08402_ _08403_ _08411_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19085_ net6794 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__clkbuf_1
X_12529_ _05707_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand2_1
X_16297_ _09372_ _09388_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5509 net631 vssd1 vssd1 vccd1 vccd1 net6036 sky130_fd_sc_hd__dlygate4sd3_1
X_18036_ _02212_ _02213_ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__o21a_1
X_15248_ _08294_ _08317_ vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4808 rbzero.spi_registers.texadd0\[20\] vssd1 vssd1 vccd1 vccd1 net5335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4819 net1001 vssd1 vssd1 vccd1 vccd1 net5346 sky130_fd_sc_hd__dlygate4sd3_1
X_15179_ _06009_ _06340_ net4180 vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19987_ net4997 _03484_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__and2_2
XFILLER_0_158_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18938_ net3320 net6878 _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
.ends

