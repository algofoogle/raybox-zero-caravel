* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd2_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_la_invalid i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_outs_enb i_reg_sclk i_reset_lock_a i_reset_lock_b i_spare_0 i_spare_1 i_test_uc2
+ i_test_wci i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3] i_vec_csb i_vec_mosi
+ i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_gpout[3] o_gpout[4] o_gpout[5] o_hsync
+ o_reset o_rgb[10] o_rgb[11] o_rgb[12] o_rgb[13] o_rgb[14] o_rgb[15] o_rgb[18] o_rgb[19]
+ o_rgb[20] o_rgb[21] o_rgb[22] o_rgb[23] o_rgb[6] o_rgb[7] o_tex_csb o_tex_oeb0 o_tex_out0
+ o_tex_sclk o_vsync ones[12] ones[13] ones[14] ones[15] ones[1] ones[2] ones[3] ones[4]
+ ones[5] ones[7] ones[8] ones[9] vccd1 vssd1 zeros[10] zeros[12] zeros[13] zeros[14]
+ zeros[15] zeros[2] zeros[3] zeros[4] zeros[5] zeros[6] zeros[7] zeros[8] zeros[9]
+ o_rgb[17] ones[11] o_rgb[16] ones[0] ones[10] ones[6] o_rgb[9] o_rgb[8] o_rgb[5]
+ o_rgb[4] o_rgb[3] o_rgb[2] o_rgb[1] o_rgb[0] zeros[1] zeros[0] zeros[11]
XFILLER_0_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18869_ rbzero.wall_tracer.rayAddendY\[2\] rbzero.wall_tracer.rayAddendY\[1\] net4708
+ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21880_ clknet_leaf_99_i_clk net1178 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22432_ clknet_leaf_40_i_clk net4544 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6700 rbzero.tex_b1\[40\] vssd1 vssd1 vccd1 vccd1 net7224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22363_ net495 net1349 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold6711 net2695 vssd1 vssd1 vccd1 vccd1 net7235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6722 rbzero.tex_r0\[6\] vssd1 vssd1 vccd1 vccd1 net7246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6733 rbzero.tex_b0\[25\] vssd1 vssd1 vccd1 vccd1 net7257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6744 net2858 vssd1 vssd1 vccd1 vccd1 net7268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21314_ clknet_leaf_73_i_clk net4276 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6755 rbzero.tex_r1\[19\] vssd1 vssd1 vccd1 vccd1 net7279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6766 net2845 vssd1 vssd1 vccd1 vccd1 net7290 sky130_fd_sc_hd__dlygate4sd3_1
X_22294_ net426 net2387 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold6777 rbzero.tex_g0\[38\] vssd1 vssd1 vccd1 vccd1 net7301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6788 _03304_ vssd1 vssd1 vccd1 vccd1 net7312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6799 _03089_ vssd1 vssd1 vccd1 vccd1 net7323 sky130_fd_sc_hd__dlygate4sd3_1
X_21245_ clknet_leaf_53_i_clk net3541 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold340 net4906 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold351 net5129 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold362 net5225 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold373 net5148 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 net4790 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
X_21176_ net4142 _04140_ _04141_ _09908_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold395 net5294 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20127_ net3590 _03676_ _03682_ _03683_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20058_ _03440_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__clkbuf_4
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 _03414_ vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 net6056 vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ _04986_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__buf_4
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1062 net5715 vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1073 net6247 vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ net3 _06007_ _06008_ clknet_leaf_67_i_clk vssd1 vssd1 vccd1 vccd1 _06038_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_198_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1084 net3950 vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__buf_4
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 net5751 vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _04984_ _04990_ _04996_ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__o211a_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _07660_ _07663_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__xnor2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ net2776 _04931_ _04929_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a21oi_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _06565_ _06587_ _06629_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__and3_1
X_10713_ net7171 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__clkbuf_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _07616_ _07630_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__nor2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ net2043 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__inv_2
X_16220_ _09294_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ _06572_ _06573_ _06576_ _06541_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__a31o_1
X_10644_ net6908 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16151_ _08633_ _09224_ _09225_ _08610_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ _06511_ _06513_ _06429_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer7 net530 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ net3047 net3233 _08219_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__mux2_1
X_12314_ _05019_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__or2_1
X_16082_ _08325_ net7444 _09154_ _09151_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__or4b_1
X_13294_ _06438_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19910_ net4355 _03530_ net2912 _03496_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__o211a_1
X_15033_ net3064 _08168_ _08026_ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__mux2_1
X_12245_ rbzero.debug_overlay.facingX\[-4\] _05383_ _05384_ rbzero.debug_overlay.facingX\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19841_ net4335 _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__nor2_1
X_12176_ _04605_ net3910 _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ net6391 net1750 _04437_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__mux2_1
X_16984_ net4507 net4579 vssd1 vssd1 vccd1 vccd1 _09996_ sky130_fd_sc_hd__or2_1
X_19772_ net6660 _03429_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15935_ _08987_ _08981_ _08986_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__nand3_1
X_11058_ net7143 net7095 _04404_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18723_ net4587 _05401_ _02700_ _08246_ _02676_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__o311a_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20721__154 clknet_1_0__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__inv_2
X_18654_ net4696 net7608 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__and2_1
X_15866_ _08837_ _08885_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__or2_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _01655_ _01656_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nand2_1
X_14817_ _07742_ _07792_ _07794_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18585_ _02594_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_120 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_120/HI zeros[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_204_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15797_ _08471_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__buf_4
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_131 vssd1 vssd1 vccd1 vccd1 ones[7] top_ew_algofoogle_131/LO sky130_fd_sc_hd__conb_1
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17536_ _09582_ _09861_ vssd1 vssd1 vccd1 vccd1 _10535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14748_ _07892_ _07898_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17467_ _10217_ _10445_ vssd1 vssd1 vccd1 vccd1 _10466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14679_ _07818_ _07829_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16418_ _09371_ _09490_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__xor2_2
X_19206_ net5151 _03078_ _03102_ _03096_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17398_ _10385_ _10397_ vssd1 vssd1 vccd1 vccd1 _10398_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19137_ _02992_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__clkbuf_4
X_16349_ _09309_ _09313_ _09307_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__a21o_1
Xhold6007 net1430 vssd1 vssd1 vccd1 vccd1 net6531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6018 rbzero.tex_g0\[57\] vssd1 vssd1 vccd1 vccd1 net6542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6029 net1513 vssd1 vssd1 vccd1 vccd1 net6553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5306 net2473 vssd1 vssd1 vccd1 vccd1 net5830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5317 rbzero.tex_b1\[2\] vssd1 vssd1 vccd1 vccd1 net5841 sky130_fd_sc_hd__dlygate4sd3_1
X_19068_ net6058 _03009_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5328 net2194 vssd1 vssd1 vccd1 vccd1 net5852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5339 _00792_ vssd1 vssd1 vccd1 vccd1 net5863 sky130_fd_sc_hd__dlygate4sd3_1
X_18019_ _01967_ _01969_ _01965_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4605 _00712_ vssd1 vssd1 vccd1 vccd1 net5129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4616 net861 vssd1 vssd1 vccd1 vccd1 net5140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4627 net987 vssd1 vssd1 vccd1 vccd1 net5151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4638 _00872_ vssd1 vssd1 vccd1 vccd1 net5162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21030_ net5334 _03519_ _04014_ _04032_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3904 net7528 vssd1 vssd1 vccd1 vccd1 net4428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4649 _00716_ vssd1 vssd1 vccd1 vccd1 net5173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3915 _02753_ vssd1 vssd1 vccd1 vccd1 net4439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3926 net7806 vssd1 vssd1 vccd1 vccd1 net4450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3937 _01024_ vssd1 vssd1 vccd1 vccd1 net4461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3948 net7819 vssd1 vssd1 vccd1 vccd1 net4472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3959 net3321 vssd1 vssd1 vccd1 vccd1 net4483 sky130_fd_sc_hd__clkbuf_2
X_21932_ clknet_leaf_8_i_clk net4842 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_20696__131 clknet_1_1__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__inv_2
XFILLER_0_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21863_ clknet_leaf_94_i_clk net3331 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21794_ clknet_leaf_11_i_clk net4221 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20338__71 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
XFILLER_0_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7220 net4422 vssd1 vssd1 vccd1 vccd1 net7744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20353__85 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__inv_2
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22415_ net143 net2264 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7242 _08427_ vssd1 vssd1 vccd1 vccd1 net7766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7253 _08389_ vssd1 vssd1 vccd1 vccd1 net7777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7264 net4385 vssd1 vssd1 vccd1 vccd1 net7788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6530 net2185 vssd1 vssd1 vccd1 vccd1 net7054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7275 _01978_ vssd1 vssd1 vccd1 vccd1 net7799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6541 rbzero.tex_r0\[5\] vssd1 vssd1 vccd1 vccd1 net7065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7286 _08369_ vssd1 vssd1 vccd1 vccd1 net7810 sky130_fd_sc_hd__dlygate4sd3_1
X_22346_ net478 net2507 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6552 _04330_ vssd1 vssd1 vccd1 vccd1 net7076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6563 net2415 vssd1 vssd1 vccd1 vccd1 net7087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6574 rbzero.tex_g0\[56\] vssd1 vssd1 vccd1 vccd1 net7098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6585 net2638 vssd1 vssd1 vccd1 vccd1 net7109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5840 rbzero.pov.mosi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5851 net1088 vssd1 vssd1 vccd1 vccd1 net6375 sky130_fd_sc_hd__dlygate4sd3_1
X_22277_ net409 net2634 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
Xhold6596 rbzero.tex_r0\[58\] vssd1 vssd1 vccd1 vccd1 net7120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5862 rbzero.tex_b1\[46\] vssd1 vssd1 vccd1 vccd1 net6386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5873 net1149 vssd1 vssd1 vccd1 vccd1 net6397 sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ net4001 net4972 net4059 vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5884 _04278_ vssd1 vssd1 vccd1 vccd1 net6408 sky130_fd_sc_hd__dlygate4sd3_1
X_21228_ clknet_leaf_57_i_clk _00397_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5895 net1179 vssd1 vssd1 vccd1 vccd1 net6419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold170 net4108 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold181 net3421 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 net4659 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
X_21159_ _04136_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20779__206 clknet_1_0__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__inv_2
X_13981_ _06781_ _06869_ _07129_ _07130_ _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__a41o_1
XFILLER_0_176_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15720_ _08794_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_52_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ net38 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__inv_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _08331_ _08454_ _08699_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__or3_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ net4060 _06012_ _06008_ _05194_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__a221o_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _07751_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__nand2_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__clkbuf_4
X_18370_ net3394 _02398_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__nand2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _08542_ _08626_ _08646_ _08645_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__or4b_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12794_ net26 _05949_ _05951_ _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a22o_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_67_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17321_ _10320_ _10321_ vssd1 vssd1 vccd1 vccd1 _10322_ sky130_fd_sc_hd__xor2_2
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _07668_ _07682_ _07683_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11745_ net1060 net1915 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__or2_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _10220_ _10252_ vssd1 vssd1 vccd1 vccd1 _10253_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_0__03990_ _03990_ vssd1 vssd1 vccd1 vccd1 clknet_0__03990_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14464_ _07595_ _07614_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ net4105 vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16203_ _09276_ net2943 vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13415_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17183_ _10182_ _10183_ _10161_ vssd1 vssd1 vccd1 vccd1 _10185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10627_ net2821 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14395_ _07525_ _07526_ _07545_ _07543_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _08449_ _08424_ _08550_ _08565_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__or4_1
X_13346_ _06455_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16065_ _09138_ _09139_ _08517_ _08874_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__or4_1
X_13277_ _06425_ _06427_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _06428_
+ sky130_fd_sc_hd__mux2_4
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15016_ _08031_ _08128_ _08141_ _08111_ net7458 net7478 vssd1 vssd1 vccd1 vccd1 _08154_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12228_ net3807 _05383_ _05384_ _05396_ _04889_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19824_ _02967_ net3926 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__and2_1
X_12159_ net4052 net4071 vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1809 _01143_ vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19755_ net3151 net4327 net3075 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__or3b_1
X_16967_ net5746 _09966_ _09965_ _09981_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a22o_1
X_18706_ _02696_ _02700_ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15918_ _08989_ _08992_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__and2_1
X_16898_ net839 _09937_ _09938_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1
+ vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
X_19686_ net3109 _03374_ net1730 _03384_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15849_ _08915_ _08922_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__or2b_1
X_18637_ _02637_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__buf_2
XFILLER_0_204_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18568_ net4690 rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _02582_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_176_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17519_ _08717_ _09477_ vssd1 vssd1 vccd1 vccd1 _10518_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18499_ net1296 net3374 _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20530_ net1018 net3800 _03889_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20461_ _03836_ net3783 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22200_ net332 net1814 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
X_20392_ net3587 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__clkbuf_1
Xhold5103 _01073_ vssd1 vssd1 vccd1 vccd1 net5627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5114 rbzero.spi_registers.texadd0\[5\] vssd1 vssd1 vccd1 vccd1 net5638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5125 net1320 vssd1 vssd1 vccd1 vccd1 net5649 sky130_fd_sc_hd__dlygate4sd3_1
X_22131_ net263 net2208 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5136 net1391 vssd1 vssd1 vccd1 vccd1 net5660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4402 net3461 vssd1 vssd1 vccd1 vccd1 net4926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5147 rbzero.pov.spi_buffer\[36\] vssd1 vssd1 vccd1 vccd1 net5671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4413 _04088_ vssd1 vssd1 vccd1 vccd1 net4937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5158 _00725_ vssd1 vssd1 vccd1 vccd1 net5682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5169 rbzero.pov.spi_buffer\[51\] vssd1 vssd1 vccd1 vccd1 net5693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4424 _00000_ vssd1 vssd1 vccd1 vccd1 net4948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4435 net662 vssd1 vssd1 vccd1 vccd1 net4959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4446 net691 vssd1 vssd1 vccd1 vccd1 net4970 sky130_fd_sc_hd__dlygate4sd3_1
X_22062_ clknet_leaf_7_i_clk net3649 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3701 _00893_ vssd1 vssd1 vccd1 vccd1 net4225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3712 _03410_ vssd1 vssd1 vccd1 vccd1 net4236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4457 net776 vssd1 vssd1 vccd1 vccd1 net4981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4468 _00870_ vssd1 vssd1 vccd1 vccd1 net4992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3723 rbzero.spi_registers.texadd0\[13\] vssd1 vssd1 vccd1 vccd1 net4247 sky130_fd_sc_hd__dlygate4sd3_1
X_21013_ _09920_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__clkbuf_4
Xhold4479 net771 vssd1 vssd1 vccd1 vccd1 net5003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3734 _03409_ vssd1 vssd1 vccd1 vccd1 net4258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3745 _00764_ vssd1 vssd1 vccd1 vccd1 net4269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3756 net7670 vssd1 vssd1 vccd1 vccd1 net4280 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3767 net7675 vssd1 vssd1 vccd1 vccd1 net4291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3778 net2947 vssd1 vssd1 vccd1 vccd1 net4302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3789 net1304 vssd1 vssd1 vccd1 vccd1 net4313 sky130_fd_sc_hd__dlygate4sd3_1
X_21915_ clknet_leaf_92_i_clk net1240 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21846_ clknet_leaf_82_i_clk net1367 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21777_ clknet_leaf_20_i_clk net2232 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ rbzero.spi_registers.texadd3\[22\] _04693_ _04692_ vssd1 vssd1 vccd1 vccd1
+ _04702_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_81_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ _04634_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlymetal6s2s_1
X_20750__180 clknet_1_0__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__inv_2
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ net2705 _06221_ _06354_ net2043 _06355_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__a221o_1
Xhold7061 _02581_ vssd1 vssd1 vccd1 vccd1 net7585 sky130_fd_sc_hd__dlygate4sd3_1
X_11392_ net6734 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
Xhold7072 _10054_ vssd1 vssd1 vccd1 vccd1 net7596 sky130_fd_sc_hd__dlygate4sd3_1
X_14180_ _07281_ _07330_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__xnor2_1
Xhold6360 net2140 vssd1 vssd1 vccd1 vccd1 net6884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6371 _04362_ vssd1 vssd1 vccd1 vccd1 net6895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13131_ net3493 vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__inv_2
X_22329_ net461 net2761 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6382 net2469 vssd1 vssd1 vccd1 vccd1 net6906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6393 _04317_ vssd1 vssd1 vccd1 vccd1 net6917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5670 rbzero.spi_registers.buf_texadd2\[7\] vssd1 vssd1 vccd1 vccd1 net6194 sky130_fd_sc_hd__dlygate4sd3_1
X_13062_ net2774 _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__nor2_1
Xhold5681 _00420_ vssd1 vssd1 vccd1 vccd1 net6205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5692 rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 net6216 sky130_fd_sc_hd__dlygate4sd3_1
X_12013_ net1524 _04998_ _04982_ rbzero.floor_leak\[1\] _05182_ vssd1 vssd1 vccd1
+ vccd1 _05183_ sky130_fd_sc_hd__a221o_1
X_17870_ _01918_ _01919_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__and2_1
Xhold4980 net1164 vssd1 vssd1 vccd1 vccd1 net5504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4991 net1114 vssd1 vssd1 vccd1 vccd1 net5515 sky130_fd_sc_hd__dlygate4sd3_1
X_16821_ _09887_ _09888_ _09890_ vssd1 vssd1 vccd1 vccd1 _09891_ sky130_fd_sc_hd__nand3_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16752_ _09820_ _09821_ vssd1 vssd1 vccd1 vccd1 _09822_ sky130_fd_sc_hd__nor2_1
X_19540_ net3864 net1571 _03298_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
X_13964_ _06865_ net541 vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__nor2_1
X_15703_ _08463_ _08508_ _08507_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__a21oi_2
X_12915_ net34 _06071_ _06065_ net43 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__a2bb2o_1
X_16683_ _09751_ _09753_ vssd1 vssd1 vccd1 vccd1 _09754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19471_ _02492_ _03238_ net3076 net6559 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__a31o_1
XFILLER_0_159_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13895_ _06941_ _06940_ _06939_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15634_ _08326_ _08708_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__nor2_1
X_18422_ _02450_ net4483 _02411_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ net4095 _05446_ net28 vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _02383_ _02384_ _02385_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15565_ _08624_ _08635_ _08627_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__a21o_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833__255 clknet_1_1__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__inv_2
X_12777_ net6355 _05894_ _05934_ net56 vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a22o_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _10177_ _10179_ _10303_ vssd1 vssd1 vccd1 vccd1 _10305_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14516_ _07651_ _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__xor2_4
X_20317__52 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_0_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ net4345 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__inv_2
X_18284_ _02166_ _02169_ _02252_ _02269_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a311oi_1
X_15496_ _08551_ _08562_ _08569_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17235_ _10130_ _09251_ vssd1 vssd1 vccd1 vccd1 _10236_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14447_ _07533_ _07535_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__nand2_2
X_11659_ net4001 _04827_ net3996 _04759_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a22o_1
X_20332__66 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
X_17166_ _06211_ _09870_ _10167_ vssd1 vssd1 vccd1 vccd1 _10168_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_25_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14378_ _07474_ _07354_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold906 net6530 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16117_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__xnor2_1
Xhold917 net5697 vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ net7770 _06430_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__nor2_1
Xhold928 net6267 vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ _09666_ _09133_ vssd1 vssd1 vccd1 vccd1 _10099_ sky130_fd_sc_hd__and2b_1
Xhold939 _01169_ vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _09074_ _09122_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3008 _03871_ vssd1 vssd1 vccd1 vccd1 net3532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3019 net3605 vssd1 vssd1 vccd1 vccd1 net3543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2307 _04341_ vssd1 vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2318 net3946 vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__buf_2
Xhold2329 _01484_ vssd1 vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1606 _01355_ vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
X_19807_ net6037 _03428_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__or2_1
Xhold1617 net5815 vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 net2517 vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_17999_ _02040_ _02047_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__xnor2_1
Xhold1639 net6921 vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19738_ net1784 _03408_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19669_ net5838 _03374_ net3012 _03371_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21700_ clknet_leaf_101_i_clk net5063 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21631_ clknet_leaf_19_i_clk net5293 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21562_ clknet_leaf_17_i_clk net5308 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20513_ net3715 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21493_ clknet_leaf_15_i_clk net2865 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20444_ net3743 net3843 _03823_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20375_ _08275_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4210 net3122 vssd1 vssd1 vccd1 vccd1 net4734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4221 _01607_ vssd1 vssd1 vccd1 vccd1 net4745 sky130_fd_sc_hd__dlygate4sd3_1
X_22114_ net246 net1802 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold4232 net2000 vssd1 vssd1 vccd1 vccd1 net4756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4243 _02664_ vssd1 vssd1 vccd1 vccd1 net4767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4254 net2834 vssd1 vssd1 vccd1 vccd1 net4778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4265 net3007 vssd1 vssd1 vccd1 vccd1 net4789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3520 _05202_ vssd1 vssd1 vccd1 vccd1 net4044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4276 _02759_ vssd1 vssd1 vccd1 vccd1 net4800 sky130_fd_sc_hd__dlygate4sd3_1
X_22045_ clknet_leaf_92_i_clk net3533 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3531 _09926_ vssd1 vssd1 vccd1 vccd1 net4055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3542 _05615_ vssd1 vssd1 vccd1 vccd1 net4066 sky130_fd_sc_hd__clkbuf_4
Xhold4287 _02690_ vssd1 vssd1 vccd1 vccd1 net4811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3553 _05187_ vssd1 vssd1 vccd1 vccd1 net4077 sky130_fd_sc_hd__clkbuf_4
Xhold4298 _06199_ vssd1 vssd1 vccd1 vccd1 net4822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3564 _08293_ vssd1 vssd1 vccd1 vccd1 net4088 sky130_fd_sc_hd__clkbuf_4
Xhold2830 _03829_ vssd1 vssd1 vccd1 vccd1 net3354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3575 net4058 vssd1 vssd1 vccd1 vccd1 net4099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3586 net7482 vssd1 vssd1 vccd1 vccd1 net4110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2841 net2911 vssd1 vssd1 vccd1 vccd1 net3365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 _02984_ vssd1 vssd1 vccd1 vccd1 net3376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3597 net7623 vssd1 vssd1 vccd1 vccd1 net4121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2863 rbzero.pov.ready_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net3387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2874 _10060_ vssd1 vssd1 vccd1 vccd1 net3398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2885 net6101 vssd1 vssd1 vccd1 vccd1 net3409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2896 net4529 vssd1 vssd1 vccd1 vccd1 net3420 sky130_fd_sc_hd__buf_1
XFILLER_0_39_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ net6982 net7183 _04355_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12700_ net13 _05856_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _06662_ _06784_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10892_ net6411 net7167 _04236_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12631_ net8 _05789_ _05791_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a22o_1
X_21829_ clknet_leaf_88_i_clk net3832 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15350_ _08394_ _08405_ _08411_ _08424_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__o22ai_1
X_12562_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _04994_ vssd1 vssd1 vccd1 vccd1 _05727_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _07450_ _07451_ _07418_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11513_ rbzero.spi_registers.texadd1\[14\] _04639_ _04638_ vssd1 vssd1 vccd1 vccd1
+ _04685_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15281_ _08354_ _08355_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12493_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _05262_ vssd1 vssd1 vccd1 vccd1 _05659_
+ sky130_fd_sc_hd__mux2_1
X_17020_ _10019_ _09281_ vssd1 vssd1 vccd1 vccd1 _10029_ sky130_fd_sc_hd__nand2_1
X_14232_ _07381_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__nand2_1
X_11444_ net3506 net3534 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _06880_ _07000_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__nand2_1
X_11375_ net7125 net7048 _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6190 net1732 vssd1 vssd1 vccd1 vccd1 net6714 sky130_fd_sc_hd__dlygate4sd3_1
X_13114_ _06269_ net4577 vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__and2_1
X_14094_ _07232_ _07242_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__o21a_1
X_18971_ net3998 net6249 _01749_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _01869_ _01871_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__o21ai_1
X_13045_ _06180_ net4823 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__or2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17853_ _01900_ _01901_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__and2_1
X_16804_ _09873_ _09738_ _08632_ vssd1 vssd1 vccd1 vccd1 _09874_ sky130_fd_sc_hd__a21oi_1
X_17784_ _01833_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__and2_1
X_14996_ net7566 _08051_ _08135_ net7836 _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__o221ai_4
X_19523_ _03287_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16735_ _09666_ vssd1 vssd1 vccd1 vccd1 _09805_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13947_ _07096_ _07097_ _07094_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19454_ net3180 net2964 _03241_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16666_ _08181_ _08184_ _08186_ net77 vssd1 vssd1 vccd1 vccd1 _09737_ sky130_fd_sc_hd__or4b_4
X_13878_ _07027_ _07026_ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_147_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15617_ _08688_ _08675_ _08690_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__nand3_1
X_18405_ _10010_ _02434_ _02435_ _10571_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_5_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12829_ net48 _05956_ _05958_ clknet_1_1__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _05988_
+ sky130_fd_sc_hd__a22o_2
X_16597_ _09664_ _09667_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19385_ net5487 _03198_ _03204_ _03194_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ rbzero.wall_tracer.visualWallDist\[-11\] _08298_ vssd1 vssd1 vccd1 vccd1
+ _08623_ sky130_fd_sc_hd__nand2_1
X_18336_ _02368_ _02369_ _02370_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__o21a_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18267_ _08793_ _09602_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15479_ _08130_ _08320_ _08552_ _08553_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17218_ _10217_ _10218_ vssd1 vssd1 vccd1 vccd1 _10219_ sky130_fd_sc_hd__nor2_2
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18198_ _02238_ _02243_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold703 net4589 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17149_ _09108_ _09595_ _09855_ _10150_ vssd1 vssd1 vccd1 vccd1 _10151_ sky130_fd_sc_hd__o31ai_4
Xhold714 net5573 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold725 net4921 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold736 _01472_ vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 net5241 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
X_20160_ net5582 _03691_ _03701_ _03696_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__o211a_1
Xhold758 net4849 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 net5545 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20091_ net3227 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__clkbuf_1
Xhold2104 rbzero.pov.spi_counter\[1\] vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 _04363_ vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2126 net5923 vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2137 _01386_ vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2148 _04389_ vssd1 vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 _04452_ vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _04308_ vssd1 vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 net5984 vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _01123_ vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1436 net4245 vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 net5954 vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1458 net2770 vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 net5812 vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21614_ clknet_leaf_25_i_clk net5348 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21545_ clknet_leaf_27_i_clk net1005 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21476_ clknet_leaf_102_i_clk net3073 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20427_ net3451 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__clkbuf_1
X_11160_ net5850 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4040 net936 vssd1 vssd1 vccd1 vccd1 net4564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4051 net3502 vssd1 vssd1 vccd1 vccd1 net4575 sky130_fd_sc_hd__buf_1
X_20862__281 clknet_1_0__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__inv_2
X_11091_ net6770 net6457 _04415_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4062 net3528 vssd1 vssd1 vccd1 vccd1 net4586 sky130_fd_sc_hd__dlygate4sd3_1
X_20289_ clknet_1_0__leaf__03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__buf_1
Xhold4073 net3566 vssd1 vssd1 vccd1 vccd1 net4597 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4084 _00873_ vssd1 vssd1 vccd1 vccd1 net4608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3350 _03588_ vssd1 vssd1 vccd1 vccd1 net3874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4095 net3717 vssd1 vssd1 vccd1 vccd1 net4619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3361 net7358 vssd1 vssd1 vccd1 vccd1 net3885 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22028_ clknet_leaf_96_i_clk net3759 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3372 _00596_ vssd1 vssd1 vccd1 vccd1 net3896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3383 _00624_ vssd1 vssd1 vccd1 vccd1 net3907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3394 _02729_ vssd1 vssd1 vccd1 vccd1 net3918 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2660 net4452 vssd1 vssd1 vccd1 vccd1 net3184 sky130_fd_sc_hd__buf_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2671 net7147 vssd1 vssd1 vccd1 vccd1 net3195 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _06678_ _07990_ _07994_ _08000_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__a31o_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold74 _03222_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2682 rbzero.wall_tracer.visualWallDist\[-7\] vssd1 vssd1 vccd1 vccd1 net3206
+ sky130_fd_sc_hd__clkbuf_2
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold85 net968 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2693 net4454 vssd1 vssd1 vccd1 vccd1 net3217 sky130_fd_sc_hd__buf_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _06922_ _06921_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__or2b_1
Xhold96 net4125 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1970 net5982 vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1981 net7059 vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _07930_ _07931_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1992 _01401_ vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ net3016 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__inv_2
X_16520_ _09583_ _09591_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__xnor2_1
X_13732_ net580 _06819_ _06796_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__nand3_1
XFILLER_0_202_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ net2125 net6551 _04344_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ _09405_ _09408_ _09523_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ _06813_ _06704_ _06677_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__mux2_1
X_10875_ net2715 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15402_ _08379_ _08476_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19170_ net1735 _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__or2_1
X_12614_ net83 _05778_ net4006 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__o21a_1
X_16382_ _08529_ _08498_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__nor2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ _06697_ _06698_ _06556_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__a21o_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _01967_ _01969_ _02067_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__o31ai_4
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ net3115 _08304_ _08306_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ rbzero.tex_b1\[57\] rbzero.tex_b1\[56\] _05541_ vssd1 vssd1 vccd1 vccd1 _05710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18052_ _01684_ _01711_ _10539_ _10520_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15264_ net7402 _06492_ _06500_ _06482_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__and4b_1
X_12476_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _05230_ vssd1 vssd1 vccd1 vccd1 _05642_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17003_ _10013_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__clkbuf_1
X_14215_ _06973_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11427_ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_5 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20945__356 clknet_1_0__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__inv_2
X_15195_ net65 net4007 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _07070_ _07024_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__and2b_1
X_11358_ net6477 net2295 _04562_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14077_ _07182_ _07181_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__nor2_1
X_18954_ _02934_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11289_ net1930 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17905_ _01953_ _01954_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__nor2_1
X_13028_ net6185 _06178_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__and2_1
X_18885_ _02870_ _02871_ _02844_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _01883_ _01884_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer17 _06896_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ _01816_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__nor2_1
Xrebuffer28 _06819_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_1
Xrebuffer39 net562 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14979_ _08101_ _08121_ _08069_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19506_ net5562 _03274_ _03278_ _03260_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__o211a_1
X_16718_ _09669_ _09786_ vssd1 vssd1 vccd1 vccd1 _09788_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17698_ _01748_ net4403 _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ net1862 _03225_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20690__126 clknet_1_1__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__inv_2
X_16649_ _08899_ _08599_ vssd1 vssd1 vccd1 vccd1 _09720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19368_ net1563 _03186_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18319_ _02360_ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19299_ net2256 _03147_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__or2_1
Xhold6904 net4300 vssd1 vssd1 vccd1 vccd1 net7428 sky130_fd_sc_hd__dlygate4sd3_1
X_21330_ clknet_leaf_57_i_clk net4253 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6915 _08119_ vssd1 vssd1 vccd1 vccd1 net7439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6926 rbzero.wall_tracer.stepDistY\[-2\] vssd1 vssd1 vccd1 vccd1 net7450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6948 net4141 vssd1 vssd1 vccd1 vccd1 net7472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6959 net4110 vssd1 vssd1 vccd1 vccd1 net7483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold500 net4249 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
X_21261_ clknet_leaf_71_i_clk net3720 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold511 _03522_ vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 net5392 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 net5399 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20212_ _03678_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__buf_2
X_21192_ net4791 _02528_ _02579_ _04148_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold544 net5496 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 net5478 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _01282_ vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 net4286 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 _01382_ vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
X_20143_ _03678_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold599 net5561 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20074_ net3809 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 net6653 vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 net6289 vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 _00934_ vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 _04485_ vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1244 net7667 vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 _01481_ vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 net7674 vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1277 _04509_ vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1288 net6961 vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _01419_ vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ net1762 net5821 _04192_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12330_ _05496_ _05497_ _04991_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21528_ clknet_leaf_28_i_clk net2954 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ net4288 _05381_ _05420_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21459_ clknet_leaf_25_i_clk net1469 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14000_ _07041_ _07068_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__xnor2_2
X_11212_ net6423 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12192_ _05356_ net3762 vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__and2b_1
X_11143_ net1927 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__clkbuf_4
Xoutput75 net140 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__buf_1
XFILLER_0_179_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15951_ _09017_ _09018_ _09024_ _09025_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__a31o_1
X_11074_ net2871 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3180 rbzero.pov.spi_buffer\[62\] vssd1 vssd1 vccd1 vccd1 net3704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3191 _03886_ vssd1 vssd1 vccd1 vccd1 net3715 sky130_fd_sc_hd__dlygate4sd3_1
X_14902_ _07995_ _07990_ _07994_ _08050_ net7891 vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__a311o_2
X_15882_ _08916_ _08920_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__xnor2_1
X_18670_ net4463 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__inv_2
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2490 net4531 vssd1 vssd1 vccd1 vccd1 net3014 sky130_fd_sc_hd__buf_4
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _10536_ _10531_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__or2b_1
X_14833_ _07578_ _07983_ vssd1 vssd1 vccd1 vccd1 _07984_ sky130_fd_sc_hd__xnor2_4
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17552_ _10548_ _10549_ vssd1 vssd1 vccd1 vccd1 _10551_ sky130_fd_sc_hd__and2_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _07905_ _07913_ _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__or3_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _05123_ _05142_ _05143_ _05145_ net3987 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__o32a_1
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _09453_ _09455_ _09452_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__a21boi_1
X_13715_ _06737_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__inv_2
X_10927_ net6752 net6930 _04333_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__mux2_1
X_17483_ _10479_ _10480_ vssd1 vssd1 vccd1 vccd1 _10482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14695_ _07534_ _07359_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__nor2_1
X_19222_ net5360 _03107_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__or2_1
X_16434_ _09348_ _09387_ _09386_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13646_ _06775_ _06778_ _06662_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_184_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10858_ net2459 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16365_ _09345_ _09417_ _09437_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19153_ net5322 _03066_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__or2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__05891_ _05891_ vssd1 vssd1 vccd1 vccd1 clknet_0__05891_ sky130_fd_sc_hd__clkbuf_16
X_13577_ _06606_ _06619_ _06621_ _06727_ _06722_ _06692_ vssd1 vssd1 vccd1 vccd1 _06728_
+ sky130_fd_sc_hd__mux4_2
X_10789_ _04243_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18104_ _02150_ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__nand2_1
X_15316_ net7777 _08390_ _08304_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__a21o_2
X_12528_ _04906_ _05693_ _04842_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a21o_1
X_16296_ net3539 _08328_ _08628_ _09226_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__or4_1
X_19084_ net57 _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18035_ _09582_ _01940_ _01938_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15247_ _08320_ net7589 vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__nor2_1
X_12459_ _05235_ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4809 rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 net5333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15178_ net4593 _08173_ _08260_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14129_ _06970_ _06867_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__or2_1
XFILLER_0_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19986_ net3849 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18937_ _02863_ net3135 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18868_ _02854_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_158_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17819_ _01867_ _01868_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18799_ net3699 rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _02792_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_178_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22431_ clknet_leaf_41_i_clk net4505 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6701 net1923 vssd1 vssd1 vccd1 vccd1 net7225 sky130_fd_sc_hd__dlygate4sd3_1
X_22362_ net494 net1902 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6712 _04307_ vssd1 vssd1 vccd1 vccd1 net7236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6723 net2682 vssd1 vssd1 vccd1 vccd1 net7247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6734 net2804 vssd1 vssd1 vccd1 vccd1 net7258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6745 rbzero.tex_b0\[52\] vssd1 vssd1 vccd1 vccd1 net7269 sky130_fd_sc_hd__dlygate4sd3_1
X_20928__340 clknet_1_0__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__inv_2
X_21313_ clknet_leaf_72_i_clk net4534 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6756 net2827 vssd1 vssd1 vccd1 vccd1 net7280 sky130_fd_sc_hd__dlygate4sd3_1
X_22293_ net425 net2716 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold6767 rbzero.tex_r0\[51\] vssd1 vssd1 vccd1 vccd1 net7291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6778 net2870 vssd1 vssd1 vccd1 vccd1 net7302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6789 _00840_ vssd1 vssd1 vccd1 vccd1 net7313 sky130_fd_sc_hd__dlygate4sd3_1
X_21244_ clknet_leaf_53_i_clk net3724 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold330 net5156 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 net5282 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 net5229 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 net5227 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold374 net5189 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
X_21175_ net4140 _04140_ _04141_ _09769_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__a22o_1
Xhold385 net4792 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 net5296 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20126_ _03440_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20057_ _02647_ _03614_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 net5988 vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _00915_ vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _00922_ vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 net4614 vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 net4747 vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 net5756 vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 net6597 vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__buf_4
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20974__382 clknet_1_0__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__inv_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20673__110 clknet_1_1__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__inv_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04929_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nor2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _06544_ _06650_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__and2_1
X_10712_ net2085 net7169 _04214_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _07616_ _07630_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__xor2_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _04821_ net2823 _04860_ _04759_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _06560_ _06577_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__nand2_1
X_10643_ net2405 net6906 _04181_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16150_ _08615_ _08173_ _08607_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__or3_1
X_13362_ rbzero.wall_tracer.rcp_sel\[2\] _06163_ _06512_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__a211o_1
Xrebuffer8 net531 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_1
X_15101_ _06344_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__clkbuf_4
X_12313_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _05456_ vssd1 vssd1 vccd1 vccd1 _05481_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16081_ _09150_ _09155_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ rbzero.debug_overlay.facingX\[-6\] net3796 vssd1 vssd1 vccd1 vccd1 _06444_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ _08166_ _08167_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__and2_1
X_12244_ rbzero.debug_overlay.facingX\[-8\] _05377_ _05378_ rbzero.debug_overlay.facingX\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19840_ _03476_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__clkbuf_4
X_12175_ _04815_ net4005 _05335_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11126_ net1889 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
X_19771_ net1727 _03427_ net1662 _03424_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__o211a_1
X_16983_ net4507 net4579 vssd1 vssd1 vccd1 vccd1 _09995_ sky130_fd_sc_hd__nand2_1
X_18722_ _02723_ _02724_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__xnor2_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ net6996 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
X_15934_ _09007_ _09008_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18653_ _02637_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02661_
+ sky130_fd_sc_hd__or2_1
X_15865_ _08833_ _08939_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__nand2_2
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _10257_ _09312_ _01654_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__o21ai_1
X_14816_ _07791_ _07840_ _07842_ _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18584_ _02595_ _02596_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__nand2_1
Xtop_ew_algofoogle_110 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_110/HI zeros[2] sky130_fd_sc_hd__conb_1
X_15796_ _08838_ _08870_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__xor2_2
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_121 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_121/HI zeros[13]
+ sky130_fd_sc_hd__conb_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_132 vssd1 vssd1 vccd1 vccd1 ones[8] top_ew_algofoogle_132/LO sky130_fd_sc_hd__conb_1
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17535_ _10532_ _10533_ vssd1 vssd1 vccd1 vccd1 _10534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14747_ _07774_ _07359_ _07893_ _07897_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11959_ net2069 _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17466_ _10442_ _10444_ vssd1 vssd1 vccd1 vccd1 _10465_ sky130_fd_sc_hd__or2_1
X_14678_ _07820_ _07827_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19205_ net1540 _03079_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16417_ net3722 _08313_ _09486_ _09489_ vssd1 vssd1 vccd1 vccd1 _09490_ sky130_fd_sc_hd__or4_2
X_13629_ _06772_ _06779_ _06659_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__a21oi_2
X_17397_ _10395_ _10396_ vssd1 vssd1 vccd1 vccd1 _10397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19136_ net5099 _03053_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__or2_1
X_16348_ _08326_ _09420_ vssd1 vssd1 vccd1 vccd1 _09421_ sky130_fd_sc_hd__or2_2
Xhold6008 _04304_ vssd1 vssd1 vccd1 vccd1 net6532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6019 net1526 vssd1 vssd1 vccd1 vccd1 net6543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5307 rbzero.tex_g1\[2\] vssd1 vssd1 vccd1 vccd1 net5831 sky130_fd_sc_hd__dlygate4sd3_1
X_16279_ _09351_ _09352_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__nand2_1
X_19067_ net6058 net2843 _03017_ _03011_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__o211a_1
Xhold5318 _04525_ vssd1 vssd1 vccd1 vccd1 net5842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5329 _00703_ vssd1 vssd1 vccd1 vccd1 net5853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18018_ _02065_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4606 net875 vssd1 vssd1 vccd1 vccd1 net5130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4617 _00871_ vssd1 vssd1 vccd1 vccd1 net5141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4628 _00698_ vssd1 vssd1 vccd1 vccd1 net5152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4639 net836 vssd1 vssd1 vccd1 vccd1 net5163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3905 net3174 vssd1 vssd1 vccd1 vccd1 net4429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3916 _01640_ vssd1 vssd1 vccd1 vccd1 net4440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3927 net3210 vssd1 vssd1 vccd1 vccd1 net4451 sky130_fd_sc_hd__buf_1
Xhold3938 net741 vssd1 vssd1 vccd1 vccd1 net4462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3949 net3315 vssd1 vssd1 vccd1 vccd1 net4473 sky130_fd_sc_hd__buf_1
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19969_ net1070 _03034_ _03483_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and3_1
X_21931_ clknet_leaf_8_i_clk net1484 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21862_ clknet_leaf_94_i_clk net1602 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20813_ clknet_1_1__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21793_ clknet_leaf_11_i_clk net3002 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22414_ net142 net1837 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7243 rbzero.wall_tracer.trackDistX\[9\] vssd1 vssd1 vccd1 vccd1 net7767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6520 net2298 vssd1 vssd1 vccd1 vccd1 net7044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7265 _02463_ vssd1 vssd1 vccd1 vccd1 net7789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6531 rbzero.tex_r1\[33\] vssd1 vssd1 vccd1 vccd1 net7055 sky130_fd_sc_hd__dlygate4sd3_1
X_22345_ net477 net2758 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
Xhold7276 rbzero.wall_tracer.stepDistY\[-4\] vssd1 vssd1 vccd1 vccd1 net7800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6542 net2385 vssd1 vssd1 vccd1 vccd1 net7066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7287 rbzero.wall_tracer.stepDistX\[3\] vssd1 vssd1 vccd1 vccd1 net7811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6553 net2247 vssd1 vssd1 vccd1 vccd1 net7077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7298 rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 net7822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6564 rbzero.tex_r1\[5\] vssd1 vssd1 vccd1 vccd1 net7088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5830 gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6575 net2659 vssd1 vssd1 vccd1 vccd1 net7099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22276_ net408 net2764 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
Xhold6586 rbzero.tex_g0\[8\] vssd1 vssd1 vccd1 vccd1 net7110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5841 net1107 vssd1 vssd1 vccd1 vccd1 net6365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5852 _04510_ vssd1 vssd1 vccd1 vccd1 net6376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6597 net2679 vssd1 vssd1 vccd1 vccd1 net7121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5863 net1138 vssd1 vssd1 vccd1 vccd1 net6387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5874 rbzero.tex_b0\[50\] vssd1 vssd1 vccd1 vccd1 net6398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5885 net1154 vssd1 vssd1 vccd1 vccd1 net6409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 rbzero.wall_tracer.visualWallDist\[4\] vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_1
X_21227_ clknet_leaf_50_i_clk _00396_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold171 rbzero.wall_tracer.visualWallDist\[-2\] vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_2
Xhold5896 rbzero.tex_b1\[36\] vssd1 vssd1 vccd1 vccd1 net6420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 net4365 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold193 net4986 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
X_21158_ _02488_ clknet_1_0__leaf__05942_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__and2_2
X_20705__139 clknet_1_1__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__inv_2
XFILLER_0_176_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20109_ net2937 net3825 _03664_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__and3_1
X_13980_ _06869_ _06990_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__nor2_1
X_21089_ net1100 net4701 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nand2_1
X_12931_ _06048_ _06083_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a21o_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _08317_ _08724_ _08702_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__o21ai_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ net4021 _05998_ _06007_ _05299_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a22o_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__buf_2
X_14601_ _07745_ _07749_ _07750_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nand3_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _08648_ _08651_ _08650_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__a21oi_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12793_ net4095 _05446_ net22 vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__mux2_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _10092_ _10197_ _10195_ vssd1 vssd1 vccd1 vccd1 _10321_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _07669_ _07681_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__nor2_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _04910_ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__nand2_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _10250_ _10251_ vssd1 vssd1 vccd1 vccd1 _10252_ sky130_fd_sc_hd__nand2_1
X_14463_ _07612_ _07613_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11675_ _04843_ net4063 net3028 _04714_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16202_ net2942 net7732 net4087 vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__mux2_1
X_13414_ _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__buf_2
X_17182_ _10161_ _10182_ _10183_ vssd1 vssd1 vccd1 vccd1 _10184_ sky130_fd_sc_hd__and3_1
X_10626_ net7272 net2820 _04170_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14394_ _07543_ _07544_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16133_ _08585_ _08589_ _08583_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _06445_ _06458_ _06456_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_109_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16064_ _09086_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__clkbuf_4
X_13276_ _06416_ _06426_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__and2_1
X_15015_ _08153_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
X_12227_ net4549 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__clkbuf_4
X_19823_ net3960 net3925 _03459_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ net4009 net3761 net4070 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__o21ai_1
X_11109_ net2741 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ net1613 _03392_ net5763 _03424_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__o211a_1
X_12089_ _05256_ _05257_ _05003_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__mux2_1
X_16966_ _09979_ _09980_ vssd1 vssd1 vccd1 vccd1 _09981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18705_ _02693_ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__xnor2_1
X_15917_ _08990_ _08989_ _08991_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__nand3_1
XFILLER_0_56_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19685_ net6622 _03375_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or2_1
X_16897_ net773 _09937_ _09938_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1
+ vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18636_ _02637_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _02645_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _08915_ _08922_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18567_ _05401_ rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _02581_
+ sky130_fd_sc_hd__nand2_1
X_15779_ _08844_ _08852_ _08853_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__a21o_1
X_17518_ _10515_ _10516_ vssd1 vssd1 vccd1 vccd1 _10517_ sky130_fd_sc_hd__xor2_2
XFILLER_0_8_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18498_ net1296 net3969 _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__nor3_1
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ _10446_ _10448_ vssd1 vssd1 vccd1 vccd1 _10449_ sky130_fd_sc_hd__xor2_4
XFILLER_0_172_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20810__234 clknet_1_1__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__inv_2
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20460_ net2887 net3782 _03845_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ net5876 _03037_ _03050_ _03048_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20391_ _03791_ net3586 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__and2_1
Xhold5104 rbzero.spi_registers.texadd2\[22\] vssd1 vssd1 vccd1 vccd1 net5628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5115 net1420 vssd1 vssd1 vccd1 vccd1 net5639 sky130_fd_sc_hd__dlygate4sd3_1
X_22130_ net262 net1811 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5126 _00715_ vssd1 vssd1 vccd1 vccd1 net5650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5137 _00751_ vssd1 vssd1 vccd1 vccd1 net5661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4403 rbzero.wall_tracer.trackDistX\[-2\] vssd1 vssd1 vccd1 vccd1 net4927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5148 _01072_ vssd1 vssd1 vccd1 vccd1 net5672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4414 _04092_ vssd1 vssd1 vccd1 vccd1 net4938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5159 net7833 vssd1 vssd1 vccd1 vccd1 net5683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4425 net3404 vssd1 vssd1 vccd1 vccd1 net4949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22061_ clknet_leaf_7_i_clk net3601 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4436 _01650_ vssd1 vssd1 vccd1 vccd1 net4960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3702 net1592 vssd1 vssd1 vccd1 vccd1 net4226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4447 gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 net4971 sky130_fd_sc_hd__buf_1
Xhold3713 _00912_ vssd1 vssd1 vccd1 vccd1 net4237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4458 rbzero.spi_registers.texadd1\[9\] vssd1 vssd1 vccd1 vccd1 net4982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4469 net737 vssd1 vssd1 vccd1 vccd1 net4993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3724 net1023 vssd1 vssd1 vccd1 vccd1 net4248 sky130_fd_sc_hd__dlygate4sd3_1
X_21012_ _04014_ _04015_ _04016_ _04017_ net4987 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3735 _00911_ vssd1 vssd1 vccd1 vccd1 net4259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3746 net2281 vssd1 vssd1 vccd1 vccd1 net4270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3757 _00497_ vssd1 vssd1 vccd1 vccd1 net4281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3768 _00768_ vssd1 vssd1 vccd1 vccd1 net4292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3779 net7677 vssd1 vssd1 vccd1 vccd1 net4303 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21914_ clknet_leaf_90_i_clk net1325 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21845_ clknet_leaf_82_i_clk net3245 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21776_ clknet_leaf_1_i_clk net4324 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _04162_ _04611_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__or2_2
X_20658_ clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__buf_1
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20785__211 clknet_1_0__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__inv_2
Xhold7051 _02798_ vssd1 vssd1 vccd1 vccd1 net7575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7062 _02583_ vssd1 vssd1 vccd1 vccd1 net7586 sky130_fd_sc_hd__dlygate4sd3_1
X_11391_ net6732 net2734 _04573_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20589_ net3385 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
Xhold7084 _02661_ vssd1 vssd1 vccd1 vccd1 net7608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6350 net2028 vssd1 vssd1 vccd1 vccd1 net6874 sky130_fd_sc_hd__dlygate4sd3_1
X_13130_ net3542 _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nor2_1
Xhold7095 _00506_ vssd1 vssd1 vccd1 vccd1 net7619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6361 _04463_ vssd1 vssd1 vccd1 vccd1 net6885 sky130_fd_sc_hd__dlygate4sd3_1
X_22328_ net460 net1553 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
Xhold6372 net2525 vssd1 vssd1 vccd1 vccd1 net6896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6383 _04188_ vssd1 vssd1 vccd1 vccd1 net6907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6394 net2111 vssd1 vssd1 vccd1 vccd1 net6918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5660 net677 vssd1 vssd1 vccd1 vccd1 net6184 sky130_fd_sc_hd__dlygate4sd3_1
X_13061_ net6251 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__buf_2
X_22259_ net391 net2127 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5671 net2455 vssd1 vssd1 vccd1 vccd1 net6195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5682 rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 net6206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5693 _06222_ vssd1 vssd1 vccd1 vccd1 net6217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12012_ rbzero.floor_leak\[1\] _04981_ _04987_ net1113 vssd1 vssd1 vccd1 vccd1 _05182_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4970 rbzero.pov.spi_buffer\[29\] vssd1 vssd1 vccd1 vccd1 net5494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4981 _00771_ vssd1 vssd1 vccd1 vccd1 net5505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4992 rbzero.pov.spi_buffer\[22\] vssd1 vssd1 vccd1 vccd1 net5516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ _09726_ _09750_ _09889_ vssd1 vssd1 vccd1 vccd1 _09890_ sky130_fd_sc_hd__a21o_1
X_16751_ _09672_ _09682_ _09680_ vssd1 vssd1 vccd1 vccd1 _09821_ sky130_fd_sc_hd__a21oi_1
X_13963_ _06888_ _07112_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15702_ _08749_ _08776_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__xor2_4
X_19470_ net3079 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__clkbuf_1
X_12914_ net44 net35 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__nand2_1
X_16682_ _09592_ _09620_ _09752_ vssd1 vssd1 vccd1 vccd1 _09753_ sky130_fd_sc_hd__a21oi_1
X_13894_ _06941_ _06939_ _06940_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__nand3_1
XFILLER_0_186_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18421_ _10010_ _02449_ _01862_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15633_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__clkbuf_4
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _06002_ net32 vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nor2_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18352_ _02389_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__clkbuf_1
X_15564_ _08590_ _08638_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__xnor2_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ net49 _05894_ _05903_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__a31o_2
XFILLER_0_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _10177_ _10179_ _10303_ vssd1 vssd1 vccd1 vccd1 _10304_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _07659_ _07665_ _07657_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__o21a_2
X_11727_ _04894_ _04759_ _04776_ _04895_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__o221a_1
X_15495_ _08551_ _08562_ _08569_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__a21o_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17234_ _09813_ _10109_ _10112_ vssd1 vssd1 vccd1 vccd1 _10235_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14446_ _07549_ _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__nand2_1
X_11658_ net3995 vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__clkbuf_4
X_17165_ net3502 _09304_ vssd1 vssd1 vccd1 vccd1 _10167_ sky130_fd_sc_hd__and2_1
X_14377_ _07514_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _04744_ _04749_ _04753_ _04758_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold907 net6532 vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16116_ _08707_ _09133_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__and2b_1
Xhold918 net6507 vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13328_ _06094_ _06130_ _06131_ _06132_ net7582 vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_126_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17096_ _10096_ _10097_ vssd1 vssd1 vccd1 vccd1 _10098_ sky130_fd_sc_hd__nor2_1
Xhold929 net6452 vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16047_ _09117_ _09113_ _09116_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__a21bo_1
X_13259_ net5510 _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__xnor2_1
Xhold3009 _01214_ vssd1 vssd1 vccd1 vccd1 net3533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2308 _01435_ vssd1 vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2319 _03008_ vssd1 vssd1 vccd1 vccd1 net2843 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19806_ net4322 _03426_ net1863 _03454_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__o211a_1
Xhold1607 net7011 vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 _01326_ vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
X_17998_ _02045_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__xor2_1
Xhold1629 _04200_ vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19737_ net3100 _03407_ net5719 _03413_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__o211a_1
X_16949_ _09960_ net4877 _09965_ _09966_ net2807 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19668_ net3011 _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _02627_ _02628_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19599_ net3112 _03327_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__or2_1
X_21630_ clknet_leaf_19_i_clk net4981 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21561_ clknet_leaf_19_i_clk net5300 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20512_ _03880_ net3714 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21492_ clknet_leaf_15_i_clk net2906 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20443_ net3730 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_51_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20374_ net3819 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__clkbuf_1
Xhold4200 _00607_ vssd1 vssd1 vccd1 vccd1 net4724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22113_ net245 net1090 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4211 rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 net4735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4222 net2910 vssd1 vssd1 vccd1 vccd1 net4746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4244 _02665_ vssd1 vssd1 vccd1 vccd1 net4768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3510 _05194_ vssd1 vssd1 vccd1 vccd1 net4034 sky130_fd_sc_hd__buf_2
Xhold4255 net680 vssd1 vssd1 vccd1 vccd1 net4779 sky130_fd_sc_hd__buf_4
Xhold4266 rbzero.wall_tracer.rayAddendX\[-6\] vssd1 vssd1 vccd1 vccd1 net4790 sky130_fd_sc_hd__dlygate4sd3_1
X_22044_ clknet_leaf_92_i_clk net3778 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3521 _05531_ vssd1 vssd1 vccd1 vccd1 net4045 sky130_fd_sc_hd__clkbuf_4
Xhold4277 _04153_ vssd1 vssd1 vccd1 vccd1 net4801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3532 _09927_ vssd1 vssd1 vccd1 vccd1 net4056 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_66_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold4288 _02691_ vssd1 vssd1 vccd1 vccd1 net4812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3543 _08280_ vssd1 vssd1 vccd1 vccd1 net4067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4299 _06200_ vssd1 vssd1 vccd1 vccd1 net4823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3554 _05779_ vssd1 vssd1 vccd1 vccd1 net4078 sky130_fd_sc_hd__clkbuf_4
Xhold2820 _03895_ vssd1 vssd1 vccd1 vccd1 net3344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3565 _00465_ vssd1 vssd1 vccd1 vccd1 net4089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2831 _01195_ vssd1 vssd1 vccd1 vccd1 net3355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3576 _03968_ vssd1 vssd1 vccd1 vccd1 net4100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3587 net700 vssd1 vssd1 vccd1 vccd1 net4111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2842 _03881_ vssd1 vssd1 vccd1 vccd1 net3366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3598 _00717_ vssd1 vssd1 vccd1 vccd1 net4122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2853 _00626_ vssd1 vssd1 vccd1 vccd1 net3377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2864 net949 vssd1 vssd1 vccd1 vccd1 net3388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2875 _10069_ vssd1 vssd1 vccd1 vccd1 net3399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2886 _00608_ vssd1 vssd1 vccd1 vccd1 net3410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2897 rbzero.pov.ready_buffer\[34\] vssd1 vssd1 vccd1 vccd1 net3421 sky130_fd_sc_hd__dlygate4sd3_1
X_10960_ net6435 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10891_ net2782 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ net4095 _05446_ net4 vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21828_ clknet_leaf_91_i_clk net4517 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12561_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _04994_ vssd1 vssd1 vccd1 vccd1 _05726_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21759_ clknet_leaf_23_i_clk net1688 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14300_ _07414_ _07449_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__and2_1
X_11512_ rbzero.spi_registers.texadd0\[14\] _04680_ vssd1 vssd1 vccd1 vccd1 _04684_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15280_ net3024 net4355 net4893 vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__o21ai_1
X_12492_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _05457_ vssd1 vssd1 vccd1 vccd1 _05658_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14231_ _07375_ _07380_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__or2_1
X_11443_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_19_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14162_ _07264_ _07265_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11374_ _04403_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6180 net1677 vssd1 vssd1 vccd1 vccd1 net6704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ net4342 vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__inv_2
Xhold6191 rbzero.tex_g0\[20\] vssd1 vssd1 vccd1 vccd1 net6715 sky130_fd_sc_hd__dlygate4sd3_1
X_14093_ _07221_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__or2b_1
X_18970_ _02261_ _09951_ _02947_ net3997 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a31o_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _01967_ _01969_ _01970_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a21o_1
X_13044_ _06182_ _06198_ net4822 vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a21o_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5490 net2917 vssd1 vssd1 vccd1 vccd1 net6014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ _01900_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16803_ net3528 _09486_ vssd1 vssd1 vccd1 vccd1 _09873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17783_ _10298_ _10299_ _01713_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__or3_1
X_14995_ _06734_ _08103_ net3457 vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__a21oi_1
X_19522_ _02492_ _02497_ _02498_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__and3_1
X_16734_ _09802_ _09803_ vssd1 vssd1 vccd1 vccd1 _09804_ sky130_fd_sc_hd__nor2_1
X_13946_ _06895_ _06876_ _06884_ _06953_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19453_ net1608 _03241_ net1596 _03233_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665_ _08180_ _09605_ net77 _09735_ vssd1 vssd1 vccd1 vccd1 _09736_ sky130_fd_sc_hd__a31o_1
X_13877_ _06837_ _06957_ _06955_ _06895_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__o22ai_1
X_18404_ _02432_ _02433_ _02425_ _02429_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _08688_ _08675_ _08690_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__a21o_1
X_19384_ net1574 _03199_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__or2_1
X_12828_ _05950_ net24 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__and2_1
X_16596_ _08326_ _09666_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18335_ _02374_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15547_ _08597_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__inv_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ net17 net18 net19 vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ _02296_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15478_ net4086 _06151_ _08294_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17217_ _10122_ _10215_ _10216_ vssd1 vssd1 vccd1 vccd1 _10218_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ _07578_ _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18197_ _02238_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17148_ _09854_ _09857_ vssd1 vssd1 vccd1 vccd1 _10150_ sky130_fd_sc_hd__or2b_1
Xhold704 net5211 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 net3274 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 net4923 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold737 net5577 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold748 net3290 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ _10081_ net4595 net4903 vssd1 vssd1 vccd1 vccd1 _10082_ sky130_fd_sc_hd__mux2_1
Xhold759 _01097_ vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20922__335 clknet_1_0__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__inv_2
XFILLER_0_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20090_ net3562 net3226 net4796 vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2105 _03657_ vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2116 _01415_ vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2127 net5925 vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2138 net7244 vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 _01391_ vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1404 _01335_ vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 net5986 vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1426 net6931 vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1437 net6975 vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1448 _01168_ vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1459 _04387_ vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21613_ clknet_leaf_23_i_clk net5340 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21544_ clknet_leaf_27_i_clk net877 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21475_ clknet_leaf_102_i_clk net2844 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20426_ _03814_ net3450 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__and2_1
XFILLER_0_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4030 net1092 vssd1 vssd1 vccd1 vccd1 net4554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4041 net7762 vssd1 vssd1 vccd1 vccd1 net4565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4052 net7750 vssd1 vssd1 vccd1 vccd1 net4576 sky130_fd_sc_hd__dlygate4sd3_1
X_11090_ net2403 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
Xhold4063 rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 net4587 sky130_fd_sc_hd__buf_2
X_20288_ clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__buf_1
XFILLER_0_80_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4074 net7432 vssd1 vssd1 vccd1 vccd1 net4598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4085 net768 vssd1 vssd1 vccd1 vccd1 net4609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3340 rbzero.spi_registers.buf_vinf vssd1 vssd1 vccd1 vccd1 net3864 sky130_fd_sc_hd__buf_1
X_20897__312 clknet_1_1__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__inv_2
X_22027_ clknet_leaf_96_i_clk net3294 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4096 rbzero.debug_overlay.vplaneY\[-8\] vssd1 vssd1 vccd1 vccd1 net4620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3351 _00989_ vssd1 vssd1 vccd1 vccd1 net3875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3362 _02980_ vssd1 vssd1 vccd1 vccd1 net3886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3373 net6264 vssd1 vssd1 vccd1 vccd1 net3897 sky130_fd_sc_hd__buf_2
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3384 net6024 vssd1 vssd1 vccd1 vccd1 net3908 sky130_fd_sc_hd__clkbuf_2
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2650 net4428 vssd1 vssd1 vccd1 vccd1 net3174 sky130_fd_sc_hd__buf_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3395 _02730_ vssd1 vssd1 vccd1 vccd1 net3919 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2661 net4430 vssd1 vssd1 vccd1 vccd1 net3185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold64 net5820 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2672 _00590_ vssd1 vssd1 vccd1 vccd1 net3196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2683 net6153 vssd1 vssd1 vccd1 vccd1 net3207 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 net3218 sky130_fd_sc_hd__buf_1
Xhold75 net4119 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1960 net7208 vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _06948_ _06949_ _06950_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a21bo_1
Xhold86 _03129_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net6323 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1971 _01551_ vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _07923_ _07929_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__nand2_1
X_11992_ net1600 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__inv_2
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1982 net7061 vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1993 rbzero.tex_r1\[36\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
X_10943_ net2046 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_1
X_13731_ net584 _06796_ _06819_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__a21o_2
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16450_ _09521_ net3004 vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__xor2_1
X_10874_ net7300 net6922 _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13662_ net539 _06688_ _06699_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _08475_ net4288 _06178_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__mux2_1
X_12613_ _04858_ _05700_ _05777_ _05696_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__o211a_1
X_16381_ _09452_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__and2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13593_ _06519_ _06667_ _06686_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__or3_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _01965_ _02167_ _02066_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a21o_1
X_12544_ _05062_ _05704_ _05708_ _04979_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a211o_1
X_15332_ _08096_ net7775 _08294_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18051_ _01684_ _10520_ _10168_ _10539_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__or4_1
X_12475_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _05457_ vssd1 vssd1 vccd1 vccd1 _05641_
+ sky130_fd_sc_hd__mux2_1
X_15263_ _06510_ _06507_ _06497_ net7401 vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__or4_1
XFILLER_0_152_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17002_ _10012_ net4689 _09966_ vssd1 vssd1 vccd1 vccd1 _10013_ sky130_fd_sc_hd__mux2_1
X_14214_ _07312_ _07320_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nor2_1
X_11426_ net4009 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15194_ net4096 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ _07294_ _07295_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__nor2_4
XFILLER_0_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11357_ net1895 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14076_ _07198_ _07226_ _07224_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__a21o_1
X_18953_ _02909_ _02921_ _02919_ _02903_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__o211a_1
X_11288_ net2034 net7087 _04448_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
X_17904_ _01798_ _01848_ _01846_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a21oi_1
X_20763__191 clknet_1_0__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__inv_2
X_13027_ net4912 vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__clkbuf_4
X_18884_ _02847_ _02851_ _02869_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ _01883_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__nor2_1
X_17766_ _01814_ _01815_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and2_1
Xrebuffer18 net541 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer29 net562 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_1
X_14978_ _07991_ _08120_ _08008_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19505_ net3093 _03275_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__or2_1
X_16717_ _09784_ _09786_ _08326_ vssd1 vssd1 vccd1 vccd1 _09787_ sky130_fd_sc_hd__or3b_2
X_13929_ _07073_ _07079_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17697_ net4902 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19436_ net5287 _03224_ _03232_ _03233_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__o211a_1
X_16648_ _09594_ _09598_ _09597_ vssd1 vssd1 vccd1 vccd1 _09719_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_190_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19367_ net4261 _03185_ net592 _03194_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16579_ net4384 _08296_ _09649_ _09650_ _08239_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18318_ _02359_ net4499 _02338_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19298_ net5022 _03146_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18249_ _02291_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6916 net4779 vssd1 vssd1 vccd1 vccd1 net7440 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6927 rbzero.wall_tracer.stepDistX\[-2\] vssd1 vssd1 vccd1 vccd1 net7451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21260_ clknet_leaf_71_i_clk net3629 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold501 net5337 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold512 _03524_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20211_ _03675_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__buf_2
Xhold523 net6340 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 net5458 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21191_ _02538_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__xnor2_1
Xhold545 net5498 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold556 net6346 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold567 net7640 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_1
Xhold578 net6398 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
X_20142_ _03675_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__clkbuf_4
Xhold589 net5512 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20073_ _03616_ net3808 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__or2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _01511_ vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 net6291 vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 net6641 vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1234 _01305_ vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1245 _03386_ vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 net5896 vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1267 _03250_ vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _01283_ vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 net6963 vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21527_ clknet_leaf_33_i_clk net5328 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12260_ _05421_ _05422_ _05424_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__or4_1
X_21458_ clknet_leaf_30_i_clk net5621 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ net2227 net6421 _04481_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20409_ net3388 net1168 _03801_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__mux2_1
X_12191_ _05343_ _05349_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nand2_1
X_21389_ clknet_leaf_52_i_clk _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11142_ net7071 net6756 _04448_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__mux2_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 o_reset sky130_fd_sc_hd__clkbuf_4
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__clkbuf_4
X_11073_ net7302 net6610 _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__mux2_1
X_15950_ _09019_ _09023_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__nor2_1
Xhold3170 rbzero.pov.ready_buffer\[33\] vssd1 vssd1 vccd1 vccd1 net3694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3181 net1253 vssd1 vssd1 vccd1 vccd1 net3705 sky130_fd_sc_hd__buf_1
X_14901_ net7438 _07995_ _08002_ vssd1 vssd1 vccd1 vccd1 _08050_ sky130_fd_sc_hd__nor3_1
Xhold3192 _01221_ vssd1 vssd1 vccd1 vccd1 net3716 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _08953_ _08954_ _08952_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _10519_ _10521_ _10523_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2480 _09522_ vssd1 vssd1 vccd1 vccd1 net3004 sky130_fd_sc_hd__buf_1
XFILLER_0_192_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _07979_ _07981_ _07982_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__o21ai_4
Xhold2491 net4533 vssd1 vssd1 vccd1 vccd1 net3015 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21001__3 clknet_1_0__leaf__03773_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _10548_ _10549_ vssd1 vssd1 vccd1 vccd1 _10550_ sky130_fd_sc_hd__nor2_1
Xhold1790 _04423_ vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _07912_ _07902_ _07910_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _05124_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__nand2_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _09572_ _09573_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__xnor2_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13714_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10926_ net2462 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkbuf_1
X_17482_ _10479_ _10480_ vssd1 vssd1 vccd1 vccd1 _10481_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14694_ _07534_ _07359_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__or3_1
X_20951__361 clknet_1_1__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__inv_2
X_19221_ net5883 _03106_ _03111_ _03096_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16433_ _09463_ _09505_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__xnor2_1
X_10857_ net7085 net6992 _04299_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__mux2_1
X_13645_ _06789_ _06792_ _06795_ _06716_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__o22a_4
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ net5733 _03065_ _03069_ _03061_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__o211a_1
X_16364_ _09421_ _09436_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__xor2_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ net1733 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__clkbuf_1
X_13576_ _06601_ _06602_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__xor2_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _02114_ _02149_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__or2_1
X_15315_ _08100_ _08105_ _08294_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19083_ _08274_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__buf_4
X_12527_ _05309_ _05318_ _05611_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__o21ai_1
X_16295_ net3722 _08328_ _08628_ _09368_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18034_ _02080_ _02081_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nor2_1
X_15246_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] _08300_
+ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__mux2_1
X_12458_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _05263_ vssd1 vssd1 vccd1 vccd1 _05624_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11409_ net6463 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
X_12389_ rbzero.tex_g1\[39\] rbzero.tex_g1\[38\] _05456_ vssd1 vssd1 vccd1 vccd1 _05556_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15177_ net4934 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14128_ _07003_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__or2_1
X_19985_ _03261_ net3848 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14059_ _06862_ _06990_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor2_1
X_18936_ _02863_ net3135 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18867_ _02854_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02855_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _01751_ _01754_ _01752_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__o21a_1
XFILLER_0_207_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18798_ net3700 rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _02791_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17749_ _01708_ _01699_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19419_ net4112 _03211_ net601 _03220_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20691_ clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__buf_1
XFILLER_0_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22430_ clknet_leaf_41_i_clk net4548 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22361_ net493 net2223 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold6702 rbzero.tex_g1\[39\] vssd1 vssd1 vccd1 vccd1 net7226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6713 net2696 vssd1 vssd1 vccd1 vccd1 net7237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6724 rbzero.tex_r1\[2\] vssd1 vssd1 vccd1 vccd1 net7248 sky130_fd_sc_hd__dlygate4sd3_1
X_21312_ clknet_leaf_49_i_clk net3994 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6735 rbzero.tex_g0\[61\] vssd1 vssd1 vccd1 vccd1 net7259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6746 net2799 vssd1 vssd1 vccd1 vccd1 net7270 sky130_fd_sc_hd__dlygate4sd3_1
X_22292_ net424 net2165 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold6757 rbzero.tex_r0\[56\] vssd1 vssd1 vccd1 vccd1 net7281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6768 net2848 vssd1 vssd1 vccd1 vccd1 net7292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6779 rbzero.tex_g1\[57\] vssd1 vssd1 vccd1 vccd1 net7303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21243_ clknet_leaf_70_i_clk _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold320 net5244 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 net5017 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold342 net5284 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold353 net5231 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 net7638 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
X_21174_ net4166 _04140_ _04141_ _09642_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a22o_1
Xhold375 net5191 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold386 net3069 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_1
Xhold397 net5101 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
X_20125_ net3641 _03679_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20056_ net3352 _03613_ net4588 _03602_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__o211a_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _03449_ vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 net5990 vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 net6113 vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 net6556 vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 net4616 vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 net4749 vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 net6569 vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 net6599 vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11760_ net923 net1569 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__nor2_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ net6522 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__clkbuf_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ net2677 _04776_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__xor2_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10642_ net6820 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__clkbuf_1
X_13430_ _06481_ _06568_ _06580_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__nand3_1
XFILLER_0_193_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13361_ net3206 net7582 vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ _06386_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__buf_2
X_12312_ _05279_ _05477_ _05479_ _05461_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer9 net532 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_1
X_16080_ _09131_ _09151_ _09154_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13292_ _06440_ _06441_ _06442_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__o21a_2
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12243_ rbzero.debug_overlay.facingX\[-2\] _05374_ _05372_ rbzero.debug_overlay.facingX\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a22o_1
X_15031_ _08150_ _08115_ _08047_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ net4009 _05342_ _04811_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ net6640 net6391 _04437_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
X_19770_ net6233 _03429_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__or2_1
X_16982_ _09994_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__clkbuf_1
X_18721_ _02647_ net6304 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__xor2_1
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ net6994 net2538 _04404_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
X_15933_ _08872_ _08874_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__nor2_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18652_ _02637_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02660_
+ sky130_fd_sc_hd__nand2_1
X_15864_ _08831_ _08832_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__or2_4
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _10257_ _09312_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__or3_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _07795_ _07879_ _07963_ _07965_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__a22o_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ net4587 rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _02596_
+ sky130_fd_sc_hd__nand2_1
X_15795_ _08855_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__and2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_100 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_100/HI o_rgb[12]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_111 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_111/HI zeros[3] sky130_fd_sc_hd__conb_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_122 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_122/HI zeros[14]
+ sky130_fd_sc_hd__conb_1
X_20875__292 clknet_1_1__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__inv_2
X_17534_ _10406_ _10407_ _10416_ _09108_ vssd1 vssd1 vccd1 vccd1 _10533_ sky130_fd_sc_hd__o22ai_2
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_133 vssd1 vssd1 vccd1 vccd1 ones[9] top_ew_algofoogle_133/LO sky130_fd_sc_hd__conb_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _07894_ _07896_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11958_ net3040 _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17465_ _10463_ _10453_ vssd1 vssd1 vccd1 vccd1 _10464_ sky130_fd_sc_hd__or2_1
X_10909_ net2762 net7229 _04321_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14677_ _07821_ _07822_ _07826_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__nand3_1
X_11889_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _05037_ vssd1 vssd1 vccd1 vccd1 _05059_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19204_ net2953 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16416_ _08633_ _09487_ _09488_ _08610_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__a31o_2
Xclkbuf_0__05942_ _05942_ vssd1 vssd1 vccd1 vccd1 clknet_0__05942_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _06662_ _06775_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__or3_1
X_17396_ _10392_ _10394_ vssd1 vssd1 vccd1 vccd1 _10396_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19135_ net5699 _03052_ net637 _03048_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__o211a_1
X_16347_ _09419_ vssd1 vssd1 vccd1 vccd1 _09420_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13559_ _06707_ _06708_ _06709_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__a21boi_1
Xhold6009 net1431 vssd1 vssd1 vccd1 vccd1 net6533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19066_ net3100 _03009_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5308 _04384_ vssd1 vssd1 vccd1 vccd1 net5832 sky130_fd_sc_hd__dlygate4sd3_1
X_16278_ _08588_ _09064_ _08969_ _08642_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5319 net2038 vssd1 vssd1 vccd1 vccd1 net5843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18017_ _01980_ _01981_ _02064_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and3_1
X_15229_ _08303_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__buf_4
Xhold4607 rbzero.spi_registers.buf_mapdx\[0\] vssd1 vssd1 vccd1 vccd1 net5131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4618 rbzero.spi_registers.texadd3\[15\] vssd1 vssd1 vccd1 vccd1 net5142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4629 net988 vssd1 vssd1 vccd1 vccd1 net5153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3906 net7918 vssd1 vssd1 vccd1 vccd1 net4430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3917 net724 vssd1 vssd1 vccd1 vccd1 net4441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3928 net7533 vssd1 vssd1 vccd1 vccd1 net4452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3939 rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 net4463 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19968_ _03577_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18919_ _02863_ net3090 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2_2
X_19899_ rbzero.debug_overlay.playerX\[5\] _03471_ vssd1 vssd1 vccd1 vccd1 _03525_
+ sky130_fd_sc_hd__nor2_1
X_20958__367 clknet_1_1__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__inv_2
X_21930_ clknet_leaf_8_i_clk net4835 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21861_ clknet_leaf_94_i_clk net2631 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21792_ clknet_leaf_11_i_clk net2930 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7200 net4283 vssd1 vssd1 vccd1 vccd1 net7724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22413_ net165 net1466 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7211 rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 net7735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7233 _06611_ vssd1 vssd1 vccd1 vccd1 net7757 sky130_fd_sc_hd__buf_4
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6510 net2045 vssd1 vssd1 vccd1 vccd1 net7034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7255 _08360_ vssd1 vssd1 vccd1 vccd1 net7779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6521 rbzero.tex_b1\[51\] vssd1 vssd1 vccd1 vccd1 net7045 sky130_fd_sc_hd__dlygate4sd3_1
X_22344_ net476 net2420 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
Xhold7266 _02464_ vssd1 vssd1 vccd1 vccd1 net7790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6532 net2343 vssd1 vssd1 vccd1 vccd1 net7056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7277 _02390_ vssd1 vssd1 vccd1 vccd1 net7801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6543 _04309_ vssd1 vssd1 vccd1 vccd1 net7067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7288 rbzero.wall_tracer.stepDistY\[3\] vssd1 vssd1 vccd1 vccd1 net7812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6554 rbzero.tex_r0\[52\] vssd1 vssd1 vccd1 vccd1 net7078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7299 net4333 vssd1 vssd1 vccd1 vccd1 net7823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6565 net1458 vssd1 vssd1 vccd1 vccd1 net7089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5820 _04378_ vssd1 vssd1 vccd1 vccd1 net6344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6576 rbzero.tex_g1\[40\] vssd1 vssd1 vccd1 vccd1 net7100 sky130_fd_sc_hd__dlygate4sd3_1
X_22275_ net407 net2248 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
Xhold5831 net1182 vssd1 vssd1 vccd1 vccd1 net6355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5842 rbzero.tex_g1\[38\] vssd1 vssd1 vccd1 vccd1 net6366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6587 net2521 vssd1 vssd1 vccd1 vccd1 net7111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5853 net1089 vssd1 vssd1 vccd1 vccd1 net6377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6598 rbzero.tex_b0\[48\] vssd1 vssd1 vccd1 vccd1 net7122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5864 _04477_ vssd1 vssd1 vccd1 vccd1 net6388 sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ clknet_leaf_58_i_clk _00395_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold150 net4168 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5875 net1102 vssd1 vssd1 vccd1 vccd1 net6399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5886 rbzero.tex_g1\[58\] vssd1 vssd1 vccd1 vccd1 net6410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 net4187 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5897 net1234 vssd1 vssd1 vccd1 vccd1 net6421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 net4131 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 net4974 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 net4988 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
X_21157_ _04135_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__buf_1
XFILLER_0_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20108_ net3827 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21088_ net1100 net4701 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20039_ net1298 _03613_ net4447 _03602_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__o211a_1
X_12930_ _06052_ _06084_ _06086_ net37 vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__o211a_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ net32 net33 _06015_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__and4b_1
XFILLER_0_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _07745_ _07749_ _07750_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__a21o_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11812_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__clkbuf_8
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _08573_ _08654_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _05950_ net26 vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _07669_ _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__xor2_4
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ net1257 net2158 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__or2_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17250_ _10221_ _10222_ _10249_ vssd1 vssd1 vccd1 vccd1 _10251_ sky130_fd_sc_hd__nand3_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _07597_ _07611_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11674_ net4020 rbzero.debug_overlay.playerY\[-1\] vssd1 vssd1 vccd1 vccd1 _04844_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ _09184_ _09275_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__xor2_4
XFILLER_0_37_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13413_ _06559_ _06563_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__xor2_1
X_17181_ _10179_ _10180_ _10181_ vssd1 vssd1 vccd1 vccd1 _10183_ sky130_fd_sc_hd__a21o_1
X_10625_ net2575 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14393_ _07528_ _07542_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ _08566_ _08568_ _08563_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13344_ _06433_ _06492_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_84_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16063_ _08584_ vssd1 vssd1 vccd1 vccd1 _09138_ sky130_fd_sc_hd__clkbuf_4
X_13275_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__or2_1
X_15014_ net4372 _08152_ _08138_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__mux2_1
X_12226_ _05393_ _05377_ _05379_ rbzero.debug_overlay.vplaneY\[-7\] _05394_ vssd1
+ vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19822_ net3962 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
X_12157_ net4037 _05325_ net3989 vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11108_ net7274 net6716 _04426_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12088_ rbzero.tex_r1\[15\] rbzero.tex_r1\[14\] _05014_ vssd1 vssd1 vccd1 vccd1 _05257_
+ sky130_fd_sc_hd__mux2_1
X_16965_ _09973_ _09977_ _09971_ vssd1 vssd1 vccd1 vccd1 _09980_ sky130_fd_sc_hd__a21o_1
X_19753_ _03294_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15916_ _08933_ _08948_ _08988_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__a21o_1
X_11039_ net2898 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__clkbuf_1
X_18704_ _02707_ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19684_ net6029 _03374_ net1860 _03384_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__o211a_1
X_16896_ net4254 _09937_ _09938_ net1495 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18635_ net1999 _02557_ _02636_ net4754 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _08916_ _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ net3241 rbzero.wall_tracer.rayAddendX\[-2\] _02571_ vssd1 vssd1 vccd1 vccd1
+ _02580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778_ _08845_ _08851_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__and2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17517_ _08872_ _09484_ vssd1 vssd1 vccd1 vccd1 _10516_ sky130_fd_sc_hd__nor2_1
X_14729_ _07876_ _07875_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18497_ net3885 net3904 net3913 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17448_ _10090_ _10322_ _10447_ vssd1 vssd1 vccd1 vccd1 _10448_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _08641_ vssd1 vssd1 vccd1 vccd1 _10379_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19118_ net5045 _03040_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20390_ net1598 net3585 _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5105 net1300 vssd1 vssd1 vccd1 vccd1 net5629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5116 _00711_ vssd1 vssd1 vccd1 vccd1 net5640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5127 rbzero.spi_registers.texadd2\[3\] vssd1 vssd1 vccd1 vccd1 net5651 sky130_fd_sc_hd__dlygate4sd3_1
X_19049_ net6172 _02990_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or2_1
Xhold5138 net1392 vssd1 vssd1 vccd1 vccd1 net5662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4404 net3416 vssd1 vssd1 vccd1 vccd1 net4928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5149 rbzero.spi_registers.texadd2\[5\] vssd1 vssd1 vccd1 vccd1 net5673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4415 _01603_ vssd1 vssd1 vccd1 vccd1 net4939 sky130_fd_sc_hd__dlygate4sd3_1
X_22060_ clknet_leaf_7_i_clk net3289 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4426 gpout0.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4437 rbzero.hsync vssd1 vssd1 vccd1 vccd1 net4961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3703 net7660 vssd1 vssd1 vccd1 vccd1 net4227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4448 _04801_ vssd1 vssd1 vccd1 vccd1 net4972 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21011_ _04597_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__clkbuf_4
Xhold3714 net613 vssd1 vssd1 vccd1 vccd1 net4238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4459 net779 vssd1 vssd1 vccd1 vccd1 net4983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3725 _00719_ vssd1 vssd1 vccd1 vccd1 net4249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3736 net615 vssd1 vssd1 vccd1 vccd1 net4260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3747 net7671 vssd1 vssd1 vccd1 vccd1 net4271 sky130_fd_sc_hd__buf_1
Xhold3758 net1394 vssd1 vssd1 vccd1 vccd1 net4282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3769 net596 vssd1 vssd1 vccd1 vccd1 net4293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21913_ clknet_leaf_90_i_clk net5207 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21844_ clknet_leaf_81_i_clk net1252 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21775_ clknet_leaf_2_i_clk net1633 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7030 net7377 vssd1 vssd1 vccd1 vccd1 net7554 sky130_fd_sc_hd__clkbuf_2
X_11390_ net2609 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7052 _02800_ vssd1 vssd1 vccd1 vccd1 net7576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20588_ _03924_ net3384 vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__and2_1
Xhold7074 _02878_ vssd1 vssd1 vccd1 vccd1 net7598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6340 net2341 vssd1 vssd1 vccd1 vccd1 net6864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7085 _02666_ vssd1 vssd1 vccd1 vccd1 net7609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6351 rbzero.tex_g1\[16\] vssd1 vssd1 vccd1 vccd1 net6875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7096 rbzero.spi_registers.buf_texadd0\[13\] vssd1 vssd1 vccd1 vccd1 net7620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6362 net2213 vssd1 vssd1 vccd1 vccd1 net6886 sky130_fd_sc_hd__dlygate4sd3_1
X_22327_ net459 net2309 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
Xhold6373 rbzero.tex_r1\[7\] vssd1 vssd1 vccd1 vccd1 net6897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6384 net2470 vssd1 vssd1 vccd1 vccd1 net6908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6395 rbzero.tex_b0\[3\] vssd1 vssd1 vccd1 vccd1 net6919 sky130_fd_sc_hd__dlygate4sd3_1
X_13060_ net6248 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__clkbuf_4
Xhold5650 net1691 vssd1 vssd1 vccd1 vccd1 net6174 sky130_fd_sc_hd__dlygate4sd3_1
X_22258_ net390 net1782 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
Xhold5661 net6208 vssd1 vssd1 vccd1 vccd1 net6185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5672 rbzero.spi_registers.spi_buffer\[9\] vssd1 vssd1 vccd1 vccd1 net6196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ net3026 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__inv_2
Xhold5683 net3917 vssd1 vssd1 vccd1 vccd1 net6207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21209_ net4965 net65 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__nor2_1
Xhold5694 _02958_ vssd1 vssd1 vccd1 vccd1 net6218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4960 rbzero.pov.spi_buffer\[26\] vssd1 vssd1 vccd1 vccd1 net5484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22189_ net321 net1334 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold4971 _01065_ vssd1 vssd1 vccd1 vccd1 net5495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4982 net1165 vssd1 vssd1 vccd1 vccd1 net5506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4993 net1288 vssd1 vssd1 vccd1 vccd1 net5517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20652__91 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__inv_2
X_16750_ _09809_ _09819_ vssd1 vssd1 vccd1 vccd1 _09820_ sky130_fd_sc_hd__xnor2_1
X_13962_ _06888_ net548 vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__nor2_1
X_15701_ _08768_ _08774_ _08775_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12913_ _06048_ _06069_ net36 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__a21bo_1
X_16681_ _09617_ _09619_ vssd1 vssd1 vccd1 vccd1 _09752_ sky130_fd_sc_hd__and2b_1
X_13893_ _06946_ _07043_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__or2b_4
X_18420_ _02447_ _02448_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__xnor2_1
X_15632_ _08706_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__buf_2
XFILLER_0_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ net31 vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__inv_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _02388_ net4485 _02338_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15563_ _08621_ _08637_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__xor2_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12775_ clknet_1_1__leaf__04800_ _05894_ _05905_ vssd1 vssd1 vccd1 vccd1 _05935_
+ sky130_fd_sc_hd__and3_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _10297_ _10302_ vssd1 vssd1 vccd1 vccd1 _10303_ sky130_fd_sc_hd__xnor2_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _07660_ _07663_ _07664_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__a21boi_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ net2825 _04602_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__xnor2_1
X_18282_ _02274_ _02326_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__or2_1
X_15494_ _08567_ _08568_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ _10232_ _10233_ vssd1 vssd1 vccd1 vccd1 _10234_ sky130_fd_sc_hd__xor2_1
X_14445_ _07525_ _07526_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11657_ net3279 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10608_ _04168_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__buf_4
X_17164_ _10162_ _10165_ vssd1 vssd1 vccd1 vccd1 _10166_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14376_ _07361_ _07403_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11588_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__buf_4
X_16115_ _09188_ _09189_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__nand2_1
Xhold908 _01468_ vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13327_ _06472_ _06477_ _06433_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a21oi_2
X_17095_ _09051_ _09662_ _10095_ vssd1 vssd1 vccd1 vccd1 _10097_ sky130_fd_sc_hd__a21oi_1
Xhold919 net6509 vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16046_ _09078_ _09079_ _09120_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ net5491 _06396_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__a21oi_1
X_12209_ _05376_ _05348_ _05357_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__and3b_2
XFILLER_0_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _04863_ _06222_ net4913 net2536 vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__a22o_1
Xhold2309 net4775 vssd1 vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19805_ net1862 _03428_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__or2_1
Xhold1608 _04390_ vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_17997_ _01812_ _09861_ _01923_ _01921_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__o31a_1
XFILLER_0_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1619 net6991 vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_19736_ net5718 _03408_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__or2_1
X_16948_ net4902 vssd1 vssd1 vccd1 vccd1 _09966_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667_ _03361_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__buf_2
X_16879_ net4275 _09934_ _09936_ _08074_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18618_ _05401_ net3838 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19598_ net5318 _03325_ _03334_ _03330_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18549_ _02561_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21560_ clknet_leaf_19_i_clk net1053 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20734__166 clknet_1_0__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__inv_2
XFILLER_0_30_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20511_ net3713 net1375 _03867_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21491_ clknet_leaf_15_i_clk net2926 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20442_ _03836_ net3729 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__and2_1
X_20323__57 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
XFILLER_0_7_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20373_ _08279_ net3818 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22112_ net244 net2868 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold4201 net1582 vssd1 vssd1 vccd1 vccd1 net4725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4212 net851 vssd1 vssd1 vccd1 vccd1 net4736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4223 rbzero.pov.ready_buffer\[8\] vssd1 vssd1 vccd1 vccd1 net4747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4234 _02881_ vssd1 vssd1 vccd1 vccd1 net4758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4245 _00587_ vssd1 vssd1 vccd1 vccd1 net4769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3500 _01256_ vssd1 vssd1 vccd1 vccd1 net4024 sky130_fd_sc_hd__dlygate4sd3_1
X_22043_ clknet_leaf_92_i_clk net3522 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3511 _01258_ vssd1 vssd1 vccd1 vccd1 net4035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4256 _08243_ vssd1 vssd1 vccd1 vccd1 net4780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4267 net908 vssd1 vssd1 vccd1 vccd1 net4791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3522 _08278_ vssd1 vssd1 vccd1 vccd1 net4046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3533 _00480_ vssd1 vssd1 vccd1 vccd1 net4057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4278 _04154_ vssd1 vssd1 vccd1 vccd1 net4802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4289 _00589_ vssd1 vssd1 vccd1 vccd1 net4813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3544 _00460_ vssd1 vssd1 vccd1 vccd1 net4068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2810 net6091 vssd1 vssd1 vccd1 vccd1 net3334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3555 _08282_ vssd1 vssd1 vccd1 vccd1 net4079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2821 _01225_ vssd1 vssd1 vccd1 vccd1 net3345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3566 net6181 vssd1 vssd1 vccd1 vccd1 net4090 sky130_fd_sc_hd__buf_2
Xhold3577 _03969_ vssd1 vssd1 vccd1 vccd1 net4101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2832 rbzero.wall_tracer.visualWallDist\[-6\] vssd1 vssd1 vccd1 vccd1 net3356
+ sky130_fd_sc_hd__clkbuf_2
Xhold2843 _03882_ vssd1 vssd1 vccd1 vccd1 net3367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3588 net7624 vssd1 vssd1 vccd1 vccd1 net4112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2854 rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1 vccd1 net3378 sky130_fd_sc_hd__buf_2
Xhold3599 net605 vssd1 vssd1 vccd1 vccd1 net4123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2865 _03815_ vssd1 vssd1 vccd1 vccd1 net3389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2876 _10075_ vssd1 vssd1 vccd1 vccd1 net3400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2887 net5687 vssd1 vssd1 vccd1 vccd1 net3411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2898 net705 vssd1 vssd1 vccd1 vccd1 net3422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10890_ net7167 net7177 _04236_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21827_ clknet_leaf_88_i_clk net3903 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12560_ _05004_ _05722_ _05724_ _05000_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__o211a_1
X_21758_ clknet_leaf_23_i_clk net1711 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _04648_ _04678_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ _05655_ _05656_ _05069_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21689_ clknet_leaf_25_i_clk net5320 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14230_ _07375_ _07380_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__nand2_1
X_11442_ _04617_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_6
XFILLER_0_145_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__06044_ clknet_0__06044_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__06044_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11373_ net6950 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
X_14161_ _07311_ _06990_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__or2_1
Xhold6170 net1709 vssd1 vssd1 vccd1 vccd1 net6694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6181 _04270_ vssd1 vssd1 vccd1 vccd1 net6705 sky130_fd_sc_hd__dlygate4sd3_1
X_13112_ net3622 net4899 vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__nor2_1
Xhold6192 net1917 vssd1 vssd1 vccd1 vccd1 net6716 sky130_fd_sc_hd__dlygate4sd3_1
X_14092_ _07218_ _07220_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5480 rbzero.map_overlay.i_othery\[1\] vssd1 vssd1 vccd1 vccd1 net6004 sky130_fd_sc_hd__dlygate4sd3_1
X_17920_ _01967_ _01969_ _06205_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__o21ai_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5491 _00657_ vssd1 vssd1 vccd1 vccd1 net6015 sky130_fd_sc_hd__dlygate4sd3_1
X_13043_ net4821 net3034 _06179_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17851_ _01777_ _01788_ _01786_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a21oi_1
Xhold4790 net964 vssd1 vssd1 vccd1 vccd1 net5314 sky130_fd_sc_hd__dlygate4sd3_1
X_16802_ net4828 _08664_ _09870_ vssd1 vssd1 vccd1 vccd1 _09872_ sky130_fd_sc_hd__or3b_1
XFILLER_0_156_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17782_ _10301_ _01713_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14994_ _08092_ _08133_ _08134_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_89_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16733_ _09800_ _09801_ vssd1 vssd1 vccd1 vccd1 _09803_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19521_ net5375 _03274_ _03286_ _03280_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13945_ _07094_ _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19452_ _02492_ _02498_ _03238_ net6245 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16664_ _08186_ vssd1 vssd1 vccd1 vccd1 _09735_ sky130_fd_sc_hd__inv_2
X_13876_ _06885_ _06929_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _08689_ _08531_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__xor2_1
X_18403_ _02425_ _02429_ _02432_ _02433_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_9_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19383_ net5523 _03198_ _03203_ _03194_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__o211a_1
X_12827_ net57 _05958_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a21o_1
X_16595_ net7441 vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _02373_ net4511 _02338_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
X_15546_ _08603_ _08620_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__xor2_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12758_ net4060 _05904_ _05905_ _05816_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18265_ _02300_ _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__xnor2_1
X_11709_ _04872_ _04873_ _04874_ _04875_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a221o_1
X_15477_ _08300_ _06489_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12689_ net14 _05847_ _05848_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17216_ _10122_ _10215_ _10216_ vssd1 vssd1 vccd1 vccd1 _10217_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14428_ _07573_ _07577_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__or2_1
X_18196_ _02241_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17147_ _10127_ _10148_ vssd1 vssd1 vccd1 vccd1 _10149_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14359_ _07473_ _07475_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__nand2_1
Xhold705 net5213 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 net5450 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 net3322 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 net5579 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17078_ _10010_ net3401 _10079_ _10080_ vssd1 vssd1 vccd1 vccd1 _10081_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold749 net5603 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16029_ _09086_ _08517_ _09085_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2106 _03662_ vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2117 net7148 vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2128 _01111_ vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2139 _04405_ vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1405 net2033 vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _01365_ vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 _04400_ vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _04546_ vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1449 net6701 vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19719_ net6202 _03395_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21612_ clknet_leaf_25_i_clk net5437 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21543_ clknet_leaf_26_i_clk net5130 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21474_ clknet_leaf_0_i_clk net3101 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20425_ net3449 net1389 _03823_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20356_ clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__buf_1
XFILLER_0_114_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4020 net1457 vssd1 vssd1 vccd1 vccd1 net4544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4031 net7549 vssd1 vssd1 vccd1 vccd1 net4555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4042 net3471 vssd1 vssd1 vccd1 vccd1 net4566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20287_ net4861 _03675_ _03772_ _08276_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4053 net3518 vssd1 vssd1 vccd1 vccd1 net4577 sky130_fd_sc_hd__clkbuf_2
Xhold4064 _03634_ vssd1 vssd1 vccd1 vccd1 net4588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3330 _02960_ vssd1 vssd1 vccd1 vccd1 net3854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4075 net3555 vssd1 vssd1 vccd1 vccd1 net4599 sky130_fd_sc_hd__buf_1
X_22026_ clknet_leaf_97_i_clk net3355 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4086 net7748 vssd1 vssd1 vccd1 vccd1 net4610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3341 _03299_ vssd1 vssd1 vccd1 vccd1 net3865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3352 rbzero.debug_overlay.facingY\[10\] vssd1 vssd1 vccd1 vccd1 net3876 sky130_fd_sc_hd__buf_2
Xhold4097 _02754_ vssd1 vssd1 vccd1 vccd1 net4621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3363 _02981_ vssd1 vssd1 vccd1 vccd1 net3887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3374 _03030_ vssd1 vssd1 vccd1 vccd1 net3898 sky130_fd_sc_hd__buf_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2640 net6068 vssd1 vssd1 vccd1 vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3385 _05331_ vssd1 vssd1 vccd1 vccd1 net3909 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2651 net3346 vssd1 vssd1 vccd1 vccd1 net3175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3396 _00593_ vssd1 vssd1 vccd1 vccd1 net3920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2662 net3577 vssd1 vssd1 vccd1 vccd1 net3186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold65 net5822 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2673 rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 net3197 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold76 net1988 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2684 _00417_ vssd1 vssd1 vccd1 vccd1 net3208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1950 _01580_ vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2695 net7319 vssd1 vssd1 vccd1 vccd1 net3219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net4150 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1961 _04213_ vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1972 rbzero.tex_g1\[56\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _03028_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_1
X_11991_ net2993 vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__inv_2
Xhold1983 _01515_ vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1994 net2152 vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_13730_ _06830_ _06832_ _06835_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__nand3_4
X_10942_ net6551 net7034 _04344_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ _06743_ _06808_ _06811_ _06659_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10873_ _04243_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15400_ _08473_ _08474_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__and2_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12612_ net4077 _05701_ _05776_ _05189_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a211o_1
X_20717__150 clknet_1_1__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__inv_2
X_16380_ _08564_ _08873_ _08565_ _08471_ vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__o22ai_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _06742_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _06156_ _06507_ net4086 vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12543_ _04984_ _05705_ _05707_ _05035_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__o211a_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18050_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15262_ rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\] _06427_
+ _06418_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__or4_1
X_12474_ _05069_ _05637_ _05639_ _05244_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17001_ _06206_ _10009_ _10011_ vssd1 vssd1 vccd1 vccd1 _10012_ sky130_fd_sc_hd__o21ai_1
X_14213_ _07324_ _07335_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__nor2_1
X_11425_ net3993 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ _08276_ net4095 vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__and2_1
X_20302__38 clknet_1_1__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XFILLER_0_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14144_ _07291_ _07293_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__and2_1
X_11356_ net6822 net6477 _04562_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14075_ _07224_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__and2b_1
X_18952_ _02932_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__nand2_1
X_11287_ net2035 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
X_17903_ _01909_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__xnor2_1
X_13026_ _06181_ _06179_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__xnor2_1
X_18883_ _02847_ _02851_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17834_ _01768_ _01769_ _01767_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17765_ _01814_ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__nor2_1
X_14977_ _07996_ _07975_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__xnor2_1
Xrebuffer19 net542 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19504_ net5367 _03274_ _03277_ _03260_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_50_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16716_ _09660_ _09689_ _09785_ vssd1 vssd1 vccd1 vccd1 _09786_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13928_ _07074_ _07075_ net571 net574 vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__a22o_1
X_17696_ _06206_ net7376 _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_187_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16647_ _09586_ _09587_ _09717_ vssd1 vssd1 vccd1 vccd1 _09718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19435_ _03141_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13859_ _07008_ _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ net7407 _09648_ _08633_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__a21o_1
X_19366_ _03141_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18317_ _02357_ _02358_ _10021_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15529_ _08068_ _08149_ _08151_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__a21oi_1
X_19297_ _03141_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18248_ _02292_ _02293_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__xor2_1
Xhold6906 _08170_ vssd1 vssd1 vccd1 vccd1 net7430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6917 _09665_ vssd1 vssd1 vccd1 vccd1 net7441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ _02219_ _02224_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 net5339 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20210_ net3530 _03717_ _03729_ _03722_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__o211a_1
Xhold513 _00968_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold524 _04158_ vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
X_21190_ _02530_ net4477 vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__and2b_1
Xhold535 net5460 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 net5466 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _04013_ vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
X_20141_ net5209 _03676_ _03690_ _03683_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold568 net4553 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 net6400 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20072_ net3807 net3189 _03580_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__mux2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 net6224 vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 net6292 vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1224 net6643 vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1235 net6743 vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1246 net6105 vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 net5898 vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1268 net6226 vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold1279 net6797 vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21526_ clknet_leaf_34_i_clk net2976 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21457_ clknet_leaf_30_i_clk net3377 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11210_ net2588 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20408_ _08275_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__buf_2
X_12190_ _05326_ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__nand2_2
X_21388_ clknet_leaf_53_i_clk _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11141_ net2617 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__clkbuf_4
X_11072_ _04403_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3160 net1224 vssd1 vssd1 vccd1 vccd1 net3684 sky130_fd_sc_hd__dlygate4sd3_1
X_14900_ net4311 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__clkbuf_1
Xhold3171 net857 vssd1 vssd1 vccd1 vccd1 net3695 sky130_fd_sc_hd__dlygate4sd3_1
X_22009_ clknet_leaf_100_i_clk net3820 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _08952_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__and3_1
Xhold3182 _03920_ vssd1 vssd1 vccd1 vccd1 net3706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3193 net4618 vssd1 vssd1 vccd1 vccd1 net3717 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2470 _00487_ vssd1 vssd1 vccd1 vccd1 net2994 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2481 net4309 vssd1 vssd1 vccd1 vccd1 net3005 sky130_fd_sc_hd__dlygate4sd3_1
X_14831_ _07502_ _07566_ _07576_ _07981_ _07979_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_203_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2492 net4316 vssd1 vssd1 vccd1 vccd1 net3016 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_192_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1780 net6771 vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
X_17550_ _10414_ _10426_ _10425_ vssd1 vssd1 vccd1 vccd1 _10549_ sky130_fd_sc_hd__a21boi_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1791 _01361_ vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
X_14762_ _07902_ _07910_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__a21oi_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _05122_ _05123_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__or2_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _08564_ _08497_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__buf_4
X_10925_ net6930 net7127 _04333_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
X_17481_ _09091_ _09666_ _10345_ _10346_ vssd1 vssd1 vccd1 vccd1 _10480_ sky130_fd_sc_hd__o31a_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14693_ _07532_ _07523_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16432_ _09502_ _09504_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__xor2_2
XFILLER_0_168_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19220_ net5302 _03107_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__or2_1
X_13644_ _06725_ _06794_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10856_ net6700 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ net5079 _03066_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__or2_1
X_16363_ _09433_ _09435_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13575_ _06721_ _06723_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__o21ai_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ net6714 net6465 _04255_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18102_ _02114_ _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__nand2_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _08300_ _06500_ _08320_ _08388_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _05690_ net4082 net4077 vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__mux2_2
X_19082_ net6033 net2842 net2949 _03022_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__o211a_1
X_16294_ _08296_ _09366_ _09367_ _08609_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18033_ _02016_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15245_ _08319_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ _05621_ _05622_ _05003_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ net6461 net2793 _04584_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__mux2_1
X_15176_ net3273 _08168_ net4933 vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__mux2_1
X_12388_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _05476_ vssd1 vssd1 vccd1 vccd1 _05555_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _06997_ _07005_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__and2b_1
X_11339_ net7030 net6888 _04551_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__mux2_1
X_19984_ rbzero.debug_overlay.facingX\[-4\] net3775 _03581_ vssd1 vssd1 vccd1 vccd1
+ _03589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14058_ _07201_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__nor2_1
X_18935_ _02529_ net4818 _02909_ net3091 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _06164_ _06099_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18866_ net4708 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17817_ _01865_ _01866_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__or2b_1
XFILLER_0_94_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18797_ net3699 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__clkbuf_1
X_17748_ _01688_ _01690_ _01692_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17679_ _01729_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19418_ net1989 _03212_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19349_ net1217 _03173_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7415 net656 vssd1 vssd1 vccd1 vccd1 net7939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22360_ net492 net2081 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6703 net2674 vssd1 vssd1 vccd1 vccd1 net7227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6714 rbzero.tex_b1\[53\] vssd1 vssd1 vccd1 vccd1 net7238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6725 net2723 vssd1 vssd1 vccd1 vccd1 net7249 sky130_fd_sc_hd__dlygate4sd3_1
X_21311_ clknet_leaf_49_i_clk net4057 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6736 net2671 vssd1 vssd1 vccd1 vccd1 net7260 sky130_fd_sc_hd__dlygate4sd3_1
X_22291_ net423 net2564 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6747 rbzero.tex_r1\[55\] vssd1 vssd1 vccd1 vccd1 net7271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6758 net2756 vssd1 vssd1 vccd1 vccd1 net7282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6769 rbzero.tex_b0\[55\] vssd1 vssd1 vccd1 vccd1 net7293 sky130_fd_sc_hd__dlygate4sd3_1
X_21242_ clknet_leaf_65_i_clk _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold310 net5096 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 net3336 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 net5019 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 net5123 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
X_21173_ net4164 _04140_ _04141_ _09521_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold354 net5082 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 net4420 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 net5258 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _03346_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
X_20124_ net3641 _03676_ net5572 _03636_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__o211a_1
Xhold398 net5103 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
X_20986__13 clknet_1_1__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
XFILLER_0_99_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20055_ net4587 _03614_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__or2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 net6301 vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1021 _00940_ vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _01447_ vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _03450_ vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 _03979_ vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 net5735 vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 net4264 vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 net6571 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 _01118_ vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ clknet_1_0__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__buf_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ net2728 net6520 _04214_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11690_ net2705 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ net2469 net6818 _04181_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ _06414_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12311_ _05229_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21509_ clknet_leaf_44_i_clk net1069 vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13291_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20659__97 clknet_1_0__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__inv_2
X_15030_ _08092_ _08163_ _08165_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__o21ai_2
X_20829__251 clknet_1_0__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__inv_2
X_12242_ _05195_ _05400_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__or3_2
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _04612_ _04615_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ net1986 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
X_16981_ _09993_ net4568 _09966_ vssd1 vssd1 vccd1 vccd1 _09994_ sky130_fd_sc_hd__mux2_1
X_18720_ _02718_ _02719_ _02717_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__o21a_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ net6576 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
X_15932_ _09004_ _09005_ _09006_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__a21oi_1
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15863_ _08890_ _08937_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__nor2_1
X_18651_ net6095 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17602_ _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__xnor2_1
X_14814_ _07795_ _07964_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _08855_ _08856_ _08867_ _08868_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__nand4_1
XFILLER_0_157_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18582_ net4587 rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _02595_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_101 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_101/HI o_rgb[13]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_112 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_112/HI zeros[4] sky130_fd_sc_hd__conb_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_123 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_123/HI zeros[15]
+ sky130_fd_sc_hd__conb_1
X_17533_ _09103_ _10406_ _10407_ _10415_ vssd1 vssd1 vccd1 vccd1 _10532_ sky130_fd_sc_hd__or4_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _07893_ _07895_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_134 vssd1 vssd1 vccd1 vccd1 ones[10] top_ew_algofoogle_134/LO sky130_fd_sc_hd__conb_1
XFILLER_0_197_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net2955 _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17464_ _10449_ vssd1 vssd1 vccd1 vccd1 _10463_ sky130_fd_sc_hd__inv_2
X_10908_ net5895 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__clkbuf_1
X_14676_ _07821_ _07822_ _07826_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11888_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _05037_ vssd1 vssd1 vccd1 vccd1 _05058_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19203_ _03088_ net2952 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16415_ _08180_ net77 vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__nand2_1
X_13627_ _06776_ _06777_ _06677_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17395_ _10392_ _10394_ vssd1 vssd1 vccd1 vccd1 _10395_ sky130_fd_sc_hd__nor2_1
X_10839_ net6676 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__clkbuf_1
X_16346_ _09305_ _09418_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__or2_1
X_19134_ net930 _03053_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or2_1
X_13558_ _06584_ _06678_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _05263_ vssd1 vssd1 vccd1 vccd1 _05675_
+ sky130_fd_sc_hd__mux2_1
X_19065_ net3100 net2843 _03016_ _03011_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__o211a_1
X_16277_ _08449_ _09064_ _08574_ _08588_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13489_ _06638_ _06600_ _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5309 net2443 vssd1 vssd1 vccd1 vccd1 net5833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18016_ _01980_ _01981_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a21oi_1
X_15228_ net3506 net3534 _06207_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__and3_2
XFILLER_0_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4608 net801 vssd1 vssd1 vccd1 vccd1 net5132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4619 net902 vssd1 vssd1 vccd1 vccd1 net5143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15159_ net4717 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
Xhold3907 net3185 vssd1 vssd1 vccd1 vccd1 net4431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3929 net3184 vssd1 vssd1 vccd1 vccd1 net4453 sky130_fd_sc_hd__buf_1
X_19967_ _03035_ _03473_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__nand2_4
XFILLER_0_120_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18918_ _02529_ net7581 net4663 net3481 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a31o_1
X_19898_ _03502_ net1036 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18849_ net1580 _02830_ _02836_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_179_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21860_ clknet_leaf_94_i_clk net3228 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21791_ clknet_leaf_11_i_clk net4302 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22412_ net164 net2429 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
Xhold7201 rbzero.texu_hot\[5\] vssd1 vssd1 vccd1 vccd1 net7725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7212 net4341 vssd1 vssd1 vccd1 vccd1 net7736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7223 rbzero.wall_tracer.trackDistX\[4\] vssd1 vssd1 vccd1 vccd1 net7747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6500 net2548 vssd1 vssd1 vccd1 vccd1 net7024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7245 _08600_ vssd1 vssd1 vccd1 vccd1 net7769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6511 rbzero.tex_r0\[22\] vssd1 vssd1 vccd1 vccd1 net7035 sky130_fd_sc_hd__dlygate4sd3_1
X_22343_ net475 net1150 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
Xhold7256 rbzero.wall_tracer.stepDistY\[-7\] vssd1 vssd1 vccd1 vccd1 net7780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6522 net2249 vssd1 vssd1 vccd1 vccd1 net7046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7267 rbzero.wall_tracer.stepDistY\[-11\] vssd1 vssd1 vccd1 vccd1 net7791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6533 rbzero.tex_r0\[16\] vssd1 vssd1 vccd1 vccd1 net7057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6544 rbzero.tex_r0\[17\] vssd1 vssd1 vccd1 vccd1 net7068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7289 net4377 vssd1 vssd1 vccd1 vccd1 net7813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6555 net1976 vssd1 vssd1 vccd1 vccd1 net7079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5810 _04587_ vssd1 vssd1 vccd1 vccd1 net6334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5821 net829 vssd1 vssd1 vccd1 vccd1 net6345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22274_ net406 net2255 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
Xhold6566 _04234_ vssd1 vssd1 vccd1 vccd1 net7090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6577 net2310 vssd1 vssd1 vccd1 vccd1 net7101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5832 gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5843 net1061 vssd1 vssd1 vccd1 vccd1 net6367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6588 rbzero.tex_g0\[40\] vssd1 vssd1 vccd1 vccd1 net7112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6599 net2502 vssd1 vssd1 vccd1 vccd1 net7123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5854 rbzero.tex_g0\[22\] vssd1 vssd1 vccd1 vccd1 net6378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5865 net1139 vssd1 vssd1 vccd1 vccd1 net6389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 net4964 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ clknet_leaf_50_i_clk _00394_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5876 _04543_ vssd1 vssd1 vccd1 vccd1 net6400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 rbzero.pov.ready_buffer\[70\] vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 rbzero.wall_tracer.visualWallDist\[1\] vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_1
Xhold5887 net1120 vssd1 vssd1 vccd1 vccd1 net6411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net3087 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5898 _04488_ vssd1 vssd1 vccd1 vccd1 net6422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 net4976 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 net7632 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ _02488_ clknet_1_0__leaf__05891_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__and2_2
X_20107_ _03667_ net3562 net3826 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__and3b_1
X_21087_ _04018_ _04079_ _04080_ _04017_ net4542 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a32o_1
XFILLER_0_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20038_ net4446 _03614_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ net4043 _06012_ _06016_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a211o_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11811_ _04953_ _04971_ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__or3_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ net25 vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__inv_2
X_21989_ net214 net2348 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _07670_ _07679_ _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__a21oi_4
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _04910_ _04911_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__xnor2_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20329__63 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _07597_ _07611_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nor2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ net3964 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__inv_2
XFILLER_0_194_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16200_ _09273_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__and2_4
XFILLER_0_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13412_ _06560_ _06561_ _06562_ _06541_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a31o_1
X_17180_ _10179_ _10180_ _10181_ vssd1 vssd1 vccd1 vccd1 _10182_ sky130_fd_sc_hd__nand3_1
X_10624_ net2820 net5828 _04170_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14392_ _07528_ _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16131_ _09185_ _09205_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13343_ net7582 _06152_ _06493_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16062_ _09129_ _09136_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13274_ rbzero.wall_tracer.visualWallDist\[-9\] _06166_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15013_ _08068_ _08149_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__a21o_4
X_12225_ rbzero.debug_overlay.vplaneY\[-9\] _05382_ _05378_ rbzero.debug_overlay.vplaneY\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a22o_1
X_19821_ _02967_ net3961 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__and2_1
X_12156_ net4037 _04615_ _05324_ _04614_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11107_ net6381 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19752_ net5762 _03394_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__or2_1
X_12087_ rbzero.tex_r1\[13\] rbzero.tex_r1\[12\] _05014_ vssd1 vssd1 vccd1 vccd1 _05256_
+ sky130_fd_sc_hd__mux2_1
X_16964_ net5746 _09968_ vssd1 vssd1 vccd1 vccd1 _09979_ sky130_fd_sc_hd__xnor2_1
X_18703_ _02647_ net4587 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__nand2_1
X_15915_ _08875_ _08983_ _08984_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__and3_1
X_11038_ net7296 net6802 _04392_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19683_ _03294_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__clkbuf_4
X_16895_ net4280 _09937_ _09938_ net1393 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _09943_ net4753 _02643_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__or3_1
XFILLER_0_189_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _08849_ _08665_ _08917_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18565_ _09935_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__clkbuf_4
X_15777_ _08845_ _08851_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__xor2_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _06140_ _06141_ _06136_ _06142_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__o221a_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ _08873_ _09595_ vssd1 vssd1 vccd1 vccd1 _10515_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14728_ _07843_ _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__and2_1
X_18496_ net3885 _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17447_ _10320_ _10321_ vssd1 vssd1 vccd1 vccd1 _10447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ _06859_ _07805_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17378_ _08701_ _08540_ _08643_ _08317_ vssd1 vssd1 vccd1 vccd1 _10378_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19117_ net5959 _03037_ _03049_ _03048_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__o211a_1
X_16329_ _09300_ _09402_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5106 _00776_ vssd1 vssd1 vccd1 vccd1 net5630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5117 rbzero.spi_registers.texadd2\[2\] vssd1 vssd1 vccd1 vccd1 net5641 sky130_fd_sc_hd__dlygate4sd3_1
X_19048_ net6172 _02988_ _03006_ _02993_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5128 net1330 vssd1 vssd1 vccd1 vccd1 net5652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5139 rbzero.pov.spi_buffer\[13\] vssd1 vssd1 vccd1 vccd1 net5663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4405 rbzero.trace_state\[1\] vssd1 vssd1 vccd1 vccd1 net4929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4416 net1887 vssd1 vssd1 vccd1 vccd1 net4940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4427 net658 vssd1 vssd1 vccd1 vccd1 net4951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4438 net650 vssd1 vssd1 vccd1 vccd1 net4962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4449 rbzero.wall_tracer.trackDistX\[-3\] vssd1 vssd1 vccd1 vccd1 net4973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3704 _00766_ vssd1 vssd1 vccd1 vccd1 net4228 sky130_fd_sc_hd__dlygate4sd3_1
X_21010_ net773 net4987 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nand2_1
Xhold3715 net7679 vssd1 vssd1 vccd1 vccd1 net4239 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3726 net1024 vssd1 vssd1 vccd1 vccd1 net4250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3737 net7668 vssd1 vssd1 vccd1 vccd1 net4261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3748 _00495_ vssd1 vssd1 vccd1 vccd1 net4272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3759 net7723 vssd1 vssd1 vccd1 vccd1 net4283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21912_ clknet_leaf_90_i_clk net1271 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21843_ clknet_leaf_81_i_clk net3178 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21774_ clknet_leaf_102_i_clk net1849 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7020 net4490 vssd1 vssd1 vccd1 vccd1 net7544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7031 _00520_ vssd1 vssd1 vccd1 vccd1 net7555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20711__145 clknet_1_0__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__inv_2
Xhold7042 _06660_ vssd1 vssd1 vccd1 vccd1 net7566 sky130_fd_sc_hd__clkbuf_4
Xhold7053 _00603_ vssd1 vssd1 vccd1 vccd1 net7577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20587_ net675 net3383 net3250 vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__mux2_1
Xhold6330 net2076 vssd1 vssd1 vccd1 vccd1 net6854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7075 _02883_ vssd1 vssd1 vccd1 vccd1 net7599 sky130_fd_sc_hd__dlygate4sd3_1
X_22326_ net458 net1820 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
Xhold6341 rbzero.tex_r0\[20\] vssd1 vssd1 vccd1 vccd1 net6865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6352 net2134 vssd1 vssd1 vccd1 vccd1 net6876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7097 rbzero.pov.ready_buffer\[36\] vssd1 vssd1 vccd1 vccd1 net7621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6363 rbzero.tex_b0\[38\] vssd1 vssd1 vccd1 vccd1 net6887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6374 net2079 vssd1 vssd1 vccd1 vccd1 net6898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5640 net3050 vssd1 vssd1 vccd1 vccd1 net6164 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6385 rbzero.tex_r1\[51\] vssd1 vssd1 vccd1 vccd1 net6909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22257_ net389 net2003 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold6396 net2370 vssd1 vssd1 vccd1 vccd1 net6920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5651 rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 net6175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5662 _06184_ vssd1 vssd1 vccd1 vccd1 net6186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5673 net3095 vssd1 vssd1 vccd1 vccd1 net6197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ _05175_ _05176_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__o21ai_1
Xhold5684 rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 net6208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4950 rbzero.pov.spi_buffer\[8\] vssd1 vssd1 vccd1 vccd1 net5474 sky130_fd_sc_hd__dlygate4sd3_1
X_21208_ _03502_ net1183 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__nor2_1
Xhold5695 gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 net6219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4961 _01062_ vssd1 vssd1 vccd1 vccd1 net5485 sky130_fd_sc_hd__dlygate4sd3_1
X_22188_ net320 net2529 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4972 rbzero.mapdxw\[0\] vssd1 vssd1 vccd1 vccd1 net5496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4983 rbzero.pov.spi_buffer\[4\] vssd1 vssd1 vccd1 vccd1 net5507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4994 _01058_ vssd1 vssd1 vccd1 vccd1 net5518 sky130_fd_sc_hd__dlygate4sd3_1
X_21139_ _04119_ _04121_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__a21oi_1
X_13961_ _07076_ _07078_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__xnor2_2
X_15700_ _08751_ _08767_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__nor2_1
X_12912_ _05201_ _06065_ _06066_ net73 _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a221o_1
X_16680_ _09726_ _09750_ vssd1 vssd1 vccd1 vccd1 _09751_ sky130_fd_sc_hd__xnor2_1
X_13892_ _06943_ _06944_ net585 _06891_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20792__217 clknet_1_0__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__inv_2
XFILLER_0_159_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15631_ _08313_ _08705_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__or2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ net4045 net4066 net4083 net4078 net28 net31 vssd1 vssd1 vccd1 vccd1 _06001_
+ sky130_fd_sc_hd__mux4_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _08624_ _08636_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__nand2_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _10010_ _02387_ _10055_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__o21ai_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ net19 net18 vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__and2b_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _10298_ _10299_ _10301_ vssd1 vssd1 vccd1 vccd1 _10302_ sky130_fd_sc_hd__o21a_2
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _07471_ _07359_ _07661_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ net2774 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__inv_2
X_15493_ _08529_ _08444_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18281_ _02274_ _02326_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__nand2_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17232_ _09133_ _09784_ vssd1 vssd1 vccd1 vccd1 _10233_ sky130_fd_sc_hd__nor2_1
X_14444_ _07592_ _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11656_ net3921 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17163_ _10163_ _10164_ vssd1 vssd1 vccd1 vccd1 _10165_ sky130_fd_sc_hd__xnor2_1
X_10607_ _04160_ _04166_ net89 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14375_ _07355_ _07360_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ _04604_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ _08724_ _08331_ _08698_ _09051_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20686__122 clknet_1_0__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__inv_2
XFILLER_0_122_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ _06473_ _06435_ _06474_ _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a311o_1
X_17094_ _09051_ _09662_ _10095_ vssd1 vssd1 vccd1 vccd1 _10096_ sky130_fd_sc_hd__and3_1
Xhold909 net5232 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16045_ _09039_ _09076_ _09119_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ net5491 _06396_ _06407_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12208_ _05362_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__nor2_2
X_13188_ _06270_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__or2_2
XFILLER_0_209_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19804_ net6104 _03442_ net1632 _03454_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__o211a_1
X_12139_ net4972 _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17996_ _02043_ _02044_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__xor2_1
Xhold1609 _01390_ vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19735_ net3070 _03407_ net1564 _03413_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__o211a_1
X_16947_ _06206_ net4902 vssd1 vssd1 vccd1 vccd1 _09965_ sky130_fd_sc_hd__nor2_2
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19666_ _03359_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__clkbuf_4
X_16878_ net4532 _09934_ _09936_ net4088 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18617_ _05401_ net3838 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__or2_1
X_15829_ _08902_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__or2b_1
X_19597_ net1727 _03327_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__or2_1
X_18548_ _02562_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18479_ net3151 net3074 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__and2b_2
X_20308__44 clknet_1_0__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20510_ net3575 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21490_ clknet_leaf_15_i_clk net2840 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20441_ net3728 net1292 _03823_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03999_ clknet_0__03999_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03999_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20372_ net3674 net3817 _03782_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22111_ net243 net2586 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4202 net7844 vssd1 vssd1 vccd1 vccd1 net4726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4213 _01597_ vssd1 vssd1 vccd1 vccd1 net4737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4224 net1598 vssd1 vssd1 vccd1 vccd1 net4748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4235 _02882_ vssd1 vssd1 vccd1 vccd1 net4759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3501 rbzero.trace_state\[0\] vssd1 vssd1 vccd1 vccd1 net4025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4246 net3553 vssd1 vssd1 vccd1 vccd1 net4770 sky130_fd_sc_hd__dlygate4sd3_1
X_22042_ clknet_leaf_92_i_clk net3668 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3512 net4069 vssd1 vssd1 vccd1 vccd1 net4036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4257 _00433_ vssd1 vssd1 vccd1 vccd1 net4781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4268 _01639_ vssd1 vssd1 vccd1 vccd1 net4792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3523 _00459_ vssd1 vssd1 vccd1 vccd1 net4047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4279 _01643_ vssd1 vssd1 vccd1 vccd1 net4803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3534 net4098 vssd1 vssd1 vccd1 vccd1 net4058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2800 _03821_ vssd1 vssd1 vccd1 vccd1 net3324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3545 gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 net4069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2811 _00416_ vssd1 vssd1 vccd1 vccd1 net3335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3556 _00462_ vssd1 vssd1 vccd1 vccd1 net4080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2822 rbzero.pov.ready_buffer\[16\] vssd1 vssd1 vccd1 vccd1 net3346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3567 _04825_ vssd1 vssd1 vccd1 vccd1 net4091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3578 rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 net4102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2833 net6144 vssd1 vssd1 vccd1 vccd1 net3357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2844 _01219_ vssd1 vssd1 vccd1 vccd1 net3368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3589 _00790_ vssd1 vssd1 vccd1 vccd1 net4113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 net6498 vssd1 vssd1 vccd1 vccd1 net3379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2866 _03816_ vssd1 vssd1 vccd1 vccd1 net3390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2877 _10078_ vssd1 vssd1 vccd1 vccd1 net3401 sky130_fd_sc_hd__buf_1
Xhold2888 net1314 vssd1 vssd1 vccd1 vccd1 net3412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2899 _03859_ vssd1 vssd1 vccd1 vccd1 net3423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21826_ clknet_leaf_91_i_clk net4409 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21757_ clknet_leaf_22_i_clk net1905 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11510_ rbzero.spi_registers.texadd2\[13\] _04679_ _04680_ rbzero.spi_registers.texadd0\[13\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _05219_ vssd1 vssd1 vccd1 vccd1 _05656_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21688_ clknet_leaf_29_i_clk net5059 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ _04165_ _04600_ _04611_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__or4_1
XFILLER_0_190_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20639_ _03083_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14160_ _06668_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__buf_2
X_11372_ net6948 net2711 _04562_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6160 net1797 vssd1 vssd1 vccd1 vccd1 net6684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _06257_ net4898 _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__and3_1
Xhold6171 rbzero.tex_b1\[17\] vssd1 vssd1 vccd1 vccd1 net6695 sky130_fd_sc_hd__dlygate4sd3_1
X_22309_ net441 net2378 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6182 net1678 vssd1 vssd1 vccd1 vccd1 net6706 sky130_fd_sc_hd__dlygate4sd3_1
X_14091_ _07207_ _07241_ _06865_ _07193_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__a2bb2o_1
Xhold6193 _04435_ vssd1 vssd1 vccd1 vccd1 net6717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5470 _00664_ vssd1 vssd1 vccd1 vccd1 net5994 sky130_fd_sc_hd__dlygate4sd3_1
X_13042_ _06195_ _06197_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__and2b_1
Xhold5481 net2905 vssd1 vssd1 vccd1 vccd1 net6005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5492 rbzero.map_overlay.i_othery\[0\] vssd1 vssd1 vccd1 vccd1 net6016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4780 net992 vssd1 vssd1 vccd1 vccd1 net5304 sky130_fd_sc_hd__dlygate4sd3_1
X_17850_ _01890_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4791 _00747_ vssd1 vssd1 vccd1 vccd1 net5315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16801_ _08755_ _09870_ _09790_ vssd1 vssd1 vccd1 vccd1 _09871_ sky130_fd_sc_hd__a21o_1
X_17781_ _01824_ _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__xnor2_1
X_14993_ net7458 _08102_ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19520_ _03000_ _03275_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__or2_1
X_16732_ _09800_ _09801_ vssd1 vssd1 vccd1 vccd1 _09802_ sky130_fd_sc_hd__nor2_1
X_13944_ _07087_ _07088_ _07093_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ net3256 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__clkbuf_1
X_16663_ _09732_ _09733_ _09096_ vssd1 vssd1 vccd1 vccd1 _09734_ sky130_fd_sc_hd__a21oi_1
X_13875_ _06826_ _06837_ _06933_ _06955_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__or4_4
XFILLER_0_186_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18402_ net4613 net4378 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__nor2_1
X_15614_ _08532_ _08530_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__nand2_1
X_12826_ net54 _05946_ _05956_ net55 vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19382_ net1537 _03199_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__or2_1
X_16594_ _09305_ _09486_ net7440 vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__or3b_1
XFILLER_0_9_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18333_ _10010_ _02372_ _10037_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15545_ _08612_ _08619_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__xor2_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ net4021 _05895_ _05903_ _05299_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a22o_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11708_ net4001 _04876_ net2705 _04605_ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a221o_1
X_15476_ _08347_ _08367_ _08542_ _08550_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__or4_2
X_18264_ _02306_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12688_ net4095 _05446_ net10 vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17215_ _10104_ _10105_ _10102_ vssd1 vssd1 vccd1 vccd1 _10216_ sky130_fd_sc_hd__a21oi_2
X_14427_ _07573_ _07577_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__nand2_2
X_11639_ net3936 net3929 net4001 net3 vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or4b_1
X_18195_ _02146_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__or3b_1
XFILLER_0_154_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17146_ _10129_ _10147_ vssd1 vssd1 vccd1 vccd1 _10148_ sky130_fd_sc_hd__xor2_2
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ net7757 net558 vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__nand2_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold706 net3659 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 net3669 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold728 net4465 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__nand2_1
X_17077_ _10019_ _09908_ vssd1 vssd1 vccd1 vccd1 _10080_ sky130_fd_sc_hd__nand2_1
Xhold739 net5519 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ _06859_ _07439_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _08449_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2107 net4798 vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2118 net7150 vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2129 net7001 vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1406 _04528_ vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 net5930 vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 _01381_ vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
X_17979_ _01836_ _01943_ _01833_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a21boi_1
Xhold1439 _01156_ vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20740__171 clknet_1_0__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__inv_2
X_19718_ net6164 _03393_ net2456 _03400_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__o211a_1
X_20990_ clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__buf_1
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19649_ net6854 _03362_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ clknet_leaf_22_i_clk net5400 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21542_ clknet_leaf_26_i_clk net1421 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21473_ clknet_leaf_0_i_clk net3071 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20424_ net3231 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20355_ clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__buf_1
XFILLER_0_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4010 net3015 vssd1 vssd1 vccd1 vccd1 net4534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4021 rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 net4545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4032 net3493 vssd1 vssd1 vccd1 vccd1 net4556 sky130_fd_sc_hd__buf_1
Xhold4043 net7460 vssd1 vssd1 vccd1 vccd1 net4567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4054 net7807 vssd1 vssd1 vccd1 vccd1 net4578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20286_ net1508 _03678_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3320 _03839_ vssd1 vssd1 vccd1 vccd1 net3844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4065 _01016_ vssd1 vssd1 vccd1 vccd1 net4589 sky130_fd_sc_hd__dlygate4sd3_1
X_20823__246 clknet_1_0__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__inv_2
X_22025_ clknet_leaf_97_i_clk net3452 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4076 rbzero.debug_overlay.facingY\[-1\] vssd1 vssd1 vccd1 vccd1 net4600 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3331 _02961_ vssd1 vssd1 vccd1 vccd1 net3855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4087 net2955 vssd1 vssd1 vccd1 vccd1 net4611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3342 _03300_ vssd1 vssd1 vccd1 vccd1 net3866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4098 _04150_ vssd1 vssd1 vccd1 vccd1 net4622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3353 _03619_ vssd1 vssd1 vccd1 vccd1 net3877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3364 _00625_ vssd1 vssd1 vccd1 vccd1 net3888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3375 net6331 vssd1 vssd1 vccd1 vccd1 net3899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2630 _00949_ vssd1 vssd1 vccd1 vccd1 net3154 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2641 _00606_ vssd1 vssd1 vccd1 vccd1 net3165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3386 _05332_ vssd1 vssd1 vccd1 vccd1 net3910 sky130_fd_sc_hd__buf_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2652 _03628_ vssd1 vssd1 vccd1 vccd1 net3176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3397 net6209 vssd1 vssd1 vccd1 vccd1 net3921 sky130_fd_sc_hd__clkbuf_4
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2663 _08222_ vssd1 vssd1 vccd1 vccd1 net3187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2674 net6305 vssd1 vssd1 vccd1 vccd1 net3198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 net5871 vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold66 _01562_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2685 net4457 vssd1 vssd1 vccd1 vccd1 net3209 sky130_fd_sc_hd__buf_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1951 net7035 vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _03223_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2696 _00522_ vssd1 vssd1 vccd1 vccd1 net3220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net3021 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net1793 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__inv_2
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1962 _01547_ vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 _00653_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1973 net7158 vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1984 net7200 vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10941_ net2738 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__clkbuf_1
Xhold1995 _04201_ vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13660_ _06809_ _06810_ _06743_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__a21oi_1
X_10872_ net2386 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _05207_ _05770_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21809_ clknet_leaf_10_i_clk net4290 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _06626_ _06649_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__or2_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _08404_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__buf_2
X_12542_ _05003_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__or2_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15261_ _06523_ _06524_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__and2_1
X_12473_ _05248_ _05638_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17000_ _10010_ _09286_ vssd1 vssd1 vccd1 vccd1 _10011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14212_ _07339_ _07341_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__or2_1
X_11424_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _08275_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _07291_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__nor2_2
X_11355_ net2620 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ _07223_ _07217_ _07221_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__or3_1
X_18951_ _02864_ net3085 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__nand2_1
X_11286_ net53 net2034 _04448_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__nor2_1
X_13025_ net3034 vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__inv_2
X_18882_ _02867_ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or2_1
X_20798__223 clknet_1_0__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__inv_2
X_17833_ _01881_ _01882_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17764_ _01685_ _01687_ _01683_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a21boi_1
X_14976_ _06664_ _08001_ _08004_ _08090_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19503_ net3050 _03275_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__or2_1
X_16715_ _09690_ _09658_ vssd1 vssd1 vccd1 vccd1 _09785_ sky130_fd_sc_hd__or2b_1
X_13927_ _07077_ _07075_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__xnor2_2
X_17695_ _09999_ _01745_ _01746_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or3_2
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19434_ net1631 _03225_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or2_1
X_16646_ _09588_ _09589_ vssd1 vssd1 vccd1 vccd1 _09717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13858_ _06963_ _06986_ _07007_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__nor3_1
XFILLER_0_187_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19365_ net2094 _03186_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__or2_1
X_12809_ net4043 _05957_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a211o_1
X_16577_ net7407 _09648_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__nor2_1
X_13789_ _06736_ _06861_ net79 _06918_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _02353_ _02356_ _01870_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ _08599_ _08602_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__nand2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19296_ net2090 _03147_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20770__197 clknet_1_1__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__inv_2
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18247_ _02217_ _02227_ _02225_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15459_ _08130_ _08137_ _08144_ vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__o21ai_1
Xhold6907 _06712_ vssd1 vssd1 vccd1 vccd1 net7431 sky130_fd_sc_hd__clkbuf_2
Xhold6918 net6134 vssd1 vssd1 vccd1 vccd1 net7442 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6929 rbzero.wall_tracer.trackDistX\[8\] vssd1 vssd1 vccd1 vccd1 net7453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18178_ _02219_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold503 net5325 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17129_ _08317_ _08548_ _08556_ _08331_ vssd1 vssd1 vccd1 vccd1 _10131_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold514 net5305 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold525 _01651_ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 net7449 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold547 net5468 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ net3585 _03679_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__or2_1
Xhold558 _01588_ vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 net6378 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ net3617 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__clkbuf_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1203 _03002_ vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__buf_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 net6613 vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1225 _01545_ vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 _04283_ vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 net6645 vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1258 _01427_ vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 net7724 vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__buf_1
XFILLER_0_212_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21525_ clknet_leaf_35_i_clk net5332 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21456_ clknet_leaf_31_i_clk net3888 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20407_ net3468 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21387_ clknet_leaf_54_i_clk _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ net7093 net7071 _04448_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20747__177 clknet_1_0__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__inv_2
XFILLER_0_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__clkbuf_4
X_11071_ net6964 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
X_20269_ net3812 _03756_ _03763_ _03761_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3150 rbzero.pov.ready_buffer\[3\] vssd1 vssd1 vccd1 vccd1 net3674 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22008_ clknet_leaf_100_i_clk net3593 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3161 _03806_ vssd1 vssd1 vccd1 vccd1 net3685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3172 _03856_ vssd1 vssd1 vccd1 vccd1 net3696 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3183 _03921_ vssd1 vssd1 vccd1 vccd1 net3707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3194 net671 vssd1 vssd1 vccd1 vccd1 net3718 sky130_fd_sc_hd__clkbuf_2
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2460 net6252 vssd1 vssd1 vccd1 vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2471 net7366 vssd1 vssd1 vccd1 vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
X_14830_ net7438 _07980_ _07493_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__o21a_2
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2482 rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 net3006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2493 net7792 vssd1 vssd1 vccd1 vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1770 _01466_ vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1781 net6773 vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
X_14761_ _07854_ _07911_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__xnor2_1
X_11973_ net3016 net1603 gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and3_1
Xhold1792 net7178 vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ _09570_ _09571_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__nand2_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ net2709 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__clkbuf_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06764_ _06766_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17480_ _10477_ _10478_ vssd1 vssd1 vccd1 vccd1 _10479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14692_ _07796_ _07838_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16431_ _09357_ _09382_ _09503_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ net6698 net2458 _04299_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
X_13643_ _06677_ _06767_ _06793_ _06717_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ net5939 _03065_ _03068_ _03061_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__o211a_1
X_16362_ _09434_ _09316_ _09315_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__a21o_1
X_13574_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__clkbuf_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ net2623 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__clkbuf_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _02115_ _02148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ net4081 net987 _05120_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__mux2_1
X_15313_ _08300_ _06162_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19081_ net2948 net2979 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__or2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _08615_ _08173_ _08607_ _08177_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__o31a_1
XFILLER_0_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18032_ _02016_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _05014_ vssd1 vssd1 vccd1 vccd1 _05622_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ net3507 _04818_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__or2_2
XFILLER_0_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11407_ net2409 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15175_ net3272 vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__inv_2
X_12387_ _05279_ _05551_ _05553_ _05244_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _07014_ _07018_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or2b_1
X_11338_ net6431 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19983_ net3874 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
X_20806__230 clknet_1_1__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__inv_2
XFILLER_0_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _07204_ _07206_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__a21oi_1
X_18934_ _04633_ _02916_ _02917_ _09933_ net3090 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a32o_1
X_11269_ net2320 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18865_ _02838_ _02849_ _02850_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ net4558 net4639 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__nand2_1
X_18796_ _02779_ _02780_ _02781_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17747_ _01763_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__xnor2_1
X_14959_ _08102_ _08103_ net7458 vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__mux2_1
X_17678_ _01727_ _01728_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19417_ net4118 _03211_ net598 _03220_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__o211a_1
X_16629_ _09698_ _09699_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20852__272 clknet_1_0__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__inv_2
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19348_ net5674 _03172_ _03183_ _03181_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7427 net6146 vssd1 vssd1 vccd1 vccd1 net7951 sky130_fd_sc_hd__dlygate4sd3_1
X_19279_ net5364 _03132_ _03144_ _03142_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__o211a_1
Xhold6704 rbzero.tex_g1\[51\] vssd1 vssd1 vccd1 vccd1 net7228 sky130_fd_sc_hd__dlygate4sd3_1
X_21310_ clknet_leaf_74_i_clk _00479_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold6715 net2743 vssd1 vssd1 vccd1 vccd1 net7239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6726 rbzero.tex_b1\[21\] vssd1 vssd1 vccd1 vccd1 net7250 sky130_fd_sc_hd__dlygate4sd3_1
X_22290_ net422 net1490 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold6737 rbzero.tex_r0\[26\] vssd1 vssd1 vccd1 vccd1 net7261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6748 net2750 vssd1 vssd1 vccd1 vccd1 net7272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6759 rbzero.tex_r0\[31\] vssd1 vssd1 vccd1 vccd1 net7283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold300 net630 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
X_21241_ clknet_leaf_65_i_clk _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold311 net5160 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 net4646 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 net3694 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold344 net5125 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
X_21172_ net4183 _04140_ _04141_ _09403_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a22o_1
Xhold355 net5084 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 rbzero.traced_texa\[-8\] vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 net5260 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20123_ net5571 _03679_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__or2_1
Xhold388 net5351 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 net7500 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20054_ net3449 _03613_ net4773 _03602_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__o211a_1
Xhold1000 net5709 vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 net6303 vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 net3099 vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 net5723 vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 _00941_ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 _01266_ vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 net5737 vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 net4864 vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _01333_ vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1099 net4728 vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10640_ net6373 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _05262_ vssd1 vssd1 vccd1 vccd1 _05478_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21508_ clknet_leaf_44_i_clk net1507 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12241_ net4666 _05371_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21439_ clknet_leaf_87_i_clk net3410 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12172_ _05335_ _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a21o_2
XFILLER_0_82_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11123_ net6892 net6640 _04437_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
X_16980_ _09987_ _09988_ _09989_ _09992_ vssd1 vssd1 vccd1 vccd1 _09993_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ net6574 net2550 _04404_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
X_15931_ _09002_ _09003_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_64_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ rbzero.wall_tracer.rayAddendX\[4\] _02658_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02659_ sky130_fd_sc_hd__mux2_1
X_15862_ _08909_ _08935_ _08936_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__a21oi_2
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _08641_ _08793_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__nor2_1
Xhold2290 _03510_ vssd1 vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14813_ _07839_ _07879_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__nor2_2
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ net7585 _02584_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _08865_ _08866_ _08861_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__a21o_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_102 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_102/HI o_rgb[16]
+ sky130_fd_sc_hd__conb_1
X_17532_ _10419_ _10420_ vssd1 vssd1 vccd1 vccd1 _10531_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_79_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_113 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_113/HI zeros[5] sky130_fd_sc_hd__conb_1
XFILLER_0_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _07774_ _07359_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__nor2_1
Xtop_ew_algofoogle_124 vssd1 vssd1 vccd1 vccd1 ones[0] top_ew_algofoogle_124/LO sky130_fd_sc_hd__conb_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ net1793 net2993 _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__or3_1
Xtop_ew_algofoogle_135 vssd1 vssd1 vccd1 vccd1 ones[11] top_ew_algofoogle_135/LO sky130_fd_sc_hd__conb_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _10446_ _10448_ vssd1 vssd1 vccd1 vccd1 _10462_ sky130_fd_sc_hd__or2_1
X_10907_ net2632 net5893 _04321_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11887_ _05004_ _05056_ _05035_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__o21a_1
X_14675_ _07823_ _07824_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_168_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19202_ net2951 net7327 _03084_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ _08180_ net77 vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10838_ net6674 net2376 _04288_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13626_ _06727_ _06667_ _06686_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_1__f__05840_ clknet_0__05840_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05840_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17394_ _10265_ _10266_ _10393_ vssd1 vssd1 vccd1 vccd1 _10394_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19133_ net4345 _03052_ net631 _03048_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ net7951 _08314_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__nand2_2
X_10769_ net6395 net1723 _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__mux2_1
X_13557_ _06565_ _06586_ _06689_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _05235_ _05671_ _05673_ _05061_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__o211a_1
X_19064_ net3070 _03009_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16276_ _09218_ _09220_ _09217_ vssd1 vssd1 vccd1 vccd1 _09350_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13488_ _06531_ _06543_ _06554_ _06635_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nor4_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18015_ _01874_ _02063_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12439_ net4303 _05062_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_17_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15227_ _08048_ net7464 _08295_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4609 _00837_ vssd1 vssd1 vccd1 vccd1 net5133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ net4716 _08117_ _08249_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__mux2_1
Xhold3908 net7741 vssd1 vssd1 vccd1 vccd1 net4432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20882__298 clknet_1_1__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__inv_2
Xhold3919 _03585_ vssd1 vssd1 vccd1 vccd1 net4443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14109_ _07013_ _07019_ _07259_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__a21bo_1
X_19966_ net3954 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__clkbuf_1
X_15089_ _08190_ _08209_ net3263 _01622_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18917_ rbzero.wall_tracer.rayAddendY\[6\] _09932_ _02901_ _04633_ vssd1 vssd1 vccd1
+ vccd1 _02902_ sky130_fd_sc_hd__a22o_1
X_19897_ _03521_ net1035 _03523_ _06226_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18848_ net1580 _02830_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or3_1
X_18779_ _02769_ _02772_ _08246_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21790_ clknet_leaf_11_i_clk net6012 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22411_ net163 net2474 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold7202 net7367 vssd1 vssd1 vccd1 vccd1 net7726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7213 rbzero.texu_hot\[3\] vssd1 vssd1 vccd1 vccd1 net7737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7224 rbzero.row_render.size\[6\] vssd1 vssd1 vccd1 vccd1 net7748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7235 _06725_ vssd1 vssd1 vccd1 vccd1 net7759 sky130_fd_sc_hd__clkbuf_2
X_22342_ net474 net1725 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
Xhold6501 rbzero.tex_r1\[62\] vssd1 vssd1 vccd1 vccd1 net7025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7246 net7554 vssd1 vssd1 vccd1 vccd1 net7770 sky130_fd_sc_hd__buf_2
Xhold6512 net2475 vssd1 vssd1 vccd1 vccd1 net7036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7257 net4381 vssd1 vssd1 vccd1 vccd1 net7781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6523 rbzero.tex_b0\[21\] vssd1 vssd1 vccd1 vccd1 net7047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7268 net4314 vssd1 vssd1 vccd1 vccd1 net7792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6534 net2010 vssd1 vssd1 vccd1 vccd1 net7058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6545 net2040 vssd1 vssd1 vccd1 vccd1 net7069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5800 net621 vssd1 vssd1 vccd1 vccd1 net6324 sky130_fd_sc_hd__dlygate4sd3_1
X_22273_ net405 net934 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
Xhold6556 _04258_ vssd1 vssd1 vccd1 vccd1 net7080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5811 net729 vssd1 vssd1 vccd1 vccd1 net6335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6567 net2383 vssd1 vssd1 vccd1 vccd1 net7091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5822 gpout5.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6578 _04342_ vssd1 vssd1 vccd1 vccd1 net7102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5833 net1135 vssd1 vssd1 vccd1 vccd1 net6357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5844 _04345_ vssd1 vssd1 vccd1 vccd1 net6368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6589 net2424 vssd1 vssd1 vccd1 vccd1 net7113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 net4941 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
X_21224_ clknet_leaf_51_i_clk _00393_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5855 net1093 vssd1 vssd1 vccd1 vccd1 net6379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold141 net4966 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5866 rbzero.tex_g0\[12\] vssd1 vssd1 vccd1 vccd1 net6390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5877 net1103 vssd1 vssd1 vccd1 vccd1 net6401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _03514_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5888 _04322_ vssd1 vssd1 vccd1 vccd1 net6412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 net4180 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5899 net1235 vssd1 vssd1 vccd1 vccd1 net6423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _03345_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 net4545 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
X_21155_ _04134_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__buf_1
Xhold196 net4642 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
X_20106_ net3825 _03664_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__or2_1
X_21086_ _04075_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20037_ net4776 _03613_ _03623_ _03602_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__o211a_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20859__278 clknet_1_0__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__inv_2
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _04945_ _04952_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ net4045 net4066 net4083 net4078 net22 net25 vssd1 vssd1 vccd1 vccd1 _05949_
+ sky130_fd_sc_hd__mux4_1
X_21988_ net213 net2504 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ net1500 net2968 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__xnor2_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14460_ _07604_ _07610_ _07602_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__o21a_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ net4092 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10623_ net5830 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__clkbuf_1
X_13411_ net6148 _06431_ _06545_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14391_ _07531_ _07540_ _07541_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16130_ _09203_ _09204_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__nand2_1
X_13342_ net6253 _06430_ _06414_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16061_ _09130_ _09135_ _09132_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__o21a_1
X_13273_ _06421_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__or2_4
XFILLER_0_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12224_ net4620 vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__clkbuf_4
X_15012_ net7457 _08078_ _08084_ _08150_ net6162 vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__a221o_1
X_19820_ net3075 net3960 _03459_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
X_12155_ net4037 net4009 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ net6379 net2740 _04426_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__mux2_1
X_19751_ net6047 _03392_ net2355 _03413_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__o211a_1
X_12086_ _05234_ _05254_ _05028_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16963_ net4922 _09966_ _09965_ _09978_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18702_ _02647_ net4587 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11037_ net6686 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__clkbuf_1
X_15914_ _08933_ _08948_ _08988_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19682_ net1859 _03375_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16894_ net4303 _09937_ _09938_ net1304 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18633_ net4752 _02639_ _02641_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__and3_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _08849_ _08665_ _08917_ _08918_ _08919_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__a32oi_4
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20918__331 clknet_1_1__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__inv_2
XFILLER_0_91_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ net6086 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__clkbuf_1
X_15776_ _08846_ _08848_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__a21o_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ net3857 net3135 _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17515_ _10512_ _10513_ vssd1 vssd1 vccd1 vccd1 _10514_ sky130_fd_sc_hd__and2_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _07875_ _07876_ _07877_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__nor3b_2
X_11939_ net7670 net7677 net7671 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__and3_1
X_18495_ net3075 _02497_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ _10217_ _10445_ vssd1 vssd1 vccd1 vccd1 _10446_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14658_ _07803_ _07807_ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_131_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _06697_ _06698_ _06669_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__a21oi_1
X_17377_ _10283_ _10288_ vssd1 vssd1 vccd1 vccd1 _10377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ _07696_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19116_ net5124 _03040_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__or2_1
X_16328_ _09301_ _09401_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__xor2_4
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5107 net1301 vssd1 vssd1 vccd1 vccd1 net5631 sky130_fd_sc_hd__dlygate4sd3_1
X_19047_ net6164 _02990_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__or2_1
X_16259_ _09331_ _09332_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__and2_1
Xhold5118 net1345 vssd1 vssd1 vccd1 vccd1 net5642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5129 _00757_ vssd1 vssd1 vccd1 vccd1 net5653 sky130_fd_sc_hd__dlygate4sd3_1
X_20964__373 clknet_1_0__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__inv_2
XFILLER_0_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4406 net3506 vssd1 vssd1 vccd1 vccd1 net4930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4417 gpout2.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4428 _01634_ vssd1 vssd1 vccd1 vccd1 net4952 sky130_fd_sc_hd__dlygate4sd3_1
X_20663__101 clknet_1_1__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__inv_2
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4439 _01621_ vssd1 vssd1 vccd1 vccd1 net4963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3705 net1657 vssd1 vssd1 vccd1 vccd1 net4229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3716 _00494_ vssd1 vssd1 vccd1 vccd1 net4240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3738 _00767_ vssd1 vssd1 vccd1 vccd1 net4262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3749 net1190 vssd1 vssd1 vccd1 vccd1 net4273 sky130_fd_sc_hd__dlygate4sd3_1
X_19949_ net668 _03480_ _03531_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21911_ clknet_leaf_90_i_clk net5195 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21842_ clknet_leaf_80_i_clk net3841 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_21773_ clknet_leaf_102_i_clk net1846 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20724_ clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__buf_1
XFILLER_0_59_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_6_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7010 rbzero.wall_tracer.trackDistY\[-4\] vssd1 vssd1 vccd1 vccd1 net7534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7021 rbzero.wall_tracer.trackDistY\[-8\] vssd1 vssd1 vccd1 vccd1 net7545 sky130_fd_sc_hd__dlygate4sd3_1
X_20586_ net3498 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6320 net2360 vssd1 vssd1 vccd1 vccd1 net6844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7065 _08321_ vssd1 vssd1 vccd1 vccd1 net7589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6331 rbzero.tex_g1\[20\] vssd1 vssd1 vccd1 vccd1 net6855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22325_ net457 net2646 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold6342 net2376 vssd1 vssd1 vccd1 vccd1 net6866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7087 _02819_ vssd1 vssd1 vccd1 vccd1 net7611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6353 rbzero.tex_g0\[50\] vssd1 vssd1 vccd1 vccd1 net6877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7098 rbzero.spi_registers.texadd3\[11\] vssd1 vssd1 vccd1 vccd1 net7622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6364 net2581 vssd1 vssd1 vccd1 vccd1 net6888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6375 _04233_ vssd1 vssd1 vccd1 vccd1 net6899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5630 rbzero.debug_overlay.playerX\[0\] vssd1 vssd1 vccd1 vccd1 net6154 sky130_fd_sc_hd__dlygate4sd3_1
X_22256_ net388 net2236 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold6386 net2137 vssd1 vssd1 vccd1 vccd1 net6910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5641 _00932_ vssd1 vssd1 vccd1 vccd1 net6165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6397 rbzero.tex_r0\[3\] vssd1 vssd1 vccd1 vccd1 net6921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5652 net3249 vssd1 vssd1 vccd1 vccd1 net6176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5663 _02735_ vssd1 vssd1 vccd1 vccd1 net6187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21207_ net4942 net6355 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__xnor2_1
Xhold5674 rbzero.debug_overlay.playerX\[-2\] vssd1 vssd1 vccd1 vccd1 net6198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4940 _00957_ vssd1 vssd1 vccd1 vccd1 net5464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5685 rbzero.debug_overlay.playerX\[3\] vssd1 vssd1 vccd1 vccd1 net6209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22187_ net319 net1946 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold4951 _01044_ vssd1 vssd1 vccd1 vccd1 net5475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5696 net3936 vssd1 vssd1 vccd1 vccd1 net6220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4962 rbzero.spi_registers.texadd2\[21\] vssd1 vssd1 vccd1 vccd1 net5486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4973 net1068 vssd1 vssd1 vccd1 vccd1 net5497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4984 _01040_ vssd1 vssd1 vccd1 vccd1 net5508 sky130_fd_sc_hd__dlygate4sd3_1
X_21138_ net4155 net4705 vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__xnor2_1
Xhold4995 rbzero.pov.spi_buffer\[23\] vssd1 vssd1 vccd1 vccd1 net5519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_205_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21069_ _04058_ _04059_ _04060_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__a21bo_1
X_13960_ _07085_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__xnor2_2
X_12911_ net52 net35 net34 _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__a31o_1
X_13891_ _07041_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15630_ net6123 _08314_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__nand2_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _05996_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__nand2_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15561_ _08624_ _08627_ _08635_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__nand3_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ net57 _05905_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a21o_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _09096_ net4954 _10300_ _10168_ vssd1 vssd1 vccd1 vccd1 _10301_ sky130_fd_sc_hd__or4_4
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _07661_ _07662_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__xnor2_2
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ net2895 vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__inv_2
X_18280_ _02275_ _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__xnor2_1
X_15492_ _08563_ _08566_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__nand2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _10230_ _10231_ vssd1 vssd1 vccd1 vccd1 _10232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14443_ _07525_ _07593_ net7757 vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__o21a_1
X_11655_ _04821_ net3279 net4090 net4010 _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a221o_1
XFILLER_0_182_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17162_ _09732_ _09733_ _09086_ vssd1 vssd1 vccd1 vccd1 _10164_ sky130_fd_sc_hd__a21oi_1
X_10606_ net47 net48 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__xor2_4
X_14374_ _07356_ _07521_ _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__nor3_1
X_11586_ _04755_ _04757_ _04727_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16113_ _09091_ _08454_ _09187_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13325_ net4406 net6304 vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__nor2_1
X_17093_ _08724_ _09537_ vssd1 vssd1 vccd1 vccd1 _10095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16044_ _09113_ _09115_ _09116_ _09118_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__o211a_1
X_13256_ net5491 _06394_ _06393_ _06408_ vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12207_ _05353_ _05359_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or2_2
X_13187_ _06297_ _06304_ _06307_ _06327_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__a41o_1
XFILLER_0_209_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19803_ _03440_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__buf_4
X_12138_ _04599_ _05305_ _05306_ _04807_ net4001 vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__o32a_1
X_17995_ _01812_ _10407_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12069_ _05068_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__or2_1
X_19734_ net1563 _03408_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__or2_1
X_16946_ _06204_ _06211_ net4901 _06391_ vssd1 vssd1 vccd1 vccd1 _09964_ sky130_fd_sc_hd__a211o_1
XFILLER_0_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19665_ net3096 _03360_ net1913 _03371_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__o211a_1
X_16877_ _09935_ vssd1 vssd1 vccd1 vccd1 _09936_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18616_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15828_ _08900_ _08901_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__xor2_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19596_ net5057 _03325_ _03333_ _03330_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__o211a_1
X_18547_ net4463 rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _02563_
+ sky130_fd_sc_hd__nand2_1
X_15759_ _08806_ _08830_ _08833_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_158_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18478_ _02497_ _02498_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17429_ _10292_ _10306_ _10304_ vssd1 vssd1 vccd1 vccd1 _10429_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20440_ _08275_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03998_ clknet_0__03998_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03998_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20371_ net3592 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22110_ net242 net2342 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold4203 net3332 vssd1 vssd1 vccd1 vccd1 net4727 sky130_fd_sc_hd__buf_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4214 net852 vssd1 vssd1 vccd1 vccd1 net4738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4225 _01026_ vssd1 vssd1 vccd1 vccd1 net4749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22041_ clknet_leaf_92_i_clk net3415 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4236 _00609_ vssd1 vssd1 vccd1 vccd1 net4760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4247 rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 net4771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3502 net3534 vssd1 vssd1 vccd1 vccd1 net4026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3513 _04598_ vssd1 vssd1 vccd1 vccd1 net4037 sky130_fd_sc_hd__clkbuf_2
Xhold4258 net3693 vssd1 vssd1 vccd1 vccd1 net4782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3524 gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 net4048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4269 net909 vssd1 vssd1 vccd1 vccd1 net4793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3535 _04804_ vssd1 vssd1 vccd1 vccd1 net4059 sky130_fd_sc_hd__clkbuf_4
Xhold2801 _03822_ vssd1 vssd1 vccd1 vccd1 net3325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3546 net4036 vssd1 vssd1 vccd1 vccd1 net4070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3557 rbzero.color_sky\[4\] vssd1 vssd1 vccd1 vccd1 net4081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 rbzero.pov.ready_buffer\[40\] vssd1 vssd1 vccd1 vccd1 net3336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2823 net3175 vssd1 vssd1 vccd1 vccd1 net3347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3568 _04841_ vssd1 vssd1 vccd1 vccd1 net4092 sky130_fd_sc_hd__buf_1
Xhold2834 _00418_ vssd1 vssd1 vccd1 vccd1 net3358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3579 net1451 vssd1 vssd1 vccd1 vccd1 net4103 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2845 net4498 vssd1 vssd1 vccd1 vccd1 net3369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2856 _00521_ vssd1 vssd1 vccd1 vccd1 net3380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2867 _01189_ vssd1 vssd1 vccd1 vccd1 net3391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2878 net4908 vssd1 vssd1 vccd1 vccd1 net3402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2889 _03861_ vssd1 vssd1 vccd1 vccd1 net3413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21825_ clknet_leaf_91_i_clk net4564 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_21756_ clknet_leaf_22_i_clk net1561 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21687_ clknet_leaf_28_i_clk net5238 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _04612_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20638_ net4002 _04802_ net4061 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11371_ net6808 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
X_20569_ net2944 net3812 _03911_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6150 net1841 vssd1 vssd1 vccd1 vccd1 net6674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6161 _04396_ vssd1 vssd1 vccd1 vccd1 net6685 sky130_fd_sc_hd__dlygate4sd3_1
X_22308_ net440 net1479 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _06263_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__nor2_1
Xhold6172 net1800 vssd1 vssd1 vccd1 vccd1 net6696 sky130_fd_sc_hd__dlygate4sd3_1
X_14090_ _07239_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6183 rbzero.tex_b1\[19\] vssd1 vssd1 vccd1 vccd1 net6707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6194 net1918 vssd1 vssd1 vccd1 vccd1 net6718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5460 rbzero.tex_g0\[35\] vssd1 vssd1 vccd1 vccd1 net5984 sky130_fd_sc_hd__dlygate4sd3_1
X_13041_ _06196_ _06179_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__xnor2_1
X_22239_ net371 net2006 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold5471 rbzero.floor_leak\[5\] vssd1 vssd1 vccd1 vccd1 net5995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5482 _00661_ vssd1 vssd1 vccd1 vccd1 net6006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5493 net2925 vssd1 vssd1 vccd1 vccd1 net6017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4770 rbzero.spi_registers.texadd0\[22\] vssd1 vssd1 vccd1 vccd1 net5294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4781 rbzero.spi_registers.texadd1\[1\] vssd1 vssd1 vccd1 vccd1 net5305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4792 net965 vssd1 vssd1 vccd1 vccd1 net5316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16800_ net3042 _09486_ _08609_ _09869_ vssd1 vssd1 vccd1 vccd1 _09870_ sky130_fd_sc_hd__a22o_2
XFILLER_0_121_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17780_ _01825_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__xnor2_1
X_14992_ _08120_ _08132_ _07993_ _08007_ _06690_ _06707_ vssd1 vssd1 vccd1 vccd1 _08133_
+ sky130_fd_sc_hd__mux4_2
X_20800__225 clknet_1_0__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__inv_2
X_16731_ _08326_ _09664_ _09666_ _09661_ vssd1 vssd1 vccd1 vccd1 _09801_ sky130_fd_sc_hd__o31a_1
XFILLER_0_156_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13943_ _07087_ _07088_ _07093_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__and3_1
X_19450_ _03088_ net3255 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__or2_1
X_16662_ net3420 _09304_ vssd1 vssd1 vccd1 vccd1 _09733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13874_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__xnor2_4
X_18401_ net4613 net4378 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15613_ _08671_ _08672_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__nand2_1
X_19381_ net4170 _03198_ net1133 _03194_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__o211a_1
X_12825_ _05975_ _05983_ net24 vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__mux2_1
X_16593_ _09661_ _09663_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18332_ _02368_ _02371_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__xnor2_1
X_15544_ _06211_ _08613_ _08618_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__and3_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ net20 _05912_ _05915_ net21 vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__and4b_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _02307_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__xnor2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ net4059 net2864 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xor2_1
X_15475_ _08548_ _08549_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ net14 net13 vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__and2b_1
X_17214_ _10124_ _10093_ vssd1 vssd1 vccd1 vccd1 _10215_ sky130_fd_sc_hd__or2b_1
X_14426_ _07567_ _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18194_ _02146_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__o21ba_1
X_11638_ _04803_ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17145_ _10136_ _10146_ vssd1 vssd1 vccd1 vccd1 _10147_ sky130_fd_sc_hd__xnor2_2
X_14357_ _07506_ _07507_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _04643_ _04687_ _04688_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold707 net5601 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ _06451_ _06455_ _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__and3_1
Xhold718 net4846 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ _10077_ _10076_ net3400 _10068_ vssd1 vssd1 vccd1 vccd1 _10079_ sky130_fd_sc_hd__o211a_1
Xhold729 net3704 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__buf_6
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16027_ _09083_ _09101_ vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__xor2_1
X_13239_ net4824 _06202_ _06393_ _06394_ net2388 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2108 net7228 vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2119 _01490_ vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1407 _01172_ vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 net5932 vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
X_17978_ _02025_ _02026_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__nand2_1
Xhold1429 net7003 vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19717_ net6195 _03395_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__or2_1
X_16929_ net3265 _09294_ vssd1 vssd1 vccd1 vccd1 _09947_ sky130_fd_sc_hd__xor2_2
X_20775__202 clknet_1_0__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__inv_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19648_ net1608 _03360_ net1653 _03354_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19579_ net1608 _03304_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
X_21610_ clknet_leaf_22_i_clk net5149 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21541_ clknet_leaf_28_i_clk net1311 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21472_ clknet_leaf_0_i_clk net3089 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20423_ _03814_ net3230 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4000 net3630 vssd1 vssd1 vccd1 vccd1 net4524 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4011 net7536 vssd1 vssd1 vccd1 vccd1 net4535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4022 net709 vssd1 vssd1 vccd1 vccd1 net4546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4033 net7408 vssd1 vssd1 vccd1 vccd1 net4557 sky130_fd_sc_hd__dlygate4sd3_1
X_20285_ net4868 _03675_ _03771_ _08276_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__o211a_1
Xhold4044 net3503 vssd1 vssd1 vccd1 vccd1 net4568 sky130_fd_sc_hd__buf_1
Xhold4055 net3492 vssd1 vssd1 vccd1 vccd1 net4579 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3310 _03848_ vssd1 vssd1 vccd1 vccd1 net3834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4066 net7557 vssd1 vssd1 vccd1 vccd1 net4590 sky130_fd_sc_hd__dlygate4sd3_1
X_22024_ clknet_leaf_98_i_clk net3232 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3321 _03840_ vssd1 vssd1 vccd1 vccd1 net3845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4077 _03615_ vssd1 vssd1 vccd1 vccd1 net4601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3332 _00619_ vssd1 vssd1 vccd1 vccd1 net3856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3343 _00836_ vssd1 vssd1 vccd1 vccd1 net3867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4088 net7526 vssd1 vssd1 vccd1 vccd1 net4612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4099 _01641_ vssd1 vssd1 vccd1 vccd1 net4623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3354 _03620_ vssd1 vssd1 vccd1 vccd1 net3878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3365 net7354 vssd1 vssd1 vccd1 vccd1 net3889 sky130_fd_sc_hd__buf_1
Xhold2620 rbzero.color_sky\[0\] vssd1 vssd1 vccd1 vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 net4402 vssd1 vssd1 vccd1 vccd1 net3155 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2642 net3473 vssd1 vssd1 vccd1 vccd1 net3166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3387 _00475_ vssd1 vssd1 vccd1 vccd1 net3911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2653 _03629_ vssd1 vssd1 vccd1 vccd1 net3177 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3398 _02957_ vssd1 vssd1 vccd1 vccd1 net3922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2664 net6261 vssd1 vssd1 vccd1 vccd1 net3188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1930 _01449_ vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2675 _00592_ vssd1 vssd1 vccd1 vccd1 net3199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net2093 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1941 net5873 vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold78 net4113 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2686 net4450 vssd1 vssd1 vccd1 vccd1 net3210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1952 _04291_ vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2697 net7530 vssd1 vssd1 vccd1 vccd1 net3221 sky130_fd_sc_hd__buf_1
Xhold1963 net7194 vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 net4237 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1974 _01450_ vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1985 _04494_ vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ net7034 net7213 _04344_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
Xhold1996 _01558_ vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ net7066 net2714 _04299_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
X_12610_ net42 _05772_ _05774_ net4077 vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a31o_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ clknet_leaf_90_i_clk net4360 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13590_ _06739_ _06740_ _06692_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__mux2_2
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _04988_ vssd1 vssd1 vccd1 vccd1 _05706_
+ sky130_fd_sc_hd__mux2_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21739_ clknet_leaf_24_i_clk net2457 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ rbzero.wall_tracer.visualWallDist\[-8\] _08334_ _08303_ vssd1 vssd1 vccd1
+ vccd1 _08335_ sky130_fd_sc_hd__mux2_1
X_12472_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _05218_ vssd1 vssd1 vccd1 vccd1 _05638_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20299__36 clknet_1_0__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14211_ _07297_ _07296_ _07346_ _07348_ _07349_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a32o_2
XFILLER_0_152_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ net4037 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__clkbuf_4
X_15191_ _08274_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11354_ net7223 net6822 _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14142_ _06985_ _07022_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11285_ net6475 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
X_14073_ _07217_ _07221_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18950_ _02864_ net3085 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5290 rbzero.tex_b1\[60\] vssd1 vssd1 vccd1 vccd1 net5814 sky130_fd_sc_hd__dlygate4sd3_1
X_17901_ _01948_ _01949_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and2_1
X_13024_ net2388 _06179_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18881_ net4634 net3807 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__and2_1
X_17832_ _10130_ _09805_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__nor2_1
X_17763_ _01811_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14975_ net4354 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__clkbuf_1
X_16714_ _09783_ vssd1 vssd1 vccd1 vccd1 _09784_ sky130_fd_sc_hd__buf_4
X_19502_ net5255 _03274_ _03276_ _03260_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13926_ _06846_ _06898_ _06864_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17694_ _01741_ _01744_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19433_ net5413 _03224_ _03231_ _03220_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__o211a_1
X_16645_ _09714_ _09715_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ _06963_ _06986_ _07007_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19364_ net4227 _03185_ net1656 _03181_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__o211a_1
X_12808_ net43 _05946_ _05956_ net46 vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__a22o_1
X_16576_ _09646_ _09647_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ _06844_ _06916_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__and2b_1
X_18315_ _02353_ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15527_ net4335 _06211_ _08601_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__o21a_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ net20 net19 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__and2b_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19295_ net5026 _03146_ _03153_ _03142_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18246_ _09375_ _09249_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15458_ _08530_ _08531_ _08532_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6908 rbzero.wall_tracer.trackDistX\[7\] vssd1 vssd1 vccd1 vccd1 net7432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _07558_ _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__nor2_1
X_18177_ _02222_ _02223_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ net4358 _08434_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17128_ _09695_ vssd1 vssd1 vccd1 vccd1 _10130_ sky130_fd_sc_hd__buf_2
Xhold504 net5327 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold515 net5307 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 net5416 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 net6366 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold548 net7712 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _09999_ _09641_ vssd1 vssd1 vccd1 vccd1 _10064_ sky130_fd_sc_hd__or2_1
Xhold559 net5727 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20070_ _03616_ net3616 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__or2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 net5785 vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 net6615 vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 net7015 vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 _01487_ vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 net6647 vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1259 rbzero.spi_registers.buf_texadd2\[16\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21524_ clknet_leaf_35_i_clk net5358 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21455_ clknet_leaf_31_i_clk net3907 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20406_ _03791_ net3467 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21386_ clknet_leaf_54_i_clk _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11070_ net6962 net2870 _04404_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__clkbuf_4
X_20268_ net4833 net4839 vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3140 net5671 vssd1 vssd1 vccd1 vccd1 net3664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3151 _03640_ vssd1 vssd1 vccd1 vccd1 net3675 sky130_fd_sc_hd__dlygate4sd3_1
X_22007_ clknet_leaf_100_i_clk net3644 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3162 _03807_ vssd1 vssd1 vccd1 vccd1 net3686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3173 _03857_ vssd1 vssd1 vccd1 vccd1 net3697 sky130_fd_sc_hd__dlygate4sd3_1
X_20199_ net5233 _03718_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or2_1
Xhold3184 _01237_ vssd1 vssd1 vccd1 vccd1 net3708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2450 net7326 vssd1 vssd1 vccd1 vccd1 net2974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3195 net6151 vssd1 vssd1 vccd1 vccd1 net3719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2461 net7726 vssd1 vssd1 vccd1 vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2472 _03092_ vssd1 vssd1 vccd1 vccd1 net2996 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 net4788 vssd1 vssd1 vccd1 vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2494 rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 net3018 sky130_fd_sc_hd__buf_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 net6053 vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1771 net6831 vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _07871_ _07870_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__and2b_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1782 _01501_ vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ net3016 net3868 net2986 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__o21a_1
Xhold1793 _04549_ vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _06861_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10923_ net7127 net2708 _04333_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _07791_ _07841_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__xnor2_2
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16430_ _09379_ _09381_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__nor2_1
X_13642_ _06616_ _06688_ _06770_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__a21o_1
X_10854_ net6439 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20912__326 clknet_1_1__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__inv_2
XFILLER_0_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _09253_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__inv_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ _06661_ _06713_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__xnor2_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ net7191 net6714 _04255_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
X_18100_ _02146_ _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__or2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _08312_ _08380_ _08382_ _08386_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__a2bb2o_4
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _05117_ _05620_ _05689_ _04909_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a2bb2o_1
X_19080_ net6047 net2842 net2980 _03022_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _08615_ _08173_ _08177_ _08607_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__nor4_4
XFILLER_0_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18031_ _08849_ _09784_ _01997_ _01995_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__o31a_1
X_15243_ _08310_ _08317_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__or2_2
X_12455_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _05072_ vssd1 vssd1 vccd1 vccd1 _05621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ net6984 net6461 _04584_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15174_ _08265_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12386_ _05229_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14125_ _07274_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__nand2_1
X_11337_ net6429 net2399 _04551_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19982_ _03261_ net3873 vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__or2_1
X_14056_ _07202_ _07203_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__nor2_1
X_18933_ _02914_ _02915_ _02912_ _02913_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o211ai_2
X_11268_ net6810 net6860 _04514_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13007_ _06098_ _06101_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__xor2_1
X_11199_ net1856 net5868 _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__mux2_1
X_18864_ _04633_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17815_ net4558 net4639 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18795_ net4799 _02778_ _04623_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a21oi_1
X_17746_ _01795_ _01796_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14958_ _07995_ _07991_ _08019_ vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__and3_1
XFILLER_0_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _07057_ net1998 _07059_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__a21oi_2
X_17677_ _01727_ _01728_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__nor2_1
X_14889_ _06678_ _08035_ _08038_ _06664_ vssd1 vssd1 vccd1 vccd1 _08039_ sky130_fd_sc_hd__a211o_1
X_16628_ _08707_ _09447_ vssd1 vssd1 vccd1 vccd1 _09699_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19416_ net2014 _03212_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16559_ _09559_ _09630_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__xnor2_1
X_19347_ net1883 _03173_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20887__303 clknet_1_0__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__inv_2
XFILLER_0_70_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19278_ net5038 _03133_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6705 net2632 vssd1 vssd1 vccd1 vccd1 net7229 sky130_fd_sc_hd__dlygate4sd3_1
X_18229_ _02236_ _02237_ _02244_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__o21a_1
Xhold6716 rbzero.tex_r1\[27\] vssd1 vssd1 vccd1 vccd1 net7240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6727 net2796 vssd1 vssd1 vccd1 vccd1 net7251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6738 net2851 vssd1 vssd1 vccd1 vccd1 net7262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6749 rbzero.tex_g0\[21\] vssd1 vssd1 vccd1 vccd1 net7273 sky130_fd_sc_hd__dlygate4sd3_1
X_21240_ clknet_leaf_64_i_clk _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold301 net7313 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold312 net5162 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold323 net5171 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 net4632 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
X_21171_ net4159 _04140_ _04141_ _09276_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold345 net7502 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold356 net5270 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 net7507 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
X_20122_ net5571 _03676_ net954 _03636_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__o211a_1
Xhold378 net5142 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 net4805 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20053_ _05401_ _03614_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__or2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1001 net5711 vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _00808_ vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _00916_ vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 net5725 vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1045 net5779 vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 net6057 vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__buf_1
XFILLER_0_139_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1078 net4866 vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 net6032 vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__buf_1
XFILLER_0_197_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21507_ clknet_leaf_15_i_clk net2727 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ _05401_ _05381_ _05402_ _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a211o_1
X_21438_ clknet_leaf_83_i_clk net4725 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_146_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _05335_ _05339_ _05326_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__o21bai_1
X_21369_ clknet_leaf_60_i_clk _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ net2272 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold890 _01075_ vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ net2663 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
X_15930_ _08514_ _08501_ _08899_ _08969_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__and4bb_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _08910_ _08934_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__nor2_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2280 net7257 vssd1 vssd1 vccd1 vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _08546_ _09251_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__nor2_1
X_20992__18 clknet_1_0__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _07881_ _07918_ _07961_ _07962_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__o31ai_2
Xhold2291 _00965_ vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _02590_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__xnor2_1
X_15792_ _08861_ _08865_ _08866_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__nand3_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _10409_ _10411_ _10408_ vssd1 vssd1 vccd1 vccd1 _10530_ sky130_fd_sc_hd__a21bo_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1590 _03401_ vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_103 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_103/HI o_rgb[17]
+ sky130_fd_sc_hd__conb_1
X_14743_ _07618_ _07524_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__nor2_1
Xtop_ew_algofoogle_114 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_114/HI zeros[6] sky130_fd_sc_hd__conb_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ net1600 _05124_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__or2_1
Xtop_ew_algofoogle_125 vssd1 vssd1 vccd1 vccd1 ones[1] top_ew_algofoogle_125/LO sky130_fd_sc_hd__conb_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_136 vssd1 vssd1 vccd1 vccd1 ones[12] top_ew_algofoogle_136/LO sky130_fd_sc_hd__conb_1
X_20836__257 clknet_1_1__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__inv_2
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10906_ net5991 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__clkbuf_1
X_17462_ _10458_ _10459_ _10333_ _10337_ vssd1 vssd1 vccd1 vccd1 _10461_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14674_ _07232_ _07774_ _07400_ _07438_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11886_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _05037_ vssd1 vssd1 vccd1 vccd1 _05056_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16413_ _08628_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__clkbuf_4
X_19201_ net5326 _03078_ _03099_ _03096_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ _06693_ _06694_ _06606_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__a21o_1
X_17393_ _10267_ _10268_ vssd1 vssd1 vccd1 vccd1 _10393_ sky130_fd_sc_hd__and2_1
X_10837_ net2476 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19132_ net824 _03053_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__or2_1
X_16344_ _09347_ _09324_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ _06692_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__clkbuf_4
X_10768_ _04243_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _05068_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19063_ net3070 net2843 _03015_ _03011_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16275_ _09210_ _09212_ _09209_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _06591_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__inv_2
XFILLER_0_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10699_ net6788 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__clkbuf_1
X_18014_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__xor2_2
X_15226_ rbzero.wall_tracer.rayAddendY\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] _08300_
+ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ net4303 _05062_ _05096_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15157_ _08256_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
X_12369_ _05069_ _05533_ _05535_ _05061_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__o211a_1
Xhold3909 net3173 vssd1 vssd1 vccd1 vccd1 net4433 sky130_fd_sc_hd__dlymetal6s2s_1
X_14108_ _07011_ _07020_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__or2_1
X_19965_ _08279_ net3953 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__and2_1
X_15088_ net3262 _08201_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ _07184_ _07183_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18916_ _02899_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__xnor2_1
X_19896_ _03470_ _03515_ _03478_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18847_ net3700 net4799 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18778_ _02769_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17729_ _08643_ _08795_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22410_ net162 net2576 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7214 net4383 vssd1 vssd1 vccd1 vccd1 net7738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22341_ net473 net1978 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6502 net2262 vssd1 vssd1 vccd1 vccd1 net7026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7247 _06717_ vssd1 vssd1 vccd1 vccd1 net7771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6513 rbzero.tex_b0\[56\] vssd1 vssd1 vccd1 vccd1 net7037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7258 _02364_ vssd1 vssd1 vccd1 vccd1 net7782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6524 net2203 vssd1 vssd1 vccd1 vccd1 net7048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7269 _02343_ vssd1 vssd1 vccd1 vccd1 net7793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6535 rbzero.tex_r0\[57\] vssd1 vssd1 vccd1 vccd1 net7059 sky130_fd_sc_hd__dlygate4sd3_1
X_22272_ net404 net1943 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
Xhold6546 rbzero.tex_g0\[5\] vssd1 vssd1 vccd1 vccd1 net7070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5812 rbzero.tex_b1\[6\] vssd1 vssd1 vccd1 vccd1 net6336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6557 net1977 vssd1 vssd1 vccd1 vccd1 net7081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6568 rbzero.tex_g0\[6\] vssd1 vssd1 vccd1 vccd1 net7092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5823 net1080 vssd1 vssd1 vccd1 vccd1 net6347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6579 net2311 vssd1 vssd1 vccd1 vccd1 net7103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5834 rbzero.tex_r1\[20\] vssd1 vssd1 vccd1 vccd1 net6358 sky130_fd_sc_hd__dlygate4sd3_1
X_21223_ clknet_leaf_60_i_clk _00392_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5845 net1062 vssd1 vssd1 vccd1 vccd1 net6369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 net4319 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5856 _04433_ vssd1 vssd1 vccd1 vccd1 net6380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 net4943 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5867 net1073 vssd1 vssd1 vccd1 vccd1 net6391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net4944 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 net6183 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5878 rbzero.tex_r0\[24\] vssd1 vssd1 vccd1 vccd1 net6402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5889 net1121 vssd1 vssd1 vccd1 vccd1 net6413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_1
X_21154_ _02488_ clknet_1_1__leaf__05840_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__and2_2
Xhold175 net4116 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
X_20941__352 clknet_1_0__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__inv_2
Xhold186 net4547 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 net7621 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
X_20105_ net3825 _03664_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_2_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21085_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20036_ _05403_ _03614_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21987_ net212 net1963 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11740_ net1257 net2158 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__nand2_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ net4091 _04830_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__or3_1
XFILLER_0_194_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20869_ clknet_1_1__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__buf_1
XFILLER_0_166_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13410_ _06547_ _06549_ _06539_ _06550_ _06541_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__a41o_2
X_10622_ net5828 net5824 _04170_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14390_ _07539_ _07537_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13341_ _06448_ _06487_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__xor2_4
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16060_ _09132_ _09134_ vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__nand2_1
X_13272_ rbzero.wall_tracer.rayAddendX\[-2\] _06422_ _06414_ vssd1 vssd1 vccd1 vccd1
+ _06423_ sky130_fd_sc_hd__mux2_4
XFILLER_0_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ _06734_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__clkbuf_4
X_12223_ net3699 _05374_ _05372_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1
+ vccd1 _05392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12154_ _04626_ _04817_ _04820_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__o22a_1
X_11105_ net1675 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
X_19750_ net6076 _03394_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__or2_1
X_12085_ _04978_ _05239_ _05243_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__o31a_1
X_16962_ _09973_ _09977_ vssd1 vssd1 vccd1 vccd1 _09978_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18701_ _02686_ _02692_ _02704_ _08246_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a31o_1
X_11036_ net6684 net2897 _04392_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__mux2_1
X_15913_ _08981_ _08986_ _08987_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__a21bo_1
X_16893_ net4271 _09937_ _09938_ net1189 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a22o_1
X_19681_ net1591 _03374_ net4224 _03371_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15844_ net3722 _08311_ _08305_ _08351_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__or4_1
X_18632_ net4752 _02639_ _02641_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a21oi_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _08849_ _08665_ _08811_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__and3_1
X_18563_ rbzero.wall_tracer.rayAddendX\[-2\] _02577_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ net4600 net3090 _06129_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__and3_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _10379_ _08705_ _10511_ vssd1 vssd1 vccd1 vccd1 _10513_ sky130_fd_sc_hd__o21ai_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07811_ _07836_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__xor2_1
X_11938_ _04999_ _04982_ _05022_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
X_18494_ _02501_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _10442_ _10444_ vssd1 vssd1 vccd1 vccd1 _10445_ sky130_fd_sc_hd__xor2_4
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _07799_ _07801_ _07802_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__a21o_1
X_11869_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _05014_ vssd1 vssd1 vccd1 vccd1 _05039_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13608_ _06606_ _06693_ _06694_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ _10264_ _10273_ _10272_ vssd1 vssd1 vccd1 vccd1 _10376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14588_ _07714_ _07737_ _07738_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__a21oi_2
X_20335__68 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16327_ _09398_ _09400_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19115_ net6005 _03037_ _03047_ _03048_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13539_ net7908 vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19046_ net6164 _02988_ _03005_ _02993_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__o211a_1
X_16258_ _08724_ _08708_ _09330_ vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5108 rbzero.spi_registers.texadd2\[4\] vssd1 vssd1 vccd1 vccd1 net5632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5119 _00756_ vssd1 vssd1 vccd1 vccd1 net5643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15209_ _04693_ net3623 net3509 vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4407 _04626_ vssd1 vssd1 vccd1 vccd1 net4931 sky130_fd_sc_hd__dlygate4sd3_1
X_16189_ _09262_ _09263_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__nor2_1
Xhold4418 net654 vssd1 vssd1 vccd1 vccd1 net4942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3706 net7721 vssd1 vssd1 vccd1 vccd1 net4230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3717 net1423 vssd1 vssd1 vccd1 vccd1 net4241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3728 net7516 vssd1 vssd1 vccd1 vccd1 net4252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3739 net593 vssd1 vssd1 vccd1 vccd1 net4263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19948_ _03560_ _03561_ _03476_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19879_ _03474_ _03504_ net3996 vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21910_ clknet_leaf_90_i_clk net5214 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_21841_ clknet_leaf_81_i_clk net950 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_21772_ clknet_leaf_5_i_clk net1568 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7000 rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1 vccd1 net7524 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_63_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold7011 net4484 vssd1 vssd1 vccd1 vccd1 net7535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7022 rbzero.wall_tracer.trackDistX\[-1\] vssd1 vssd1 vccd1 vccd1 net7546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7033 rbzero.wall_tracer.trackDistY\[-7\] vssd1 vssd1 vccd1 vccd1 net7557 sky130_fd_sc_hd__dlygate4sd3_1
X_20585_ _03924_ net3497 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7044 _06788_ vssd1 vssd1 vccd1 vccd1 net7568 sky130_fd_sc_hd__buf_1
Xhold6310 net2296 vssd1 vssd1 vccd1 vccd1 net6834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6321 rbzero.tex_b0\[54\] vssd1 vssd1 vccd1 vccd1 net6845 sky130_fd_sc_hd__dlygate4sd3_1
X_22324_ net456 net2847 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7066 _08322_ vssd1 vssd1 vccd1 vccd1 net7590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6332 net2240 vssd1 vssd1 vccd1 vccd1 net6856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7077 _02602_ vssd1 vssd1 vccd1 vccd1 net7601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6343 rbzero.tex_r1\[9\] vssd1 vssd1 vccd1 vccd1 net6867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7088 _02822_ vssd1 vssd1 vccd1 vccd1 net7612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6354 net1995 vssd1 vssd1 vccd1 vccd1 net6878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7099 rbzero.spi_registers.texadd0\[11\] vssd1 vssd1 vccd1 vccd1 net7623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6365 rbzero.tex_g1\[34\] vssd1 vssd1 vccd1 vccd1 net6889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5620 _08208_ vssd1 vssd1 vccd1 vccd1 net6144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5631 net3821 vssd1 vssd1 vccd1 vccd1 net6155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22255_ net387 net1682 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold6376 net2080 vssd1 vssd1 vccd1 vccd1 net6900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6387 rbzero.tex_b1\[35\] vssd1 vssd1 vccd1 vccd1 net6911 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_78_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold5642 net2072 vssd1 vssd1 vccd1 vccd1 net6166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6398 net2163 vssd1 vssd1 vccd1 vccd1 net6922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5653 _01249_ vssd1 vssd1 vccd1 vccd1 net6177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5664 _02737_ vssd1 vssd1 vccd1 vccd1 net6188 sky130_fd_sc_hd__dlygate4sd3_1
X_21206_ net4942 net65 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_1
Xhold5675 net3028 vssd1 vssd1 vccd1 vccd1 net6199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4930 rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 net5454 sky130_fd_sc_hd__dlygate4sd3_1
X_22186_ net318 net2130 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold4941 net2934 vssd1 vssd1 vccd1 vccd1 net5465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5686 net3921 vssd1 vssd1 vccd1 vccd1 net6210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4952 rbzero.spi_registers.texadd1\[3\] vssd1 vssd1 vccd1 vccd1 net5476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5697 rbzero.wall_tracer.rayAddendY\[-4\] vssd1 vssd1 vccd1 vccd1 net6221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4963 net1096 vssd1 vssd1 vccd1 vccd1 net5487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4974 _00678_ vssd1 vssd1 vccd1 vccd1 net5498 sky130_fd_sc_hd__dlygate4sd3_1
X_21137_ _09920_ _04121_ _04122_ _03083_ net4679 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a32o_1
Xhold4985 rbzero.wall_tracer.mapY\[10\] vssd1 vssd1 vccd1 vccd1 net5509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4996 net1263 vssd1 vssd1 vccd1 vccd1 net5520 sky130_fd_sc_hd__dlygate4sd3_1
X_21068_ net4173 net4546 vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__nand2_1
X_20019_ rbzero.debug_overlay.facingY\[-2\] net3833 _03594_ vssd1 vssd1 vccd1 vccd1
+ _03611_ sky130_fd_sc_hd__mux2_1
X_12910_ net34 net35 net51 vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__and3b_1
X_13890_ _07031_ _07039_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _05997_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and2_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15560_ _08630_ net7444 _08632_ _08634_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__o22ai_2
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ net54 _05895_ _05903_ net55 vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a22o_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _07366_ _07358_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__nor2_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ net3619 vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__inv_2
X_15491_ _08564_ _08424_ _08565_ _08449_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__o22ai_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _10228_ _10229_ vssd1 vssd1 vccd1 vccd1 _10231_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _07356_ _07524_ _07521_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__o21a_1
XFILLER_0_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11654_ _04801_ _04822_ _04823_ _04602_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17161_ _09863_ _09864_ _08584_ vssd1 vssd1 vccd1 vccd1 _10163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10605_ _04162_ net3993 _04165_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__and3b_2
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14373_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11585_ _04159_ _04666_ _04756_ _04714_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _08698_ _08701_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__nand2_1
X_20948__358 clknet_1_1__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__inv_2
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ net4406 net4787 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and2_1
X_17092_ _09849_ _09830_ vssd1 vssd1 vccd1 vccd1 _10094_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _09074_ _09117_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__and2_1
X_13255_ _06406_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12206_ rbzero.debug_overlay.facingY\[-3\] _05373_ _05374_ rbzero.debug_overlay.facingY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a22o_1
X_13186_ _06290_ _06341_ _06275_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__o21a_1
XFILLER_0_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19802_ net6111 _03443_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__or2_1
X_12137_ _05194_ _04759_ _05300_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_209_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17994_ _02041_ _02042_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19733_ net3088 _03407_ net2095 _03413_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12068_ rbzero.tex_r1\[35\] rbzero.tex_r1\[34\] _05077_ vssd1 vssd1 vccd1 vccd1 _05237_
+ sky130_fd_sc_hd__mux2_1
X_16945_ net4900 _09962_ _06203_ vssd1 vssd1 vccd1 vccd1 _09963_ sky130_fd_sc_hd__a21oi_1
X_11019_ net2771 net6485 _04310_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__mux2_1
X_19664_ net6285 _03362_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__or2_1
X_16876_ _04632_ _09930_ vssd1 vssd1 vccd1 vccd1 _09935_ sky130_fd_sc_hd__nor2_4
X_18615_ net3797 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
X_15827_ _08444_ _08501_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__or2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ net3940 _03327_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__or2_1
X_20693__128 clknet_1_0__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__inv_2
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15758_ _08831_ _08832_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__nand2_2
X_18546_ net4463 rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _02562_
+ sky130_fd_sc_hd__nor2_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14709_ _07825_ _07824_ _07823_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__a21o_1
X_15689_ _08529_ _08587_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__nor2_1
X_18477_ net3074 net3150 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__nor2_4
XFILLER_0_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17428_ _10414_ _10427_ vssd1 vssd1 vccd1 vccd1 _10428_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17359_ _08849_ _09306_ _10358_ vssd1 vssd1 vccd1 vccd1 _10359_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03997_ clknet_0__03997_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03997_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20370_ _08279_ net3591 vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19029_ net1572 _02990_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__or2_1
Xhold4204 rbzero.pov.ready_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net4728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4215 rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 net4739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4226 net1599 vssd1 vssd1 vccd1 vccd1 net4750 sky130_fd_sc_hd__dlygate4sd3_1
X_22040_ clknet_leaf_92_i_clk net3425 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4237 net3446 vssd1 vssd1 vccd1 vccd1 net4761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4248 net4690 vssd1 vssd1 vccd1 vccd1 net4772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3503 _04627_ vssd1 vssd1 vccd1 vccd1 net4027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3514 _05326_ vssd1 vssd1 vccd1 vccd1 net4038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4259 net686 vssd1 vssd1 vccd1 vccd1 net4783 sky130_fd_sc_hd__clkbuf_2
Xhold3525 net3868 vssd1 vssd1 vccd1 vccd1 net4049 sky130_fd_sc_hd__buf_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3536 _05193_ vssd1 vssd1 vccd1 vccd1 net4060 sky130_fd_sc_hd__buf_4
XFILLER_0_167_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2802 _01192_ vssd1 vssd1 vccd1 vccd1 net3326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3547 _05327_ vssd1 vssd1 vccd1 vccd1 net4071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3558 _05691_ vssd1 vssd1 vccd1 vccd1 net4082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2813 net845 vssd1 vssd1 vccd1 vccd1 net3337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 _03819_ vssd1 vssd1 vccd1 vccd1 net3348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3569 _04907_ vssd1 vssd1 vccd1 vccd1 net4093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2835 rbzero.pov.ready_buffer\[53\] vssd1 vssd1 vccd1 vccd1 net3359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2857 net4496 vssd1 vssd1 vccd1 vccd1 net3381 sky130_fd_sc_hd__buf_1
XFILLER_0_208_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2868 net7468 vssd1 vssd1 vccd1 vccd1 net3392 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2879 _04625_ vssd1 vssd1 vccd1 vccd1 net3403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21824_ clknet_leaf_87_i_clk net3789 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21755_ clknet_leaf_22_i_clk net5765 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21686_ clknet_leaf_29_i_clk net5228 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20637_ _04802_ net4061 _03971_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20314__49 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ net6806 net2030 _04562_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20568_ _08274_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__clkbuf_2
Xhold6140 net1674 vssd1 vssd1 vccd1 vccd1 net6664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6151 _04292_ vssd1 vssd1 vccd1 vccd1 net6675 sky130_fd_sc_hd__dlygate4sd3_1
X_22307_ net439 net2561 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6162 net1798 vssd1 vssd1 vccd1 vccd1 net6686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6173 rbzero.tex_r0\[13\] vssd1 vssd1 vccd1 vccd1 net6697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6184 net1838 vssd1 vssd1 vccd1 vccd1 net6708 sky130_fd_sc_hd__dlygate4sd3_1
X_20499_ _03858_ net3302 vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5450 _00659_ vssd1 vssd1 vccd1 vccd1 net5974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6195 rbzero.spi_registers.buf_texadd3\[4\] vssd1 vssd1 vccd1 vccd1 net6719 sky130_fd_sc_hd__dlygate4sd3_1
X_13040_ net4821 vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__inv_2
X_22238_ net370 net1743 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold5461 net1938 vssd1 vssd1 vccd1 vccd1 net5985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5472 net4076 vssd1 vssd1 vccd1 vccd1 net5996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5483 rbzero.pov.ready_buffer\[63\] vssd1 vssd1 vccd1 vccd1 net6007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5494 _00660_ vssd1 vssd1 vccd1 vccd1 net6018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4760 _00850_ vssd1 vssd1 vccd1 vccd1 net5284 sky130_fd_sc_hd__dlygate4sd3_1
X_21004__6 clknet_1_0__leaf__03773_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
Xhold4771 net919 vssd1 vssd1 vccd1 vccd1 net5295 sky130_fd_sc_hd__dlygate4sd3_1
X_22169_ net301 net2523 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold4782 net1038 vssd1 vssd1 vccd1 vccd1 net5306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4793 rbzero.spi_registers.buf_texadd0\[5\] vssd1 vssd1 vccd1 vccd1 net5317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14991_ _07583_ _07978_ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16730_ _09795_ _09799_ vssd1 vssd1 vccd1 vccd1 _09800_ sky130_fd_sc_hd__xor2_1
X_13942_ _07089_ _07091_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16661_ _09610_ _09489_ _09304_ vssd1 vssd1 vccd1 vccd1 _09732_ sky130_fd_sc_hd__a21o_2
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _06913_ _07023_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15612_ _08681_ _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__nand2_1
X_18400_ _02431_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__clkbuf_1
X_12824_ net26 _05979_ _05982_ _05973_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a22o_1
X_16592_ _09133_ _09662_ _09540_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__a21bo_1
X_19380_ net1638 _03199_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15543_ net3063 _08379_ _08609_ _08617_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__a22o_4
X_18331_ _02369_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__or2b_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ net4043 _05904_ _05913_ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18262_ _08643_ _09805_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__nor2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ net2823 vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__inv_2
X_15474_ net3065 _08327_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ net4045 net4066 net4083 net4078 net10 net13 vssd1 vssd1 vccd1 vccd1 _05847_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17213_ _10087_ _10200_ vssd1 vssd1 vccd1 vccd1 _10214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14425_ net7438 _07574_ _07575_ _07494_ _07566_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__o311a_2
XFILLER_0_154_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18193_ _02122_ _02124_ _02126_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__o21ba_1
X_11637_ net4059 _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__or2_1
XFILLER_0_182_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17144_ _10144_ _10145_ vssd1 vssd1 vccd1 vccd1 _10146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14356_ net3246 _07468_ _07465_ _07311_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11568_ _04715_ _04728_ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold708 net5250 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ _06456_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nor2_4
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17075_ _10068_ net3400 _10076_ _10077_ vssd1 vssd1 vccd1 vccd1 _10078_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold719 net3736 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14287_ _07405_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__xnor2_4
X_11499_ _04652_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__nand2_1
X_16026_ _09089_ _09099_ _09100_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__a21oi_1
X_13238_ _06392_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _06320_ net3554 _06324_ net3314 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__o22a_1
Xhold2109 net5894 vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1408 net7017 vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
X_17977_ _01836_ _02024_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__or2_1
Xhold1419 _01441_ vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19716_ net3112 _03393_ net5793 _03400_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16928_ net2807 _09294_ vssd1 vssd1 vccd1 vccd1 _09946_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19647_ net6602 _03362_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__or2_1
X_16859_ net4038 _09920_ vssd1 vssd1 vccd1 vccd1 _09922_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19578_ net5243 _03302_ _03321_ _03314_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18529_ net1076 _02528_ _02529_ net4479 _02546_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21540_ clknet_leaf_28_i_clk net1594 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21471_ clknet_leaf_0_i_clk net3039 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20422_ net3229 net1294 _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4001 _00513_ vssd1 vssd1 vccd1 vccd1 net4525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4012 net3054 vssd1 vssd1 vccd1 vccd1 net4536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4023 _01599_ vssd1 vssd1 vccd1 vccd1 net4547 sky130_fd_sc_hd__dlygate4sd3_1
X_20284_ net1302 _03678_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4034 net3472 vssd1 vssd1 vccd1 vccd1 net4558 sky130_fd_sc_hd__buf_1
XFILLER_0_105_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3300 _00615_ vssd1 vssd1 vccd1 vccd1 net3824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4045 net7834 vssd1 vssd1 vccd1 vccd1 net4569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3311 _03849_ vssd1 vssd1 vccd1 vccd1 net3835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4056 _08251_ vssd1 vssd1 vccd1 vccd1 net4580 sky130_fd_sc_hd__dlygate4sd3_1
X_22023_ clknet_leaf_98_i_clk net3326 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4067 net3542 vssd1 vssd1 vccd1 vccd1 net4591 sky130_fd_sc_hd__buf_1
Xhold3322 _01200_ vssd1 vssd1 vccd1 vccd1 net3846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4078 _01004_ vssd1 vssd1 vccd1 vccd1 net4602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3333 rbzero.debug_overlay.facingY\[0\] vssd1 vssd1 vccd1 vccd1 net3857 sky130_fd_sc_hd__clkbuf_2
Xhold4089 net3554 vssd1 vssd1 vccd1 vccd1 net4613 sky130_fd_sc_hd__buf_1
Xhold3344 net4048 vssd1 vssd1 vccd1 vccd1 net3868 sky130_fd_sc_hd__buf_2
Xhold2610 net4628 vssd1 vssd1 vccd1 vccd1 net3134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3355 _01006_ vssd1 vssd1 vccd1 vccd1 net3879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3366 _02971_ vssd1 vssd1 vccd1 vccd1 net3890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2621 _03085_ vssd1 vssd1 vccd1 vccd1 net3145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3377 net7343 vssd1 vssd1 vccd1 vccd1 net3901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2632 rbzero.pov.ready_buffer\[73\] vssd1 vssd1 vccd1 vccd1 net3156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3388 rbzero.spi_registers.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 net3912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2643 _08227_ vssd1 vssd1 vccd1 vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2654 _01012_ vssd1 vssd1 vccd1 vccd1 net3178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3399 net6218 vssd1 vssd1 vccd1 vccd1 net3923 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1920 _01396_ vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2665 rbzero.pov.ready_buffer\[5\] vssd1 vssd1 vccd1 vccd1 net3189 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2676 net3794 vssd1 vssd1 vccd1 vccd1 net3200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 net6194 vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1942 _01295_ vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 _03193_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2687 net3912 vssd1 vssd1 vccd1 vccd1 net3211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net5120 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1953 _01480_ vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2698 net684 vssd1 vssd1 vccd1 vccd1 net3222 sky130_fd_sc_hd__clkbuf_2
Xhold1964 _03381_ vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1975 net7232 vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1986 _01297_ vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1997 net7110 vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ net2683 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21807_ clknet_leaf_10_i_clk net6193 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12540_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _04989_ vssd1 vssd1 vccd1 vccd1 _05705_
+ sky130_fd_sc_hd__mux2_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21738_ clknet_leaf_24_i_clk net2089 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _05219_ vssd1 vssd1 vccd1 vccd1 _05637_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21669_ clknet_leaf_13_i_clk net899 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ _07355_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__and2b_1
X_11422_ net4036 vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15190_ net89 vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14141_ _07023_ _06913_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__or2b_1
X_11353_ _04403_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14072_ _07165_ _07222_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__xnor2_1
X_11284_ net6473 net2037 _04169_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5280 net5941 vssd1 vssd1 vccd1 vccd1 net5804 sky130_fd_sc_hd__dlygate4sd3_1
X_17900_ _01948_ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__nor2_1
X_13023_ _06178_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__clkbuf_4
Xhold5291 _04462_ vssd1 vssd1 vccd1 vccd1 net5815 sky130_fd_sc_hd__dlygate4sd3_1
X_18880_ net4634 net3807 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nor2_1
Xhold4590 net1278 vssd1 vssd1 vccd1 vccd1 net5114 sky130_fd_sc_hd__dlygate4sd3_1
X_17831_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__nand2_1
X_17762_ _01812_ _09484_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__nor2_1
X_14974_ net4353 _08117_ _08027_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19501_ net3112 _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or2_1
X_16713_ net4828 _09305_ _09486_ vssd1 vssd1 vccd1 vccd1 _09783_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _06966_ _06862_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nor2_8
XFILLER_0_89_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17693_ _01741_ _01744_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19432_ net1847 _03225_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644_ _09692_ _09713_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__or2_1
X_13856_ _06995_ _07006_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12807_ net44 _05958_ _05945_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__a21bo_1
X_19363_ net1655 _03186_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or2_1
X_16575_ _09521_ net3004 _09524_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13787_ _06915_ _06919_ _06917_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__a21o_1
X_10999_ net2479 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18314_ _02354_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15526_ _08311_ net7769 vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ net4045 net4066 net4083 net4078 net16 net19 vssd1 vssd1 vccd1 vccd1 _05898_
+ sky130_fd_sc_hd__mux4_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ net2274 _03147_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15457_ _08353_ _08373_ _08405_ _08422_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__or4_1
X_18245_ _02289_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ net3930 _05795_ _05799_ net3937 _05830_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14408_ _07548_ _07557_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__and2_1
Xhold6909 _06733_ vssd1 vssd1 vccd1 vccd1 net7433 sky130_fd_sc_hd__buf_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ _08318_ _08462_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__xnor2_4
X_18176_ _01778_ _09310_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17127_ _09852_ _09859_ _10128_ vssd1 vssd1 vccd1 vccd1 _10129_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ _07268_ _07468_ _07472_ _07489_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__a211o_1
Xhold505 net5412 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 net6370 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold527 net5418 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 net6368 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ _10058_ _10061_ _10019_ vssd1 vssd1 vccd1 vccd1 _10063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 net6390 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16009_ _08587_ _08874_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__or2_1
X_20998__24 clknet_1_1__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_0_110_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 net6621 vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _01162_ vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
X_20699__134 clknet_1_1__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__inv_2
XFILLER_0_139_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _04445_ vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1238 rbzero.tex_r1\[39\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _01411_ vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21523_ clknet_leaf_34_i_clk net2998 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21454_ clknet_leaf_31_i_clk net3916 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20405_ net1298 net3466 _03801_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__mux2_1
X_21385_ clknet_leaf_56_i_clk _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 o_gpout[0] sky130_fd_sc_hd__buf_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__clkbuf_4
X_20267_ net4833 _03756_ _03762_ _03761_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__o211a_1
Xhold3130 _01203_ vssd1 vssd1 vccd1 vccd1 net3654 sky130_fd_sc_hd__dlygate4sd3_1
X_22006_ clknet_leaf_99_i_clk net3271 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3141 net1370 vssd1 vssd1 vccd1 vccd1 net3665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3152 _03641_ vssd1 vssd1 vccd1 vccd1 net3676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3163 _01185_ vssd1 vssd1 vccd1 vccd1 net3687 sky130_fd_sc_hd__dlygate4sd3_1
X_20198_ net5233 _03717_ _03723_ _03722_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__o211a_1
Xhold3174 _01208_ vssd1 vssd1 vccd1 vccd1 net3698 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2440 rbzero.spi_registers.buf_sky\[2\] vssd1 vssd1 vccd1 vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3185 rbzero.pov.ready_buffer\[32\] vssd1 vssd1 vccd1 vccd1 net3709 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2451 _03098_ vssd1 vssd1 vccd1 vccd1 net2975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3196 _00430_ vssd1 vssd1 vccd1 vccd1 net3720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2462 net4890 vssd1 vssd1 vccd1 vccd1 net2986 sky130_fd_sc_hd__buf_2
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2473 _03093_ vssd1 vssd1 vccd1 vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2484 net6129 vssd1 vssd1 vccd1 vccd1 net3008 sky130_fd_sc_hd__clkbuf_2
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2495 net6320 vssd1 vssd1 vccd1 vccd1 net3019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1750 net6729 vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1761 net6971 vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _04776_ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__or2_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1772 net6833 vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1783 net7172 vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1794 _01153_ vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__clkbuf_4
X_10922_ net5846 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14690_ _07790_ _07840_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__nor2_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13641_ _06662_ _06791_ _06589_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__a21o_1
XFILLER_0_212_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10853_ net6437 net2063 _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _09423_ _09432_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13572_ _06591_ _06595_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10784_ net2170 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__clkbuf_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _08381_ _08385_ _08327_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ _05654_ _05688_ _04975_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__mux2_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _08626_ _09364_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15242_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__clkbuf_4
X_18030_ _02018_ _01987_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or2b_1
X_12454_ net3378 _05448_ _05617_ _05208_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ net2216 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
X_15173_ net4417 _08160_ _08260_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__mux2_1
X_12385_ rbzero.tex_g1\[35\] rbzero.tex_g1\[34\] _05262_ vssd1 vssd1 vccd1 vccd1 _05552_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14124_ _07262_ _07263_ _07273_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__nand3_1
X_11336_ net1825 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
X_19981_ rbzero.debug_overlay.facingX\[-5\] net3519 _03581_ vssd1 vssd1 vccd1 vccd1
+ _03587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _07205_ _06869_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nor2_1
X_18932_ _02912_ _02913_ _02914_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a211o_1
X_11267_ net2859 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
X_13006_ _06160_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18863_ _02838_ _02850_ _02849_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a21o_1
X_11198_ _04332_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17814_ _01864_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ net4799 net4640 _05393_ net4438 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17745_ _01695_ _01764_ _01794_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__nand3_1
X_14957_ _08082_ _08101_ _08069_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__mux2_1
X_13908_ _07044_ _07056_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17676_ _10505_ _10557_ _10555_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a21oi_1
X_14888_ _06678_ _08036_ _08037_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__nor3_1
XFILLER_0_187_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19415_ net4999 _03211_ _03221_ _03220_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16627_ _09696_ _09697_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__or2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _06929_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ net5633 _03172_ _03182_ _03181_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__o211a_1
X_16558_ _09627_ _09629_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15509_ _08559_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19277_ net5295 _03132_ _03143_ _03142_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__o211a_1
X_16489_ _09464_ _09473_ _09472_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7418 rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 net7942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18228_ _02272_ _02273_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__xnor2_1
Xhold6706 _04329_ vssd1 vssd1 vccd1 vccd1 net7230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6717 net2556 vssd1 vssd1 vccd1 vccd1 net7241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6728 rbzero.tex_b1\[15\] vssd1 vssd1 vccd1 vccd1 net7252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6739 rbzero.tex_b0\[5\] vssd1 vssd1 vccd1 vccd1 net7263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18159_ _02108_ _02090_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or2b_1
Xhold302 net5116 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold313 net5086 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 net5173 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
X_21170_ net4190 _04140_ _04141_ _09281_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold335 net5167 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 net5177 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 net5272 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20121_ net5598 _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__or2_1
Xhold368 net5157 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03779_ _03779_ vssd1 vssd1 vccd1 vccd1 clknet_0__03779_ sky130_fd_sc_hd__clkbuf_16
Xhold379 net5144 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20707__141 clknet_1_0__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__inv_2
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20052_ net3244 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__clkbuf_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 net6542 vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 net7658 vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 net6042 vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 net6297 vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 net5781 vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 net7627 vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1068 net4225 vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 net4274 vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__buf_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20753__183 clknet_1_1__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__inv_2
XFILLER_0_181_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21506_ clknet_leaf_44_i_clk net2792 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21437_ clknet_leaf_83_i_clk net3165 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ net4004 _05338_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21368_ clknet_leaf_60_i_clk _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ net7050 net6892 _04437_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__mux2_1
X_21299_ clknet_leaf_43_i_clk _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold880 net5673 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 net5689 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ net7245 net6574 _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _08910_ _08934_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__xor2_2
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2270 _04592_ vssd1 vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2281 _04570_ vssd1 vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14811_ _07882_ _07917_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__nand2_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2292 net7184 vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _08458_ _08864_ _08863_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__a21o_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1580 net6779 vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _10506_ _10528_ vssd1 vssd1 vccd1 vccd1 _10529_ sky130_fd_sc_hd__xnor2_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _07232_ _07354_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__or2_1
X_11954_ _05122_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nand2_1
Xhold1591 _00905_ vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_104 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_104/HI o_rgb[18]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_115 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_115/HI zeros[7] sky130_fd_sc_hd__conb_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_126 vssd1 vssd1 vccd1 vccd1 ones[2] top_ew_algofoogle_126/LO sky130_fd_sc_hd__conb_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_137 vssd1 vssd1 vccd1 vccd1 ones[13] top_ew_algofoogle_137/LO sky130_fd_sc_hd__conb_1
XFILLER_0_212_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10905_ net5893 net5989 _04321_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17461_ _10333_ _10337_ _10458_ _10459_ vssd1 vssd1 vccd1 vccd1 _10460_ sky130_fd_sc_hd__a211oi_1
X_14673_ _07774_ _07400_ _07439_ _07232_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__o22ai_2
X_11885_ _04984_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19200_ net1615 _03079_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16412_ _09096_ _09484_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13624_ _06676_ _06773_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10836_ net7036 net6674 _04288_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__mux2_1
X_17392_ _10390_ _10391_ vssd1 vssd1 vccd1 vccd1 _10392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19131_ net5950 _03052_ _03057_ _03048_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__o211a_1
X_16343_ _09323_ _09392_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__nand2_1
X_13555_ _06663_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__or2_1
X_10767_ net2419 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _05071_ vssd1 vssd1 vccd1 vccd1 _05672_
+ sky130_fd_sc_hd__mux2_1
X_16274_ _09324_ _09347_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__xnor2_1
X_19062_ net3088 _03009_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13486_ _06622_ _06634_ _06636_ _06616_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__and4b_1
X_10698_ net2007 net6786 _04214_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18013_ _01876_ _01956_ _01955_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a21oi_2
X_15225_ net4086 vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__clkbuf_4
X_12437_ _05105_ _05115_ _05103_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__or3b_1
XFILLER_0_113_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15156_ net4399 _08106_ _08249_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12368_ _05248_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14107_ _07071_ _07155_ _07254_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__a2bb2o_4
X_11319_ net2347 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19964_ net3952 _03569_ _03574_ _03529_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a22o_1
X_15087_ net4560 net4491 _08191_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__mux2_1
X_12299_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _05218_ vssd1 vssd1 vccd1 vccd1 _05467_
+ sky130_fd_sc_hd__mux2_1
X_14038_ _07188_ _07186_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__xnor2_1
X_18915_ _02867_ _02885_ _02887_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
X_19895_ net1034 _03485_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18846_ _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18777_ _02770_ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__or2b_1
X_15989_ _08424_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17728_ _10259_ _01778_ _01676_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17659_ _10168_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__buf_2
XFILLER_0_203_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19329_ _03084_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7215 rbzero.texu_hot\[2\] vssd1 vssd1 vccd1 vccd1 net7739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22340_ net472 net2850 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
Xhold7226 rbzero.wall_tracer.trackDistX\[10\] vssd1 vssd1 vccd1 vccd1 net7750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7237 _08335_ vssd1 vssd1 vccd1 vccd1 net7761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6503 rbzero.tex_g0\[36\] vssd1 vssd1 vccd1 vccd1 net7027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6514 net2160 vssd1 vssd1 vccd1 vccd1 net7038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6525 rbzero.tex_g0\[15\] vssd1 vssd1 vccd1 vccd1 net7049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22271_ net403 net2398 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
Xhold6536 net2505 vssd1 vssd1 vccd1 vccd1 net7060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6547 net1926 vssd1 vssd1 vccd1 vccd1 net7071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5802 _02625_ vssd1 vssd1 vccd1 vccd1 net6326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5813 net760 vssd1 vssd1 vccd1 vccd1 net6337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6558 rbzero.tex_g0\[25\] vssd1 vssd1 vccd1 vccd1 net7082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6569 net2616 vssd1 vssd1 vccd1 vccd1 net7093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5824 gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5835 net995 vssd1 vssd1 vccd1 vccd1 net6359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold110 net6317 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
X_21222_ clknet_leaf_58_i_clk _00391_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold121 rbzero.wall_tracer.visualWallDist\[-4\] vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_2
Xhold5846 rbzero.tex_r1\[50\] vssd1 vssd1 vccd1 vccd1 net6370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 rbzero.wall_tracer.visualWallDist\[-1\] vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_1
Xhold5857 net1094 vssd1 vssd1 vccd1 vccd1 net6381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5868 _04444_ vssd1 vssd1 vccd1 vccd1 net6392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 net4946 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5879 net1159 vssd1 vssd1 vccd1 vccd1 net6403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 rbzero.wall_tracer.visualWallDist\[7\] vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_1
Xhold165 net4156 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
X_21153_ _09486_ net3981 _04133_ _01622_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__o31a_1
Xhold176 net7483 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold187 net4394 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ net3330 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__clkbuf_1
Xhold198 net4522 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
X_21084_ _04075_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20035_ net3545 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ net211 net1388 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _04832_ _04833_ _04835_ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__or4_1
X_20868_ clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__buf_1
XFILLER_0_138_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10621_ net5826 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _06430_ _06151_ _06490_ _04635_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_10_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__mux2_4
X_22469_ clknet_leaf_79_i_clk net4808 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15010_ _08122_ _08148_ _08092_ vssd1 vssd1 vccd1 vccd1 _08149_ sky130_fd_sc_hd__mux2_2
X_12222_ net4625 vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__buf_2
XFILLER_0_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _04858_ _05296_ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a21oi_1
X_11104_ net6664 net6379 _04426_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12084_ _05244_ _05247_ _05252_ _05022_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a211o_1
X_16961_ net4875 _09975_ _09976_ vssd1 vssd1 vccd1 vccd1 _09977_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18700_ _02686_ _02692_ _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a21oi_1
X_11035_ net2660 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__clkbuf_1
X_15912_ _08967_ _08980_ _08949_ _08950_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__o211ai_2
X_19680_ net4223 _03375_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__or2_1
X_16892_ net4239 _09937_ _09938_ net1422 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18631_ _02605_ _02616_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a21o_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _08372_ _08632_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__or2_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _02569_ _02570_ _02576_ _04624_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _08351_ _08352_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__nand2_8
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12986_ net3876 net3085 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__nor2_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _10379_ _08705_ _10511_ vssd1 vssd1 vccd1 vccd1 _10512_ sky130_fd_sc_hd__or3_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _07814_ _07833_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__xnor2_1
X_11937_ _05104_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__nand2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ net3960 net3925 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__and2b_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _10219_ _10319_ _10443_ vssd1 vssd1 vccd1 vccd1 _10444_ sky130_fd_sc_hd__a21oi_2
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11868_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _05037_ vssd1 vssd1 vccd1 vccd1 _05038_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14656_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__and2b_1
XFILLER_0_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10819_ net6796 net6744 _04277_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__mux2_1
X_13607_ _06730_ _06757_ _06676_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__a21oi_1
X_17375_ _10343_ _10374_ vssd1 vssd1 vccd1 vccd1 _10375_ sky130_fd_sc_hd__xnor2_2
X_11799_ _04914_ _04917_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__o21a_1
X_14587_ _07715_ _07736_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19114_ _02992_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__clkbuf_4
X_16326_ _08802_ _09267_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13538_ _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19045_ net3112 _02990_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__or2_1
X_16257_ _08724_ _08707_ _09330_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__or3_1
X_13469_ _06540_ net82 _06424_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__o21a_2
XFILLER_0_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5109 net1368 vssd1 vssd1 vccd1 vccd1 net5633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ net3508 _06384_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16188_ _08742_ _09248_ _09261_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__and3_1
X_20925__337 clknet_1_0__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__inv_2
Xhold4408 _08247_ vssd1 vssd1 vccd1 vccd1 net4932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4419 _01646_ vssd1 vssd1 vccd1 vccd1 net4943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15139_ _06386_ net2960 net4829 _08239_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3707 net1500 vssd1 vssd1 vccd1 vccd1 net4231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3718 rbzero.spi_registers.buf_texadd2\[11\] vssd1 vssd1 vccd1 vccd1 net4242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3729 net774 vssd1 vssd1 vccd1 vccd1 net4253 sky130_fd_sc_hd__dlygate4sd3_1
X_19947_ net3880 _03553_ net4387 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19878_ net2812 _03485_ _03474_ _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18829_ net4708 rbzero.wall_tracer.rayAddendY\[1\] vssd1 vssd1 vccd1 vccd1 _02819_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21840_ clknet_leaf_81_i_clk net4449 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20819__242 clknet_1_1__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__inv_2
XFILLER_0_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21771_ clknet_leaf_5_i_clk net1545 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20971__379 clknet_1_1__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__inv_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20670__107 clknet_1_1__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__inv_2
XFILLER_0_72_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7001 rbzero.wall_tracer.trackDistX\[3\] vssd1 vssd1 vccd1 vccd1 net7525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7012 rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1 vccd1 net7536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7023 net4594 vssd1 vssd1 vccd1 vccd1 net7547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20584_ net2812 net3496 net3250 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
Xhold7034 rbzero.wall_tracer.trackDistX\[0\] vssd1 vssd1 vccd1 vccd1 net7558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6300 net2107 vssd1 vssd1 vccd1 vccd1 net6824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7045 rbzero.traced_texa\[2\] vssd1 vssd1 vccd1 vccd1 net7569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6311 rbzero.tex_g1\[25\] vssd1 vssd1 vccd1 vccd1 net6835 sky130_fd_sc_hd__dlygate4sd3_1
X_22323_ net455 net1155 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7056 _02890_ vssd1 vssd1 vccd1 vccd1 net7580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6322 net2146 vssd1 vssd1 vccd1 vccd1 net6846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6333 _04364_ vssd1 vssd1 vccd1 vccd1 net6857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7078 _02605_ vssd1 vssd1 vccd1 vccd1 net7602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6344 net1900 vssd1 vssd1 vccd1 vccd1 net6868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7089 rbzero.wall_tracer.rayAddendX\[-9\] vssd1 vssd1 vccd1 vccd1 net7613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6355 rbzero.tex_r1\[13\] vssd1 vssd1 vccd1 vccd1 net6879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5610 net3633 vssd1 vssd1 vccd1 vccd1 net6134 sky130_fd_sc_hd__buf_1
X_22254_ net386 net1699 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold6366 net2125 vssd1 vssd1 vccd1 vccd1 net6890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5621 rbzero.spi_registers.spi_buffer\[18\] vssd1 vssd1 vccd1 vccd1 net6145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6377 rbzero.tex_r1\[61\] vssd1 vssd1 vccd1 vccd1 net6901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5632 _00964_ vssd1 vssd1 vccd1 vccd1 net6156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6388 net2227 vssd1 vssd1 vccd1 vccd1 net6912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5643 rbzero.trace_state\[2\] vssd1 vssd1 vccd1 vccd1 net6167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5654 net2939 vssd1 vssd1 vccd1 vccd1 net6178 sky130_fd_sc_hd__dlygate4sd3_1
X_20865__284 clknet_1_1__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__inv_2
Xhold6399 rbzero.tex_g0\[31\] vssd1 vssd1 vccd1 vccd1 net6923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4920 rbzero.pov.spi_buffer\[49\] vssd1 vssd1 vccd1 vccd1 net5444 sky130_fd_sc_hd__dlygate4sd3_1
X_21205_ _03502_ net1921 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5665 _02738_ vssd1 vssd1 vccd1 vccd1 net6189 sky130_fd_sc_hd__dlygate4sd3_1
X_22185_ net317 net2362 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5676 _00962_ vssd1 vssd1 vccd1 vccd1 net6200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4931 net1016 vssd1 vssd1 vccd1 vccd1 net5455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4942 rbzero.pov.ready vssd1 vssd1 vccd1 vccd1 net5466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5687 _00967_ vssd1 vssd1 vccd1 vccd1 net6211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5698 net2884 vssd1 vssd1 vccd1 vccd1 net6222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4953 net1078 vssd1 vssd1 vccd1 vccd1 net5477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4964 _00775_ vssd1 vssd1 vccd1 vccd1 net5488 sky130_fd_sc_hd__dlygate4sd3_1
X_21136_ _04120_ _04119_ _04118_ _04115_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__a211o_1
Xhold4975 rbzero.pov.spi_buffer\[16\] vssd1 vssd1 vccd1 vccd1 net5499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4986 net1064 vssd1 vssd1 vccd1 vccd1 net5510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4997 _01059_ vssd1 vssd1 vccd1 vccd1 net5521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21067_ net4173 net4546 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or2_1
X_20018_ net888 _03578_ net4419 _03602_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__o211a_1
X_12840_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nor2_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _05922_ _05930_ net18 vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__mux2_1
X_21969_ net194 net2297 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14510_ _07367_ _07353_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__or2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _04882_ _04885_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__and3b_1
XFILLER_0_189_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15490_ _08557_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _07587_ _07591_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__nand2_1
X_11653_ net4090 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__inv_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ net4053 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__clkbuf_4
X_17160_ _08587_ _09861_ vssd1 vssd1 vccd1 vccd1 _10162_ sky130_fd_sc_hd__nor2_1
X_14372_ _07306_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__or2_2
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11584_ _04665_ _04658_ _04663_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__nand3_1
XFILLER_0_107_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16111_ _08572_ _08533_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13323_ net4561 net7146 _06465_ _06468_ _06466_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17091_ _09807_ _09824_ _09822_ vssd1 vssd1 vccd1 vccd1 _10093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16042_ _09067_ _09073_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__nand2_1
X_13254_ _06401_ _06404_ _06399_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ _05341_ _05343_ _05357_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__and3b_2
XFILLER_0_202_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13185_ _06300_ _06302_ _06339_ _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19801_ net3109 _03442_ net1848 _03441_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__o211a_1
X_12136_ _04831_ _04776_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__a21o_1
X_17993_ _01684_ _10539_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__nor2_1
X_19732_ _03294_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__clkbuf_4
X_12067_ rbzero.tex_r1\[33\] rbzero.tex_r1\[32\] _05072_ vssd1 vssd1 vccd1 vccd1 _05236_
+ sky130_fd_sc_hd__mux2_1
X_16944_ _06383_ _06344_ vssd1 vssd1 vccd1 vccd1 _09962_ sky130_fd_sc_hd__nand2_1
X_11018_ net2772 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19663_ net6172 _03360_ net2257 _03371_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__o211a_1
X_16875_ _09933_ vssd1 vssd1 vccd1 vccd1 _09934_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18614_ net3796 _02624_ _02557_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
X_15826_ _08405_ _08455_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__nor2_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19594_ net5236 _03325_ _03332_ _03330_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18545_ _02549_ _02550_ _02551_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__o21a_1
X_15757_ _08332_ _08526_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__xor2_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _06117_ _06121_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ _07825_ _07823_ _07824_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__nand3_1
XFILLER_0_158_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18476_ net7315 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__clkbuf_4
X_15688_ _08761_ _08762_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _10425_ _10426_ vssd1 vssd1 vccd1 vccd1 _10427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _07743_ _07789_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17358_ _08556_ _09251_ vssd1 vssd1 vccd1 vccd1 _10358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03996_ clknet_0__03996_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03996_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _09357_ _09382_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _10281_ _10289_ vssd1 vssd1 vccd1 vccd1 _10290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19028_ net3949 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4205 net1623 vssd1 vssd1 vccd1 vccd1 net4729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4216 net2931 vssd1 vssd1 vccd1 vccd1 net4740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4238 rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 net4762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4249 _03633_ vssd1 vssd1 vccd1 vccd1 net4773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3504 _04126_ vssd1 vssd1 vccd1 vccd1 net4028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3515 _09922_ vssd1 vssd1 vccd1 vccd1 net4039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3526 _04159_ vssd1 vssd1 vccd1 vccd1 net4050 sky130_fd_sc_hd__clkbuf_2
Xhold3537 _03967_ vssd1 vssd1 vccd1 vccd1 net4061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2803 net4474 vssd1 vssd1 vccd1 vccd1 net3327 sky130_fd_sc_hd__buf_1
Xhold3548 _05334_ vssd1 vssd1 vccd1 vccd1 net4072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 _03872_ vssd1 vssd1 vccd1 vccd1 net3338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3559 _05698_ vssd1 vssd1 vccd1 vccd1 net4083 sky130_fd_sc_hd__clkbuf_4
Xhold2825 _03820_ vssd1 vssd1 vccd1 vccd1 net3349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2836 net2892 vssd1 vssd1 vccd1 vccd1 net3360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2847 net6094 vssd1 vssd1 vccd1 vccd1 net3371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2858 rbzero.pov.spi_buffer\[70\] vssd1 vssd1 vccd1 vccd1 net3382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2869 _02392_ vssd1 vssd1 vccd1 vccd1 net3393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21823_ clknet_leaf_91_i_clk net4647 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21754_ clknet_leaf_21_i_clk net2356 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21685_ clknet_leaf_28_i_clk net5074 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20636_ _03083_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20567_ net3734 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6130 net1724 vssd1 vssd1 vccd1 vccd1 net6654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22306_ net438 net2042 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold6141 rbzero.tex_g0\[26\] vssd1 vssd1 vccd1 vccd1 net6665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6152 net1842 vssd1 vssd1 vccd1 vccd1 net6676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6163 rbzero.tex_r1\[43\] vssd1 vssd1 vccd1 vccd1 net6687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20498_ net3301 net1284 _03867_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__mux2_1
Xhold6174 net2063 vssd1 vssd1 vccd1 vccd1 net6698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6185 _04507_ vssd1 vssd1 vccd1 vccd1 net6709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5440 net2183 vssd1 vssd1 vccd1 vccd1 net5964 sky130_fd_sc_hd__dlygate4sd3_1
X_22237_ net369 net1517 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold5451 rbzero.tex_r1\[12\] vssd1 vssd1 vccd1 vccd1 net5975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6196 net1871 vssd1 vssd1 vccd1 vccd1 net6720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5462 _04419_ vssd1 vssd1 vccd1 vccd1 net5986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5473 _00687_ vssd1 vssd1 vccd1 vccd1 net5997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5484 net3732 vssd1 vssd1 vccd1 vccd1 net6008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5495 rbzero.pov.ready_buffer\[10\] vssd1 vssd1 vccd1 vccd1 net6019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4750 rbzero.spi_registers.texadd1\[19\] vssd1 vssd1 vccd1 vccd1 net5274 sky130_fd_sc_hd__dlygate4sd3_1
X_22168_ net300 net1796 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold4761 net866 vssd1 vssd1 vccd1 vccd1 net5285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4772 _00728_ vssd1 vssd1 vccd1 vccd1 net5296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4783 _00731_ vssd1 vssd1 vccd1 vccd1 net5307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4794 net939 vssd1 vssd1 vccd1 vccd1 net5318 sky130_fd_sc_hd__dlygate4sd3_1
X_21119_ _04018_ _04106_ _04107_ _03083_ net4653 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a32o_1
X_22099_ net231 net2039 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
X_14990_ _08131_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13941_ _06844_ _07090_ _06881_ _06923_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__nand4_2
X_16660_ _09729_ _09730_ vssd1 vssd1 vccd1 vccd1 _09731_ sky130_fd_sc_hd__xnor2_1
X_13872_ _06985_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15611_ _08683_ _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12823_ _05980_ _05981_ net25 vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16591_ _09305_ _09418_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18330_ net4511 net4374 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__nand2_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15542_ _08166_ _08167_ _08614_ _08616_ _08296_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__a311o_1
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ net43 _05895_ _05903_ net46 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a22o_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _02208_ _02211_ _02209_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__o21a_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11705_ _04831_ net2925 vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
X_15473_ _08299_ _08546_ _08547_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__a21o_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _05842_ _05845_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nand2_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17212_ _10198_ _10199_ vssd1 vssd1 vccd1 vccd1 _10213_ sky130_fd_sc_hd__or2_1
X_14424_ _07474_ _07509_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__nor2_1
X_11636_ net4033 net4013 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__or2_1
X_18192_ _02148_ _02115_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17143_ _10137_ _10138_ _10143_ vssd1 vssd1 vccd1 vccd1 _10145_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14355_ _07485_ _07505_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__or2_1
X_11567_ _04718_ _04733_ _04738_ _04727_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__03781_ clknet_0__03781_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03781_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13306_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__nor2_1
X_17074_ net4595 net4362 vssd1 vssd1 vccd1 vccd1 _10077_ sky130_fd_sc_hd__nor2_1
X_14286_ _07406_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__xnor2_4
Xhold709 net5252 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ rbzero.texu_hot\[4\] _04651_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16025_ _09095_ _09098_ _09093_ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__a21oi_1
X_13237_ _06206_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ net3474 vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__inv_2
X_12119_ rbzero.tex_r1\[29\] rbzero.tex_r1\[28\] _05070_ vssd1 vssd1 vccd1 vccd1 _05288_
+ sky130_fd_sc_hd__mux2_1
X_17976_ _01836_ _02024_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__nand2_1
X_13099_ net4779 net3633 _06252_ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or4_1
Xhold1409 net5805 vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_19715_ net5792 _03395_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_62_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16927_ net3219 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20701__136 clknet_1_0__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__inv_2
X_19646_ net1572 _03360_ net1704 _03354_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__o211a_1
X_16858_ net4011 _09919_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__nor2_1
X_15809_ _08838_ _08870_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19577_ net1572 _03304_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ _09853_ _09858_ vssd1 vssd1 vccd1 vccd1 _09859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18528_ _02545_ _08195_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18459_ _06269_ net3060 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21470_ clknet_leaf_0_i_clk net3023 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20421_ net3250 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20782__208 clknet_1_0__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__inv_2
XFILLER_0_109_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4002 net1145 vssd1 vssd1 vccd1 vccd1 net4526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold4013 net7538 vssd1 vssd1 vccd1 vccd1 net4537 sky130_fd_sc_hd__dlygate4sd3_1
X_20283_ net4881 _03675_ _03770_ _03761_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4024 net710 vssd1 vssd1 vccd1 vccd1 net4548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4035 net7550 vssd1 vssd1 vccd1 vccd1 net4559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22022_ clknet_leaf_99_i_clk net3350 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3301 net7347 vssd1 vssd1 vccd1 vccd1 net3825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4046 net3470 vssd1 vssd1 vccd1 vccd1 net4570 sky130_fd_sc_hd__buf_1
Xhold3312 _01204_ vssd1 vssd1 vccd1 vccd1 net3836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4057 net4285 vssd1 vssd1 vccd1 vccd1 net4581 sky130_fd_sc_hd__buf_2
Xhold4068 net7924 vssd1 vssd1 vccd1 vccd1 net4592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3334 _03617_ vssd1 vssd1 vccd1 vccd1 net3858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4079 net2888 vssd1 vssd1 vccd1 vccd1 net4603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2600 _03257_ vssd1 vssd1 vccd1 vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3345 _04719_ vssd1 vssd1 vccd1 vccd1 net3869 sky130_fd_sc_hd__clkbuf_2
Xhold2611 rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 net3135 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3356 net4674 vssd1 vssd1 vccd1 vccd1 net3880 sky130_fd_sc_hd__buf_2
Xhold3367 _02972_ vssd1 vssd1 vccd1 vccd1 net3891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 _03086_ vssd1 vssd1 vccd1 vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3378 _03600_ vssd1 vssd1 vccd1 vccd1 net3902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2633 _03526_ vssd1 vssd1 vccd1 vccd1 net3157 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2644 net4583 vssd1 vssd1 vccd1 vccd1 net3168 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1910 net6815 vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3389 net3211 vssd1 vssd1 vccd1 vccd1 net3913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2655 net4436 vssd1 vssd1 vccd1 vccd1 net3179 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1921 net6943 vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2666 _03794_ vssd1 vssd1 vccd1 vccd1 net3190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold69 net4262 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 _03404_ vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2677 _08213_ vssd1 vssd1 vccd1 vccd1 net3201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 net5882 vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__buf_1
Xhold2688 _02509_ vssd1 vssd1 vccd1 vccd1 net3212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 net7104 vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
X_20977__385 clknet_1_0__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__inv_2
Xhold2699 net6099 vssd1 vssd1 vccd1 vccd1 net3223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 _00892_ vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1976 _04262_ vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
X_20676__113 clknet_1_0__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__inv_2
Xhold1987 net6969 vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1998 _04449_ vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21806_ clknet_leaf_90_i_clk net2891 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21737_ clknet_leaf_23_i_clk net1885 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12470_ _05630_ _05632_ _05635_ _05010_ _05030_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21668_ clknet_leaf_14_i_clk net5134 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _04597_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_8
X_20619_ _05825_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__inv_2
X_21599_ clknet_leaf_1_i_clk net4293 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14140_ _07260_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11352_ net6874 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14071_ _07178_ _07177_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nor2_1
X_11283_ net5843 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__buf_4
Xhold5270 rbzero.spi_registers.buf_texadd2\[12\] vssd1 vssd1 vccd1 vccd1 net5794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5281 _04247_ vssd1 vssd1 vccd1 vccd1 net5805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5292 net2141 vssd1 vssd1 vccd1 vccd1 net5816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17830_ _10383_ _09420_ _01766_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__or3_1
Xhold4580 net922 vssd1 vssd1 vccd1 vccd1 net5104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4591 _01067_ vssd1 vssd1 vccd1 vccd1 net5115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17761_ _08717_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__buf_2
Xhold3890 _01001_ vssd1 vssd1 vccd1 vccd1 net4414 sky130_fd_sc_hd__dlygate4sd3_1
X_14973_ _08108_ _08109_ _08110_ _08116_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__a31o_2
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19500_ _02492_ _02495_ _03238_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nand3_4
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16712_ _09766_ _09654_ vssd1 vssd1 vccd1 vccd1 _09782_ sky130_fd_sc_hd__or2b_2
Xclkbuf_1_0__f__03999_ clknet_0__03999_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03999_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13924_ _06796_ _06896_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__nor2_1
X_17692_ _10463_ _10453_ _10568_ _01743_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19431_ net5003 _03224_ _03230_ _03220_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__o211a_1
X_16643_ _09692_ _09713_ vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13855_ _06997_ _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19362_ net1959 _03185_ net4244 _03181_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__o211a_1
X_12806_ _05950_ _05960_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a21boi_1
X_16574_ _09644_ _09645_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__or2b_1
X_10998_ net6343 net7105 _04366_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
X_13786_ _06928_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__xor2_2
X_18313_ net4499 net4435 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ net4355 rbzero.wall_tracer.visualWallDist\[-9\] _08297_ vssd1 vssd1 vccd1
+ vccd1 _08600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _05893_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__nand2_1
X_19293_ net5136 _03146_ _03152_ _03142_ vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18244_ _08540_ _09784_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__nor2_1
X_15456_ _08394_ _08444_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ _04802_ _05786_ _05796_ net4002 vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ _07548_ _07557_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__nor2_1
X_18175_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11619_ _04637_ _04614_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__and3_1
X_15387_ _08325_ _08331_ vssd1 vssd1 vccd1 vccd1 _08462_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12599_ rbzero.tex_b1\[15\] rbzero.tex_b1\[14\] _04987_ vssd1 vssd1 vccd1 vccd1 _05764_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ _09853_ _09858_ vssd1 vssd1 vccd1 vccd1 _10128_ sky130_fd_sc_hd__or2b_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14338_ _07474_ net558 vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold506 net5414 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold517 net6372 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold528 net5363 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _01432_ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _10058_ _10061_ vssd1 vssd1 vccd1 vccd1 _10062_ sky130_fd_sc_hd__nor2_1
X_14269_ _06931_ _06859_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16008_ _09054_ _09059_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__xnor2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _03385_ vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 net6767 vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _01341_ vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ _01914_ _01918_ _02006_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__and3_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 net5799 vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19629_ net5161 net799 _03351_ _03343_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21522_ clknet_leaf_28_i_clk net5070 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21453_ clknet_leaf_31_i_clk net3892 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20404_ net3662 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21384_ clknet_leaf_55_i_clk _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20266_ net3705 _03757_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__buf_1
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3120 _01176_ vssd1 vssd1 vccd1 vccd1 net3644 sky130_fd_sc_hd__dlygate4sd3_1
X_22005_ clknet_leaf_10_i_clk net5469 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
Xhold3142 _03863_ vssd1 vssd1 vccd1 vccd1 net3666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3153 _01021_ vssd1 vssd1 vccd1 vccd1 net3677 sky130_fd_sc_hd__dlygate4sd3_1
X_20197_ net5049 _03718_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2430 _00697_ vssd1 vssd1 vccd1 vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3175 rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 net3699 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2441 net7323 vssd1 vssd1 vccd1 vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3186 _03854_ vssd1 vssd1 vccd1 vccd1 net3710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2452 _00695_ vssd1 vssd1 vccd1 vccd1 net2976 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2463 _04854_ vssd1 vssd1 vccd1 vccd1 net2987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2474 _00692_ vssd1 vssd1 vccd1 vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1740 _01584_ vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 _09643_ vssd1 vssd1 vccd1 vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2496 _00614_ vssd1 vssd1 vccd1 vccd1 net3020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1751 _03369_ vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1762 net6973 vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _05125_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1773 _01138_ vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _04273_ vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ net2708 net5844 _04333_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__mux2_1
Xhold1795 net6859 vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10852_ _04243_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__clkbuf_4
X_13640_ _06790_ _06740_ _06677_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ net7203 net7191 _04255_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__mux2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _06695_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__buf_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _08383_ _08384_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _05028_ _05662_ _05670_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _06211_ _08618_ _09363_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ _08313_ _08315_ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20730__162 clknet_1_0__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__inv_2
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11404_ net7010 net6984 _04584_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__mux2_1
X_12384_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _05457_ vssd1 vssd1 vccd1 vccd1 _05551_
+ sky130_fd_sc_hd__mux2_1
X_15172_ _08264_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11335_ net6592 net6429 _04551_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14123_ _07262_ _07263_ _07273_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19980_ net721 _03578_ net4521 _03550_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18931_ _02897_ _02898_ _02900_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__and3_1
X_11266_ net6860 net7268 _04514_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__mux2_1
X_14054_ _06862_ _06864_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__nor2_1
X_13005_ _06153_ _06159_ _06107_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a21oi_1
X_18862_ _02830_ _02836_ _02824_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_203_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11197_ net5906 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17813_ _01863_ net4433 _01749_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
X_18793_ net6089 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
X_17744_ _01695_ _01764_ _01794_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a21o_1
X_14956_ _08013_ _08010_ vssd1 vssd1 vccd1 vccd1 _08101_ sky130_fd_sc_hd__or2_1
X_13907_ _07037_ _07038_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__xor2_2
X_17675_ _01671_ _01726_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ net7908 _08012_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__nor2_1
X_19414_ net647 _03212_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__or2_1
X_16626_ _08701_ _08849_ _09563_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13838_ _06957_ _06987_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__o21a_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19345_ net2113 _03173_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__or2_1
X_16557_ _09463_ _09505_ _09628_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_175_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13769_ _06915_ _06917_ _06919_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__nand3_4
XFILLER_0_128_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15508_ _08559_ _08560_ _08574_ _08582_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19276_ net5095 _03133_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16488_ _09451_ _09460_ _09458_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18227_ _02212_ _02213_ _02214_ _02215_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__o22a_1
X_15439_ net3471 _08328_ _08325_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_116_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6707 net2763 vssd1 vssd1 vccd1 vccd1 net7231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6718 rbzero.tex_r0\[55\] vssd1 vssd1 vccd1 vccd1 net7242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6729 net2866 vssd1 vssd1 vccd1 vccd1 net7253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18158_ _02128_ _02144_ _02142_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold303 net5118 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17109_ _09328_ _09312_ vssd1 vssd1 vccd1 vccd1 _10111_ sky130_fd_sc_hd__nor2_1
Xhold314 net5088 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 net5221 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18089_ _02130_ _02038_ _02136_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 net5169 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 net5179 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20120_ _03678_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold358 net5185 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 net5159 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03778_ _03778_ vssd1 vssd1 vccd1 vccd1 clknet_0__03778_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20051_ _03616_ net3243 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 net6544 vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894__309 clknet_1_0__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__inv_2
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _03420_ vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 net6044 vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1036 _03430_ vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 net6270 vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__buf_1
XFILLER_0_198_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1058 net4724 vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1069 net5742 vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20788__214 clknet_1_1__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__inv_2
X_21505_ clknet_leaf_14_i_clk net2790 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21436_ clknet_leaf_83_i_clk net4712 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_146_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21367_ clknet_leaf_53_i_clk _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11120_ net6968 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
Xhold870 net4281 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_21298_ clknet_leaf_43_i_clk _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold881 net5675 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__clkbuf_4
Xhold892 net5691 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
X_20249_ net3598 _03744_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__or2_1
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20760__188 clknet_1_0__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__inv_2
Xhold2260 net7186 vssd1 vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2271 _01114_ vssd1 vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
X_14810_ _07884_ _07916_ _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__o21ai_1
Xhold2282 _01134_ vssd1 vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _08458_ _08863_ _08864_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__nand3_1
Xhold2293 _04580_ vssd1 vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1570 net591 vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1581 _04523_ vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _07861_ _07864_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__xnor2_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1592 net6979 vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ net3016 net1603 vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_105 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_105/HI o_rgb[19]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_116 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_116/HI zeros[8] sky130_fd_sc_hd__conb_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_127 vssd1 vssd1 vccd1 vccd1 ones[3] top_ew_algofoogle_127/LO sky130_fd_sc_hd__conb_1
X_10904_ net2335 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__clkbuf_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ net4501 net4417 vssd1 vssd1 vccd1 vccd1 _10459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_138 vssd1 vssd1 vccd1 vccd1 ones[14] top_ew_algofoogle_138/LO sky130_fd_sc_hd__conb_1
XFILLER_0_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _07618_ _07354_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_212_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _05037_ vssd1 vssd1 vccd1 vccd1 _05054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16411_ _09483_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13623_ _06697_ _06698_ _06627_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17391_ _10388_ _10389_ vssd1 vssd1 vccd1 vccd1 _10391_ sky130_fd_sc_hd__or2_1
X_10835_ net6634 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ net5155 _03053_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__or2_1
X_16342_ _09389_ _09391_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__or2_1
X_13554_ _06703_ _06704_ _06692_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__mux2_1
X_10766_ net7243 net6395 _04244_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _05219_ vssd1 vssd1 vccd1 vccd1 _05671_
+ sky130_fd_sc_hd__mux2_1
X_19061_ net3088 net2843 _03014_ _03011_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16273_ _09345_ _09346_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__nand2_1
X_10697_ net6644 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__clkbuf_1
X_13485_ _06531_ _06635_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18012_ _01986_ _02060_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__xnor2_2
X_15224_ _08298_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__clkbuf_8
X_12436_ _05568_ _05602_ _04975_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__mux2_2
XFILLER_0_125_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _08255_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
X_12367_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _05218_ vssd1 vssd1 vccd1 vccd1 _05534_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14106_ _07071_ _07256_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11318_ net7135 net7123 _04540_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__mux2_1
X_12298_ _04993_ _05465_ _04999_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__o21a_1
X_19963_ net3483 _03471_ _03568_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a22o_1
X_15086_ _08190_ _08207_ net3357 _01622_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ net6696 net6758 _04503_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__mux2_1
X_14037_ net528 _07185_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__nand2_1
X_18914_ _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19894_ _03483_ _03520_ _03474_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_207_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18845_ net4709 _02823_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18776_ net3807 net2884 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15988_ _09055_ _09056_ _09057_ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__o21a_1
XFILLER_0_207_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17727_ _08630_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14939_ _08080_ _08085_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__nand2_2
XFILLER_0_171_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17658_ _10302_ _10544_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_212_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ _09673_ _09679_ vssd1 vssd1 vccd1 vccd1 _09680_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20737__168 clknet_1_1__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__inv_2
XFILLER_0_212_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17589_ _10130_ _09420_ _09538_ _09562_ vssd1 vssd1 vccd1 vccd1 _10587_ sky130_fd_sc_hd__o22a_1
XFILLER_0_175_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19328_ _03035_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7216 net4312 vssd1 vssd1 vccd1 vccd1 net7740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19259_ _03039_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__clkbuf_4
Xhold7227 net4576 vssd1 vssd1 vccd1 vccd1 net7751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7238 rbzero.wall_tracer.stepDistX\[-11\] vssd1 vssd1 vccd1 vccd1 net7762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6504 net2237 vssd1 vssd1 vccd1 vccd1 net7028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7249 _08451_ vssd1 vssd1 vccd1 vccd1 net7773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6515 _04536_ vssd1 vssd1 vccd1 vccd1 net7039 sky130_fd_sc_hd__dlygate4sd3_1
X_22270_ net402 net2710 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
Xhold6526 net2271 vssd1 vssd1 vccd1 vccd1 net7050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6537 _04252_ vssd1 vssd1 vccd1 vccd1 net7061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5803 rbzero.spi_registers.mosi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6548 rbzero.tex_r1\[8\] vssd1 vssd1 vccd1 vccd1 net7072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5814 _04521_ vssd1 vssd1 vccd1 vccd1 net6338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6559 net2128 vssd1 vssd1 vccd1 vccd1 net7083 sky130_fd_sc_hd__dlygate4sd3_1
X_21221_ clknet_leaf_43_i_clk net1065 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold100 net6321 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5825 net1127 vssd1 vssd1 vccd1 vccd1 net6349 sky130_fd_sc_hd__buf_1
Xhold5836 _04219_ vssd1 vssd1 vccd1 vccd1 net6360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _01362_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5847 net1040 vssd1 vssd1 vccd1 vccd1 net6371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 net4153 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5858 rbzero.tex_g0\[52\] vssd1 vssd1 vccd1 vccd1 net6382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold133 net4174 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 rbzero.pov.ready_buffer\[55\] vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5869 net1074 vssd1 vssd1 vccd1 vccd1 net6393 sky130_fd_sc_hd__dlygate4sd3_1
X_21152_ _04626_ _04818_ net4910 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o21ai_1
Xhold155 net4177 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 net4967 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 net7613 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 net4396 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ _03664_ _03661_ net3329 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__and3b_1
Xhold199 net7615 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkdlybuf4s25_1
X_21083_ _04070_ _04074_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20034_ _03616_ net3544 vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__or2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ net210 net1755 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ net5824 net2427 _04170_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270_ rbzero.wall_tracer.rayAddendX\[-3\] _06420_ _06414_ vssd1 vssd1 vccd1 vccd1
+ _06421_ sky130_fd_sc_hd__mux2_4
X_22468_ clknet_leaf_80_i_clk net4660 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ _04881_ _04806_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__or3_1
X_21419_ clknet_leaf_85_i_clk net4699 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_22399_ net151 net2381 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
X_12152_ net4092 _04906_ _05320_ net4065 vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ net2361 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12083_ _05248_ _05249_ _05251_ _05009_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__o211a_1
X_16960_ net2611 net2807 _09968_ vssd1 vssd1 vccd1 vccd1 _09976_ sky130_fd_sc_hd__o21a_1
X_20842__263 clknet_1_0__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__inv_2
X_11034_ net7099 net6684 _04392_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
X_15911_ _08983_ _08985_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__xnor2_1
X_16891_ net4109 _09937_ _09938_ _08155_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18630_ net3796 rbzero.wall_tracer.rayAddendX\[1\] net4666 vssd1 vssd1 vccd1 vccd1
+ _02640_ sky130_fd_sc_hd__o21a_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _08372_ _08663_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__nor2_2
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2090 _04537_ vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _02571_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _08811_ _08847_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__xnor2_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ _06129_ _06126_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__nand2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _10509_ _10510_ vssd1 vssd1 vccd1 vccd1 _10511_ sky130_fd_sc_hd__xnor2_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _07851_ _07873_ _07874_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__a21oi_1
X_11936_ net4239 _05000_ _04984_ _05037_ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a41o_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ net3904 _02503_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _10316_ _10318_ vssd1 vssd1 vccd1 vccd1 _10443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14655_ _07471_ _07805_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__nor2_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11867_ _05014_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _06666_ _06628_ _06686_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__or3_1
X_17374_ _10372_ _10373_ vssd1 vssd1 vccd1 vccd1 _10374_ sky130_fd_sc_hd__nand2_1
X_10818_ net2669 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14586_ _07715_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__xor2_4
X_11798_ _04914_ _04917_ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19113_ net5406 _03040_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__or2_1
X_16325_ _09265_ _09266_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ _06687_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__clkbuf_4
X_10749_ net2368 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ net3112 _02988_ _03004_ _02993_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__o211a_1
X_16256_ _09327_ _09329_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__nand2_1
X_13468_ _06617_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_211_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15207_ _08284_ net1068 net3622 vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__mux2_1
X_12419_ rbzero.tex_g1\[27\] rbzero.tex_g1\[26\] _05456_ vssd1 vssd1 vccd1 vccd1 _05586_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16187_ _08742_ _09248_ _09261_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__a21oi_4
X_13399_ _06433_ _06535_ _06527_ _06537_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4409 _08248_ vssd1 vssd1 vccd1 vccd1 net4933 sky130_fd_sc_hd__clkbuf_2
X_15138_ net4828 _06386_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3719 net4235 vssd1 vssd1 vccd1 vccd1 net4243 sky130_fd_sc_hd__dlygate4sd3_1
X_15069_ net4507 net4467 _08191_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__mux2_1
X_19946_ net4387 net4675 _03553_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__or3_1
X_19877_ net3995 _03503_ _03484_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o21ai_1
X_18828_ net4708 rbzero.wall_tracer.rayAddendY\[1\] vssd1 vssd1 vccd1 vccd1 _02818_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18759_ net4439 net4621 _02752_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21770_ clknet_leaf_4_i_clk net2157 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7002 rbzero.wall_tracer.trackDistY\[3\] vssd1 vssd1 vccd1 vccd1 net7526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7013 rbzero.traced_texa\[9\] vssd1 vssd1 vccd1 vccd1 net7537 sky130_fd_sc_hd__dlygate4sd3_1
X_20583_ net3516 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7024 rbzero.wall_tracer.trackDistX\[-8\] vssd1 vssd1 vccd1 vccd1 net7548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6301 _04305_ vssd1 vssd1 vccd1 vccd1 net6825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6312 net1821 vssd1 vssd1 vccd1 vccd1 net6836 sky130_fd_sc_hd__dlygate4sd3_1
X_22322_ net454 net2447 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7057 _02891_ vssd1 vssd1 vccd1 vccd1 net7581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6323 rbzero.tex_r1\[41\] vssd1 vssd1 vccd1 vccd1 net6847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6334 net2241 vssd1 vssd1 vccd1 vccd1 net6858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6345 _04231_ vssd1 vssd1 vccd1 vccd1 net6869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22253_ net385 net1208 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold6356 net1683 vssd1 vssd1 vccd1 vccd1 net6880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5611 _08241_ vssd1 vssd1 vccd1 vccd1 net6135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5622 net3772 vssd1 vssd1 vccd1 vccd1 net6146 sky130_fd_sc_hd__clkbuf_4
Xhold6367 rbzero.tex_g0\[14\] vssd1 vssd1 vccd1 vccd1 net6891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6378 net1835 vssd1 vssd1 vccd1 vccd1 net6902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5633 net746 vssd1 vssd1 vccd1 vccd1 net6157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6389 rbzero.tex_g0\[30\] vssd1 vssd1 vccd1 vccd1 net6913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21204_ net660 net6555 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__xnor2_1
Xhold5644 net2982 vssd1 vssd1 vccd1 vccd1 net6168 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4910 rbzero.spi_registers.texadd3\[3\] vssd1 vssd1 vccd1 vccd1 net5434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5655 rbzero.spi_registers.buf_texadd1\[8\] vssd1 vssd1 vccd1 vccd1 net6179 sky130_fd_sc_hd__dlygate4sd3_1
X_22184_ net316 net1676 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4921 _01085_ vssd1 vssd1 vccd1 vccd1 net5445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5666 rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 net6190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4932 _01595_ vssd1 vssd1 vccd1 vccd1 net5456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5677 rbzero.spi_registers.buf_texadd2\[8\] vssd1 vssd1 vccd1 vccd1 net6201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4943 net1070 vssd1 vssd1 vccd1 vccd1 net5467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5688 rbzero.debug_overlay.playerY\[3\] vssd1 vssd1 vccd1 vccd1 net6212 sky130_fd_sc_hd__dlygate4sd3_1
X_21135_ _04115_ _04118_ _04119_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__o211ai_2
Xhold5699 _02776_ vssd1 vssd1 vccd1 vccd1 net6223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4954 _00733_ vssd1 vssd1 vccd1 vccd1 net5478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4965 net1097 vssd1 vssd1 vccd1 vccd1 net5489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4976 net1105 vssd1 vssd1 vccd1 vccd1 net5500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4987 _00390_ vssd1 vssd1 vccd1 vccd1 net5511 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__05840_ clknet_0__05840_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05840_
+ sky130_fd_sc_hd__clkbuf_16
Xhold4998 rbzero.spi_registers.texadd2\[20\] vssd1 vssd1 vccd1 vccd1 net5522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21066_ _04018_ _04061_ _04062_ _04017_ net4395 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a32o_1
X_20017_ rbzero.debug_overlay.facingY\[-3\] _03582_ vssd1 vssd1 vccd1 vccd1 _03610_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_154_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ net20 _05926_ _05929_ _05920_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21968_ net193 net2432 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _04831_ _04886_ _04888_ net2726 _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__o221a_1
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20872__289 clknet_1_1__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__inv_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ clknet_leaf_95_i_clk net5051 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _07356_ _07590_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ net3893 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ net4052 vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__buf_2
X_14371_ _07302_ _07305_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _04724_ _04669_ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16110_ _08730_ _08740_ _08738_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13322_ net4406 net4787 vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__or2_1
X_17090_ _10090_ _10091_ vssd1 vssd1 vccd1 vccd1 _10092_ sky130_fd_sc_hd__nor2_2
XFILLER_0_122_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16041_ _09075_ _09072_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13253_ net5491 _06396_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__xnor2_1
X_20340__73 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_0_161_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _05341_ _05365_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__and2b_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13184_ _06304_ _06306_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20766__194 clknet_1_1__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__inv_2
XFILLER_0_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19800_ net6722 _03443_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__or2_1
X_12135_ net4033 _04759_ _04606_ net4014 vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a22o_1
X_17992_ _10520_ _10416_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19731_ net2094 _03408_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__or2_1
X_16943_ _09946_ net4876 vssd1 vssd1 vccd1 vccd1 _09961_ sky130_fd_sc_hd__nand2_1
X_12066_ _05002_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__buf_4
XFILLER_0_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ net52 net2771 _04310_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
X_16874_ _09932_ vssd1 vssd1 vccd1 vccd1 _09933_ sky130_fd_sc_hd__clkbuf_8
X_19662_ net6180 _03362_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__or2_1
X_15825_ _08899_ _08490_ _08491_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__and3_1
X_18613_ _02618_ _02623_ _04632_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ net3933 _03327_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__or2_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _08806_ _08830_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__xor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ net4446 _02548_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _06122_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14707_ _07849_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _04987_ vssd1 vssd1 vccd1 vccd1 _05089_
+ sky130_fd_sc_hd__mux2_1
X_18475_ net3925 net3960 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15687_ _08564_ _08560_ _08565_ _08559_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__o22ai_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _06052_ _06046_ net6347 vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _10422_ _10423_ _10424_ vssd1 vssd1 vccd1 vccd1 _10426_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14638_ _07763_ _07787_ _07788_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _08556_ _08795_ vssd1 vssd1 vccd1 vccd1 _10357_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14569_ _07672_ _07677_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03995_ clknet_0__03995_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03995_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _09379_ _09381_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__xor2_2
X_17288_ _10283_ _10288_ vssd1 vssd1 vccd1 vccd1 _10289_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20849__269 clknet_1_1__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__inv_2
XFILLER_0_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19027_ net1572 _02988_ net1468 _02993_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__o211a_1
X_16239_ _08325_ _09312_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4206 _01019_ vssd1 vssd1 vccd1 vccd1 net4730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4217 _01608_ vssd1 vssd1 vccd1 vccd1 net4741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4228 _02638_ vssd1 vssd1 vccd1 vccd1 net4752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4239 net979 vssd1 vssd1 vccd1 vccd1 net4763 sky130_fd_sc_hd__buf_1
Xhold3505 _04129_ vssd1 vssd1 vccd1 vccd1 net4029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3516 _00478_ vssd1 vssd1 vccd1 vccd1 net4040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3527 gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 net4051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3538 _01260_ vssd1 vssd1 vccd1 vccd1 net4062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2804 net7324 vssd1 vssd1 vccd1 vccd1 net3328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3549 _05352_ vssd1 vssd1 vccd1 vccd1 net4073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 _03873_ vssd1 vssd1 vccd1 vccd1 net3339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2826 _01191_ vssd1 vssd1 vccd1 vccd1 net3350 sky130_fd_sc_hd__dlygate4sd3_1
X_19929_ net6191 _03530_ net2957 _03496_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__o211a_1
Xhold2837 _03900_ vssd1 vssd1 vccd1 vccd1 net3361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2848 _00586_ vssd1 vssd1 vccd1 vccd1 net3372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2859 net1220 vssd1 vssd1 vccd1 vccd1 net3383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21822_ clknet_leaf_91_i_clk net3142 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21753_ clknet_leaf_21_i_clk net1576 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21684_ clknet_leaf_28_i_clk net5089 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20635_ _04802_ net4061 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20566_ _03902_ net3733 vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6120 net1748 vssd1 vssd1 vccd1 vccd1 net6644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6131 rbzero.tex_g0\[9\] vssd1 vssd1 vccd1 vccd1 net6655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22305_ net437 net2012 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold6142 net1944 vssd1 vssd1 vccd1 vccd1 net6666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20908__322 clknet_1_1__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__inv_2
Xhold6153 rbzero.tex_g0\[41\] vssd1 vssd1 vccd1 vccd1 net6677 sky130_fd_sc_hd__dlygate4sd3_1
X_20497_ net3307 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6164 net1853 vssd1 vssd1 vccd1 vccd1 net6688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5430 _04533_ vssd1 vssd1 vccd1 vccd1 net5954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6175 _04301_ vssd1 vssd1 vccd1 vccd1 net6699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5441 rbzero.map_overlay.i_mapdx\[0\] vssd1 vssd1 vccd1 vccd1 net5965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6186 net1839 vssd1 vssd1 vccd1 vccd1 net6710 sky130_fd_sc_hd__dlygate4sd3_1
X_22236_ net368 net2878 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold5452 net5927 vssd1 vssd1 vccd1 vccd1 net5976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6197 rbzero.spi_registers.buf_texadd3\[18\] vssd1 vssd1 vccd1 vccd1 net6721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5463 net1939 vssd1 vssd1 vccd1 vccd1 net5987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5474 rbzero.map_overlay.i_mapdx\[1\] vssd1 vssd1 vccd1 vccd1 net5998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5485 _03492_ vssd1 vssd1 vccd1 vccd1 net6009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4740 _00778_ vssd1 vssd1 vccd1 vccd1 net5264 sky130_fd_sc_hd__dlygate4sd3_1
X_22167_ net299 net2618 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold5496 net2900 vssd1 vssd1 vccd1 vccd1 net6020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4751 net943 vssd1 vssd1 vccd1 vccd1 net5275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4762 rbzero.spi_registers.texadd3\[19\] vssd1 vssd1 vccd1 vccd1 net5286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4773 rbzero.spi_registers.texadd1\[0\] vssd1 vssd1 vccd1 vccd1 net5297 sky130_fd_sc_hd__dlygate4sd3_1
X_21118_ _04104_ _04105_ _04103_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o21ai_1
Xhold4784 net1039 vssd1 vssd1 vccd1 vccd1 net5308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4795 _00858_ vssd1 vssd1 vccd1 vccd1 net5319 sky130_fd_sc_hd__dlygate4sd3_1
X_22098_ net230 net1482 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13940_ _06844_ _07090_ _06881_ _06923_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__a22o_1
X_21049_ _04043_ _04044_ _04045_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _07010_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_202_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15610_ _08411_ _08684_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__nor2_1
X_12822_ _04159_ net4891 _04726_ _04777_ net22 net23 vssd1 vssd1 vccd1 vccd1 _05981_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_202_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16590_ _09419_ _09540_ _09133_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__or3b_1
X_20954__364 clknet_1_0__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__inv_2
XFILLER_0_55_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _08152_ _08155_ _08160_ _08575_ _08615_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__o41a_1
XFILLER_0_16_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12753_ net44 _05905_ _05894_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18260_ _02302_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__xnor2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _04831_ net2925 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__or2_1
X_15472_ net3161 _08298_ _06209_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__o21ai_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12684_ _05843_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__and2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _10209_ _10210_ _10084_ net7824 vssd1 vssd1 vccd1 vccd1 _10212_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _07467_ _07493_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18191_ _02236_ _02237_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__xor2_1
X_11635_ net4032 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _10137_ _10138_ _10143_ vssd1 vssd1 vccd1 vccd1 _10144_ sky130_fd_sc_hd__a21oi_1
X_14354_ _07478_ _07484_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__03780_ clknet_0__03780_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03780_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11566_ _04724_ _04734_ _04735_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a31o_1
X_13305_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17073_ net4595 net4362 vssd1 vssd1 vccd1 vccd1 _10076_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14285_ _07407_ _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_40_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _04656_ _04666_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a21o_1
X_16024_ _09093_ _09095_ _09098_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__nand3_1
X_13236_ _06204_ _06211_ _06388_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__a211o_2
XFILLER_0_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _06312_ net3795 _06321_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ rbzero.tex_r1\[31\] rbzero.tex_r1\[30\] _05262_ vssd1 vssd1 vccd1 vccd1 _05287_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17975_ _02020_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__xnor2_1
X_13098_ net656 net695 net692 _06253_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__or4_1
X_19714_ net1727 _03393_ net1884 _03400_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__o211a_1
X_12049_ _05070_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__clkbuf_8
X_16926_ _04692_ net3218 _09943_ vssd1 vssd1 vccd1 vccd1 _09945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19645_ net6300 _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or2_1
X_16857_ net3762 _09919_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__nor2_1
X_15808_ _08879_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__xnor2_2
X_16788_ _09854_ _09857_ vssd1 vssd1 vccd1 vccd1 _09858_ sky130_fd_sc_hd__xnor2_1
X_19576_ net5283 _03302_ _03320_ _03314_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15739_ net3722 _08379_ _08546_ _08547_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__or4_2
X_18527_ net4424 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18458_ _02476_ _02478_ net3059 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _10406_ _09861_ _10407_ _09108_ vssd1 vssd1 vccd1 vccd1 _10409_ sky130_fd_sc_hd__o22ai_1
X_18389_ _02419_ _02420_ _02414_ net3235 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20420_ net3325 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20304__40 clknet_1_1__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4003 net7548 vssd1 vssd1 vccd1 vccd1 net4527 sky130_fd_sc_hd__dlygate4sd3_1
X_20282_ net3383 _03678_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__or2_1
Xhold4014 net3233 vssd1 vssd1 vccd1 vccd1 net4538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4025 rbzero.debug_overlay.vplaneY\[-5\] vssd1 vssd1 vccd1 vccd1 net4549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4036 net3500 vssd1 vssd1 vccd1 vccd1 net4560 sky130_fd_sc_hd__buf_1
X_22021_ clknet_leaf_99_i_clk net3456 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3302 _03668_ vssd1 vssd1 vccd1 vccd1 net3826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4047 _08252_ vssd1 vssd1 vccd1 vccd1 net4571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3313 rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 net3837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4058 _08228_ vssd1 vssd1 vccd1 vccd1 net4582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4069 net3537 vssd1 vssd1 vccd1 vccd1 net4593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3324 net7345 vssd1 vssd1 vccd1 vccd1 net3848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3335 _03618_ vssd1 vssd1 vccd1 vccd1 net3859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2601 _03258_ vssd1 vssd1 vccd1 vccd1 net3125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3346 _04720_ vssd1 vssd1 vccd1 vccd1 net3870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2612 net7321 vssd1 vssd1 vccd1 vccd1 net3136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3357 _06232_ vssd1 vssd1 vccd1 vccd1 net3881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3368 _00622_ vssd1 vssd1 vccd1 vccd1 net3892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2623 _00688_ vssd1 vssd1 vccd1 vccd1 net3147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3379 _00996_ vssd1 vssd1 vccd1 vccd1 net3903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 _03527_ vssd1 vssd1 vccd1 vccd1 net3158 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1900 net7112 vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2645 net7744 vssd1 vssd1 vccd1 vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1911 _01318_ vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2656 net3956 vssd1 vssd1 vccd1 vccd1 net3180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1922 net6945 vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2667 _03795_ vssd1 vssd1 vccd1 vccd1 net3191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1933 _00908_ vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2678 _00421_ vssd1 vssd1 vccd1 vccd1 net3202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1944 net5884 vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2689 _02522_ vssd1 vssd1 vccd1 vccd1 net3213 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold1955 _04376_ vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1966 net7182 vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1977 _01506_ vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1988 _04578_ vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1999 _01338_ vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21805_ clknet_leaf_89_i_clk net4296 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21736_ clknet_leaf_23_i_clk net2115 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21667_ clknet_leaf_27_i_clk net3867 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11420_ _04241_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20618_ net3965 net4018 net3966 _08276_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21598_ clknet_leaf_1_i_clk net4263 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11351_ net6872 net2619 _04551_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20549_ net3249 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__clkbuf_4
X_14070_ _07218_ _07220_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__nor2_1
X_11282_ net2037 net5841 _04169_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5260 _03272_ vssd1 vssd1 vccd1 vccd1 net5784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _06133_ _06176_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__or2_2
X_22219_ net351 net2441 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold5271 net1655 vssd1 vssd1 vccd1 vccd1 net5795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5282 net1933 vssd1 vssd1 vccd1 vccd1 net5806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5293 rbzero.tex_b0\[58\] vssd1 vssd1 vccd1 vccd1 net5817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4570 rbzero.spi_registers.buf_texadd0\[22\] vssd1 vssd1 vccd1 vccd1 net5094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4581 rbzero.spi_registers.texadd3\[20\] vssd1 vssd1 vccd1 vccd1 net5105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4592 rbzero.color_sky\[1\] vssd1 vssd1 vccd1 vccd1 net5116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3880 net7839 vssd1 vssd1 vccd1 vccd1 net4404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17760_ _01809_ _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__xnor2_1
Xhold3891 net1099 vssd1 vssd1 vccd1 vccd1 net4415 sky130_fd_sc_hd__dlygate4sd3_1
X_14972_ _08068_ _08115_ net6162 vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16711_ _09652_ _09779_ _09780_ vssd1 vssd1 vccd1 vccd1 _09781_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_1_0__f__03998_ clknet_0__03998_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03998_
+ sky130_fd_sc_hd__clkbuf_16
X_13923_ _06865_ net564 vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__nor2_1
X_17691_ _10462_ _01742_ _10567_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20878__295 clknet_1_0__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__inv_2
XFILLER_0_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16642_ _09711_ _09712_ vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__and2_1
X_19430_ net1844 _03225_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ _07003_ _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12805_ net25 _05961_ _05963_ net24 vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a31o_1
X_16573_ _09642_ net3009 vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__or2_1
X_19361_ net4243 _03186_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _06930_ _06935_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__xnor2_2
X_10997_ net7024 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15524_ _08596_ _08597_ _08598_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__a21o_1
X_18312_ net4499 net4435 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__nor2_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _05894_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and2_1
X_19292_ net1604 _03147_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18243_ _02228_ _02229_ _02288_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__o21a_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _08353_ _08405_ _08424_ _08529_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ net5957 vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14406_ _07550_ _07556_ _07554_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18174_ _08793_ _09375_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _04759_ _04776_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__or2_2
X_15386_ _08397_ _08446_ _08460_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__a21o_1
X_12598_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _05014_ vssd1 vssd1 vccd1 vccd1 _05763_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17125_ _09838_ _09845_ _10126_ vssd1 vssd1 vccd1 vccd1 _10127_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ _07361_ _07403_ _07487_ _07486_ _07443_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__a32o_1
XFILLER_0_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11549_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 net6350 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _01572_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _10059_ net3398 vssd1 vssd1 vccd1 vccd1 _10061_ sky130_fd_sc_hd__or2b_1
Xhold529 net5365 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ _06867_ _06880_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16007_ _09080_ _09081_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ rbzero.map_rom.f4 net4896 _06186_ _06216_ vssd1 vssd1 vccd1 vccd1 _06375_
+ sky130_fd_sc_hd__a22o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _07348_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__xor2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _00895_ vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _04372_ vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
X_17958_ _01914_ _01918_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a21oi_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1229 net6723 vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16909_ net4173 _09939_ _09940_ net6281 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__a22o_1
X_17889_ _09108_ _10406_ _01711_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_178_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19628_ net642 _03340_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19559_ net5099 _03303_ _03311_ _03295_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21521_ clknet_leaf_34_i_clk net2967 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21452_ clknet_leaf_31_i_clk net3750 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20403_ _03791_ net3661 vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21383_ clknet_leaf_56_i_clk _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20265_ net3705 _03756_ net4851 _03761_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3110 net6135 vssd1 vssd1 vccd1 vccd1 net3634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3121 net5778 vssd1 vssd1 vccd1 vccd1 net3645 sky130_fd_sc_hd__dlygate4sd3_1
X_22004_ net229 net2036 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3132 net7333 vssd1 vssd1 vccd1 vccd1 net3656 sky130_fd_sc_hd__dlygate4sd3_1
X_20196_ net5049 _03717_ _03721_ _03722_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__o211a_1
Xhold3143 _03864_ vssd1 vssd1 vccd1 vccd1 net3667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3154 net4856 vssd1 vssd1 vccd1 vccd1 net3678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3165 _02685_ vssd1 vssd1 vccd1 vccd1 net3689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2420 rbzero.pov.ready_buffer\[64\] vssd1 vssd1 vccd1 vccd1 net2944 sky130_fd_sc_hd__buf_1
XFILLER_0_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3176 _02790_ vssd1 vssd1 vccd1 vccd1 net3700 sky130_fd_sc_hd__buf_2
Xhold2431 net4610 vssd1 vssd1 vccd1 vccd1 net2955 sky130_fd_sc_hd__buf_2
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2442 _03090_ vssd1 vssd1 vccd1 vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3187 _03855_ vssd1 vssd1 vccd1 vccd1 net3711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3198 net6133 vssd1 vssd1 vccd1 vccd1 net3722 sky130_fd_sc_hd__clkbuf_4
Xhold2453 rbzero.spi_registers.sclk_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net2977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 _03951_ vssd1 vssd1 vccd1 vccd1 net2988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 _04331_ vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2475 rbzero.pov.ready_buffer\[66\] vssd1 vssd1 vccd1 vccd1 net2999 sky130_fd_sc_hd__buf_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1741 net7094 vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2486 rbzero.spi_registers.buf_texadd1\[10\] vssd1 vssd1 vccd1 vccd1 net3010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1752 _00883_ vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2497 net6234 vssd1 vssd1 vccd1 vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1763 _01315_ vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 net7043 vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
X_10920_ net5933 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__clkbuf_1
Xhold1785 _01496_ vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1796 _04518_ vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10851_ net1974 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _06707_ _06688_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__xnor2_2
X_10782_ net2500 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12521_ _05023_ _05674_ _05678_ _05686_ _05051_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__o311a_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21719_ clknet_leaf_8_i_clk net1649 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ net7552 _08314_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__nand2_2
XFILLER_0_137_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _05111_ net3014 net3378 vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11403_ net6600 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__buf_1
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15171_ net4349 _08155_ _08260_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__mux2_1
X_12383_ _04978_ _05536_ _05540_ _05545_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__o32a_1
X_14122_ _07266_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__xnor2_1
X_11334_ net2391 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14053_ _07202_ _07203_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__nand2_1
X_18930_ _02893_ net3700 _02894_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__and3_1
X_11265_ net7189 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_76_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold5090 net1377 vssd1 vssd1 vccd1 vccd1 net5614 sky130_fd_sc_hd__dlygate4sd3_1
X_13004_ _06153_ _06159_ _06107_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__and3_1
X_18861_ _02847_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11196_ net5868 net5904 _04470_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17812_ _06206_ _01755_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__o21ai_1
X_18792_ rbzero.wall_tracer.rayAddendY\[-3\] _02785_ _02714_ vssd1 vssd1 vccd1 vccd1
+ _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17743_ _01776_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__xnor2_2
X_14955_ net7891 _08098_ _08099_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13906_ _07044_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__xnor2_2
X_17674_ _01724_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__xor2_1
X_14886_ net7434 _08009_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__nor2_1
X_19413_ net5102 _03211_ _03219_ _03220_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16625_ _08317_ _09695_ _09562_ _08331_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__o22a_1
X_13837_ _06668_ _06957_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16556_ _09502_ _09504_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19344_ net5652 _03172_ _03180_ _03181_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__o211a_1
X_13768_ _06736_ _06918_ _06861_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__o21ai_2
X_15507_ _08581_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__clkbuf_4
X_12719_ _05871_ _05879_ net12 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__mux2_1
X_16487_ _09533_ _09558_ vssd1 vssd1 vccd1 vccd1 _09559_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19275_ net5076 _03132_ _03140_ _03142_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13699_ _06733_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15438_ _08502_ _08505_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__xnor2_1
X_18226_ _02080_ _02248_ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_29_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6708 rbzero.tex_r0\[48\] vssd1 vssd1 vccd1 vccd1 net7232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6719 net2418 vssd1 vssd1 vccd1 vccd1 net7243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18157_ _02202_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _08312_ _08438_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__o21ai_4
X_17108_ _09813_ _10109_ vssd1 vssd1 vccd1 vccd1 _10110_ sky130_fd_sc_hd__xor2_1
Xhold304 net6342 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold315 rbzero.traced_texa\[-10\] vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _02134_ _02135_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 net5223 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 net5139 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold348 net5333 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _10041_ _10044_ _10019_ vssd1 vssd1 vccd1 vccd1 _10046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03777_ _03777_ vssd1 vssd1 vccd1 vccd1 clknet_0__03777_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold359 net5187 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20050_ net3242 net3229 _03580_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _01387_ vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 net4329 vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1026 net6045 vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 _00925_ vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 _02986_ vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__buf_4
Xhold1059 net4468 vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__buf_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20714__147 clknet_1_1__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__inv_2
X_21504_ clknet_leaf_14_i_clk net2880 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21435_ clknet_leaf_82_i_clk net3727 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21366_ clknet_leaf_53_i_clk _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 _04499_ vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
X_21297_ clknet_leaf_41_i_clk _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[0\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold871 net3434 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 net1783 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 net6476 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _04242_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__buf_4
X_20248_ net3598 _03743_ _03751_ _03748_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__o211a_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20179_ net3843 _03704_ _03712_ _03709_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__o211a_1
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 net5965 vssd1 vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2261 net7188 vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2272 net7250 vssd1 vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2283 net7653 vssd1 vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__clkbuf_2
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 _01125_ vssd1 vssd1 vccd1 vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1560 _01563_ vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _07889_ _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__xnor2_1
Xhold1571 _03412_ vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ net1673 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__inv_2
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1582 _01270_ vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 _04446_ vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_106 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_106/HI o_rgb[20]
+ sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_117 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_117/HI zeros[9] sky130_fd_sc_hd__conb_1
X_10903_ net5989 net6904 _04321_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__mux2_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_128 vssd1 vssd1 vccd1 vccd1 ones[4] top_ew_algofoogle_128/LO sky130_fd_sc_hd__conb_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _07776_ _07775_ _07773_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__a21o_1
Xtop_ew_algofoogle_139 vssd1 vssd1 vccd1 vccd1 ones[15] top_ew_algofoogle_139/LO sky130_fd_sc_hd__conb_1
XFILLER_0_169_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11883_ _04975_ _05029_ _05052_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__or3_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _09375_ _09482_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__and2_1
X_13622_ _06600_ _06667_ _06686_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__or3_1
X_17390_ _10388_ _10389_ vssd1 vssd1 vccd1 vccd1 _10390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ net6632 net2475 _04288_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20347__79 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
XFILLER_0_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16341_ _08799_ _09258_ _09322_ _09320_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13553_ _06543_ _06554_ _06687_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__mux2_1
X_10765_ net2757 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _05035_ _05665_ _05669_ _05030_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a211o_1
X_19060_ net3038 _03009_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__or2_1
X_16272_ _09325_ _09326_ _09344_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__nand3_1
X_13484_ _06556_ _06595_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__or2_1
X_10696_ net2328 net6642 _04214_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__mux2_1
X_18011_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__xor2_2
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15223_ _08297_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__clkbuf_8
X_12435_ _05028_ _05576_ _05584_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ net4719 _08096_ _08249_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__mux2_1
X_12366_ rbzero.tex_g1\[55\] rbzero.tex_g1\[54\] _05219_ vssd1 vssd1 vccd1 vccd1 _05533_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14105_ _07255_ _07155_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ net6401 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19962_ net3952 _03471_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__nor2_1
X_15085_ net3356 _08201_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__or2_1
X_12297_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _05456_ vssd1 vssd1 vccd1 vccd1 _05465_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14036_ net528 _07185_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__and3_1
X_18913_ _02863_ net4459 net3700 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__or3b_1
X_11248_ net6710 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
X_19893_ net3853 _03515_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18844_ net4708 rbzero.wall_tracer.rayAddendY\[2\] vssd1 vssd1 vccd1 vccd1 _02833_
+ sky130_fd_sc_hd__xor2_1
X_11179_ net6816 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18775_ net3807 net2884 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15987_ _09042_ _09043_ _09061_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ _01652_ _01653_ _01655_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14938_ _08068_ _08084_ _08047_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__a21oi_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17657_ _01699_ _01708_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14869_ net7434 _08019_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16608_ _09674_ _09678_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _10130_ _09538_ vssd1 vssd1 vccd1 vccd1 _10586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19327_ net5158 _03159_ _03171_ _03168_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__o211a_1
X_16539_ _09610_ _09489_ _08632_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7217 rbzero.wall_tracer.trackDistX\[5\] vssd1 vssd1 vccd1 vccd1 net7741 sky130_fd_sc_hd__dlygate4sd3_1
X_19258_ _03036_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__clkbuf_4
Xhold7228 rbzero.debug_overlay.playerX\[-8\] vssd1 vssd1 vccd1 vccd1 net7752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6505 rbzero.tex_b0\[39\] vssd1 vssd1 vccd1 vccd1 net7029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ net3780 net4605 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__nand2_1
Xhold6516 net2161 vssd1 vssd1 vccd1 vccd1 net7040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6527 rbzero.tex_g1\[19\] vssd1 vssd1 vccd1 vccd1 net7051 sky130_fd_sc_hd__dlygate4sd3_1
X_19189_ net2995 net4081 _03084_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
Xhold6538 net2506 vssd1 vssd1 vccd1 vccd1 net7062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6549 net2221 vssd1 vssd1 vccd1 vccd1 net7073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5804 net627 vssd1 vssd1 vccd1 vccd1 net6328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5815 net761 vssd1 vssd1 vccd1 vccd1 net6339 sky130_fd_sc_hd__dlygate4sd3_1
X_21220_ clknet_leaf_43_i_clk net5493 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5826 rbzero.tex_b0\[20\] vssd1 vssd1 vccd1 vccd1 net6350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 _03469_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_1
Xhold112 net929 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5837 net996 vssd1 vssd1 vccd1 vccd1 net6361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 net7659 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5848 _04186_ vssd1 vssd1 vccd1 vccd1 net6372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5859 net1110 vssd1 vssd1 vccd1 vccd1 net6383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 net4950 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _03563_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__dlygate4sd3_1
X_21151_ net2983 _04132_ _04633_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a21oi_1
Xhold156 rbzero.wall_tracer.visualWallDist\[9\] vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_1
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold167 net4969 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 net4426 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
X_20102_ net1601 _03658_ net3328 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a21o_1
X_21082_ net4179 net4542 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__nand2_1
Xhold189 net3295 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20033_ net4424 net3543 _03594_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21984_ net209 net2318 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20935_ clknet_1_0__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__buf_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22467_ clknet_leaf_80_i_clk net4427 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12220_ net3876 _05371_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a21oi_1
X_21418_ clknet_leaf_85_i_clk net4770 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_22398_ net150 net1630 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12151_ _05297_ _05309_ _05318_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a31o_1
X_21349_ clknet_leaf_39_i_clk net4135 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11102_ net6844 net6664 _04426_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__mux2_1
X_20655__94 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__inv_2
X_12082_ _04982_ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__or2_1
Xhold690 net5717 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11033_ net6545 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__clkbuf_1
X_15910_ _08875_ _08984_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__nand2_1
X_16890_ net4509 _09937_ _09938_ _08152_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _08393_ _08625_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__nor2_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 _01574_ vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2091 _01164_ vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _02573_ _02574_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__or2_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ net3539 _08311_ _08305_ _08351_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__or4_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _06117_ _06121_ _06124_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1390 _00886_ vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
X_17511_ _08317_ _08634_ vssd1 vssd1 vccd1 vccd1 _10510_ sky130_fd_sc_hd__nor2_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935_ net3014 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__inv_2
X_14723_ _07852_ _07872_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ net3211 _02504_ _02508_ _02510_ _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a32o_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _10342_ _10441_ vssd1 vssd1 vccd1 vccd1 _10442_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_157_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14654_ _07304_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__clkbuf_4
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _04984_ _05031_ _05033_ _05035_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o211a_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _06754_ _06755_ _06661_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ net7284 net6796 _04277_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17373_ _10276_ _10344_ _10371_ vssd1 vssd1 vccd1 vccd1 _10373_ sky130_fd_sc_hd__nand3_1
X_14585_ _07717_ _07734_ _07735_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__a21oi_2
X_11797_ _04962_ _04965_ _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19112_ net6017 _03037_ _03046_ _03022_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__o211a_1
X_16324_ _09262_ _09397_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13536_ _06667_ _06686_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__nor2_8
XFILLER_0_83_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10748_ net51 net2367 _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ _08316_ _09328_ _09051_ _08701_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__a2bb2o_1
X_19043_ net1727 _02990_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__or2_1
X_13467_ _06424_ _06428_ _06540_ net82 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__o22a_2
XFILLER_0_168_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10679_ net6419 net7175 _04203_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _06381_ _08283_ _06267_ net1054 vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__a2bb2o_1
X_12418_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _05476_ vssd1 vssd1 vccd1 vccd1 _05585_
+ sky130_fd_sc_hd__mux2_1
X_16186_ _09259_ _09260_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13398_ _06545_ _06548_ _06540_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15137_ net4577 _06343_ net4342 vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__o21a_1
X_12349_ _05515_ _05516_ _04991_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3709 net7513 vssd1 vssd1 vccd1 vccd1 net4233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _08190_ _08192_ net3723 _01622_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__o211a_1
X_19945_ net4675 _03532_ net640 _03559_ _03083_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__a221o_1
X_14019_ _06895_ _06861_ _06885_ _06918_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__o22ai_2
X_19876_ net6155 _03479_ net745 _03502_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a211o_1
X_18827_ net6120 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18758_ net4620 net738 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__or2_1
X_17709_ _01668_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_136_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18689_ _02693_ _02694_ _02678_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20651_ net1578 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7003 rbzero.wall_tracer.trackDistY\[7\] vssd1 vssd1 vccd1 vccd1 net7527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7014 rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 net7538 sky130_fd_sc_hd__dlygate4sd3_1
X_20582_ _03924_ net3515 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7025 rbzero.wall_tracer.trackDistX\[-6\] vssd1 vssd1 vccd1 vccd1 net7549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22321_ net453 net2643 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold7036 rbzero.wall_tracer.trackDistX\[-7\] vssd1 vssd1 vccd1 vccd1 net7560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6302 net2108 vssd1 vssd1 vccd1 vccd1 net6826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7047 _02673_ vssd1 vssd1 vccd1 vccd1 net7571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6313 rbzero.tex_b0\[34\] vssd1 vssd1 vccd1 vccd1 net6837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7058 net4732 vssd1 vssd1 vccd1 vccd1 net7582 sky130_fd_sc_hd__buf_4
Xhold6324 net2082 vssd1 vssd1 vccd1 vccd1 net6848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6335 rbzero.tex_b1\[9\] vssd1 vssd1 vccd1 vccd1 net6859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22252_ net384 net2492 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold6346 net1901 vssd1 vssd1 vccd1 vccd1 net6870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5601 _08210_ vssd1 vssd1 vccd1 vccd1 net6125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6357 _04226_ vssd1 vssd1 vccd1 vccd1 net6881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5612 net3634 vssd1 vssd1 vccd1 vccd1 net6136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6368 net1985 vssd1 vssd1 vccd1 vccd1 net6892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5623 _08238_ vssd1 vssd1 vccd1 vccd1 net6147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6379 rbzero.tex_g1\[54\] vssd1 vssd1 vccd1 vccd1 net6903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5634 rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 net6158 sky130_fd_sc_hd__dlygate4sd3_1
X_21203_ net4956 net65 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__nor2_1
Xhold5645 rbzero.spi_registers.buf_texadd1\[7\] vssd1 vssd1 vccd1 vccd1 net6169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4900 net998 vssd1 vssd1 vccd1 vccd1 net5424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4911 net1043 vssd1 vssd1 vccd1 vccd1 net5435 sky130_fd_sc_hd__dlygate4sd3_1
X_22183_ net315 net1095 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold5656 net2256 vssd1 vssd1 vccd1 vccd1 net6180 sky130_fd_sc_hd__dlygate4sd3_1
X_20826__248 clknet_1_1__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__inv_2
Xhold5667 net4063 vssd1 vssd1 vccd1 vccd1 net6191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4922 rbzero.mapdxw\[1\] vssd1 vssd1 vccd1 vccd1 net5446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5678 net2533 vssd1 vssd1 vccd1 vccd1 net6202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4933 net1017 vssd1 vssd1 vccd1 vccd1 net5457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4944 _01174_ vssd1 vssd1 vccd1 vccd1 net5468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5689 net3893 vssd1 vssd1 vccd1 vccd1 net6213 sky130_fd_sc_hd__dlygate4sd3_1
X_21134_ net4136 net4679 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2_1
Xhold4955 net1079 vssd1 vssd1 vccd1 vccd1 net5479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4966 rbzero.wall_tracer.mapY\[9\] vssd1 vssd1 vccd1 vccd1 net5490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4977 _01052_ vssd1 vssd1 vccd1 vccd1 net5501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4988 rbzero.floor_leak\[0\] vssd1 vssd1 vccd1 vccd1 net5512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4999 net1118 vssd1 vssd1 vccd1 vccd1 net5523 sky130_fd_sc_hd__dlygate4sd3_1
X_21065_ _04059_ _04060_ _04058_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20016_ net1098 _03578_ net4413 _03602_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ net192 net2279 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _04836_ net2791 net2802 net4014 vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ clknet_leaf_95_i_clk net1279 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ net4001 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ net3992 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14370_ _06859_ _07359_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__or2_1
X_11582_ _04656_ _04666_ _04668_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ net4406 net6304 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__nand2_2
XFILLER_0_190_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16040_ _09107_ _09114_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ net4887 _06394_ _06393_ _06405_ vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12203_ _05341_ _05362_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nor2_2
XFILLER_0_161_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6880 _08341_ vssd1 vssd1 vccd1 vccd1 net7404 sky130_fd_sc_hd__buf_1
X_13183_ _06338_ _06307_ _06304_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_62_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12134_ _05194_ _05299_ _05200_ _05300_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17991_ _02038_ _02039_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19730_ net3038 _03407_ net5796 _03400_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12065_ _04978_ _05217_ _05223_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__o31a_1
X_16942_ _09946_ net4876 vssd1 vssd1 vccd1 vccd1 _09960_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ net6483 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__clkbuf_1
X_19661_ net6164 _03360_ net2091 _03371_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__o211a_1
X_16873_ _09931_ vssd1 vssd1 vccd1 vccd1 _09932_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18612_ _02607_ _02622_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__xnor2_1
X_15824_ _08422_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__inv_2
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ net5226 _03325_ _03331_ _03330_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__o211a_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ net4446 _02548_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__nand2_1
X_15755_ _08827_ _08828_ _08829_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__a21oi_2
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ net4600 net3090 vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__or2_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11918_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _05077_ vssd1 vssd1 vccd1 vccd1 _05088_
+ sky130_fd_sc_hd__mux2_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _07847_ _07848_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__or2_1
X_18474_ net3075 net3151 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__and2_2
X_15686_ _08347_ _08353_ _08367_ _08557_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ net141 _06052_ _06046_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _10422_ _10423_ _10424_ vssd1 vssd1 vccd1 vccd1 _10425_ sky130_fd_sc_hd__nand3_1
X_20931__343 clknet_1_1__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__inv_2
X_11849_ _04982_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__clkbuf_8
X_14637_ _07764_ _07786_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _09813_ _10236_ _10239_ _10237_ vssd1 vssd1 vccd1 vccd1 _10356_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14568_ _07704_ _07710_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__xor2_2
Xclkbuf_1_1__f__03994_ clknet_0__03994_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03994_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16307_ _09221_ _09233_ _09380_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__a21oi_2
X_13519_ _06519_ _06530_ _06631_ _06632_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__and4_1
X_17287_ _10286_ _10287_ vssd1 vssd1 vccd1 vccd1 _10288_ sky130_fd_sc_hd__xnor2_1
X_14499_ _07592_ _07594_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19026_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__buf_2
X_16238_ _09311_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4207 net1624 vssd1 vssd1 vccd1 vccd1 net4731 sky130_fd_sc_hd__dlygate4sd3_1
X_16169_ _08697_ _08745_ _09243_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__a21oi_1
Xhold4218 net2932 vssd1 vssd1 vccd1 vccd1 net4742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4229 _02642_ vssd1 vssd1 vccd1 vccd1 net4753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3506 _04130_ vssd1 vssd1 vccd1 vccd1 net4030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3517 net4051 vssd1 vssd1 vccd1 vccd1 net4041 sky130_fd_sc_hd__clkbuf_2
Xhold3528 net4041 vssd1 vssd1 vccd1 vccd1 net4052 sky130_fd_sc_hd__clkbuf_2
Xhold3539 net6190 vssd1 vssd1 vccd1 vccd1 net4063 sky130_fd_sc_hd__buf_2
XFILLER_0_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2805 _03665_ vssd1 vssd1 vccd1 vccd1 net3329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2816 _01215_ vssd1 vssd1 vccd1 vccd1 net3340 sky130_fd_sc_hd__dlygate4sd3_1
X_19928_ net2956 _03477_ _03532_ _03546_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2827 rbzero.pov.ready_buffer\[20\] vssd1 vssd1 vccd1 vccd1 net3351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2838 _03901_ vssd1 vssd1 vccd1 vccd1 net3362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2849 net7544 vssd1 vssd1 vccd1 vccd1 net3373 sky130_fd_sc_hd__dlygate4sd3_1
X_19859_ net2944 _08420_ _03484_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21821_ clknet_leaf_87_i_clk net3850 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21752_ clknet_leaf_1_i_clk net4330 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21683_ clknet_leaf_35_i_clk net5281 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdyw\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20634_ net4101 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20565_ net3732 net1209 _03911_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6110 net1778 vssd1 vssd1 vccd1 vccd1 net6634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6121 rbzero.tex_g1\[17\] vssd1 vssd1 vccd1 vccd1 net6645 sky130_fd_sc_hd__dlygate4sd3_1
X_22304_ net436 net1975 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6132 net1715 vssd1 vssd1 vccd1 vccd1 net6656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6143 _04429_ vssd1 vssd1 vccd1 vccd1 net6667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6154 net1765 vssd1 vssd1 vccd1 vccd1 net6678 sky130_fd_sc_hd__dlygate4sd3_1
X_20496_ _03858_ net3306 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6165 _04194_ vssd1 vssd1 vccd1 vccd1 net6689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5420 net2705 vssd1 vssd1 vccd1 vccd1 net5944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5431 net1971 vssd1 vssd1 vccd1 vccd1 net5955 sky130_fd_sc_hd__dlygate4sd3_1
X_22235_ net367 net2549 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold6176 net2064 vssd1 vssd1 vccd1 vccd1 net6700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6187 rbzero.tex_r0\[25\] vssd1 vssd1 vccd1 vccd1 net6711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5442 net2774 vssd1 vssd1 vccd1 vccd1 net5966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6198 net1847 vssd1 vssd1 vccd1 vccd1 net6722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5453 rbzero.map_overlay.i_mapdy\[2\] vssd1 vssd1 vccd1 vccd1 net5977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5464 rbzero.tex_g1\[53\] vssd1 vssd1 vccd1 vccd1 net5988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4730 rbzero.spi_registers.buf_otherx\[0\] vssd1 vssd1 vccd1 vccd1 net5254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5475 net2895 vssd1 vssd1 vccd1 vccd1 net5999 sky130_fd_sc_hd__dlygate4sd3_1
X_22166_ net298 net1928 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold5486 _03493_ vssd1 vssd1 vccd1 vccd1 net6010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4741 net990 vssd1 vssd1 vccd1 vccd1 net5265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5497 _01028_ vssd1 vssd1 vccd1 vccd1 net6021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4752 _00749_ vssd1 vssd1 vccd1 vccd1 net5276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4763 net1002 vssd1 vssd1 vccd1 vccd1 net5287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4774 net956 vssd1 vssd1 vccd1 vccd1 net5298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21117_ _04103_ _04104_ _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__or3_1
Xhold4785 rbzero.traced_texa\[-5\] vssd1 vssd1 vccd1 vccd1 net5309 sky130_fd_sc_hd__dlygate4sd3_1
X_22097_ clknet_leaf_6_i_clk net1579 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4796 net940 vssd1 vssd1 vccd1 vccd1 net5320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21048_ net5455 _03519_ _04014_ _04047_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a22o_1
X_13870_ _07011_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12821_ _04162_ net3993 net22 vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ net19 _05907_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__o21ai_1
X_15540_ _08166_ _08167_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__nand2_2
XFILLER_0_189_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ net2839 _04164_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _08295_ _08543_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__o21a_4
XFILLER_0_189_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ net11 net10 vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _10084_ _10086_ _10209_ _10210_ vssd1 vssd1 vccd1 vccd1 _10211_ sky130_fd_sc_hd__a211o_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _07568_ _07570_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nor2_1
X_11634_ net4099 vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18190_ _02112_ _02113_ _02150_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17141_ _10141_ _10142_ vssd1 vssd1 vccd1 vccd1 _10143_ sky130_fd_sc_hd__xnor2_1
X_14353_ _07502_ _07503_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11565_ _04724_ _04736_ _04691_ _04718_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ _06453_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17072_ net3399 _10067_ vssd1 vssd1 vccd1 vccd1 _10075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14284_ _07391_ _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11496_ _04654_ _04667_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16023_ _08493_ _09096_ _09095_ _09097_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_150_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ net4918 net3508 net4900 _04621_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ _06319_ net3209 vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ _05284_ _05285_ _05068_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__mux2_1
X_17974_ _01825_ _02022_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__xnor2_4
X_13097_ net4524 net4581 net4783 net673 vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19713_ net6236 _03395_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__or2_1
X_12048_ _05069_ _05214_ _05216_ _05061_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__o211a_1
X_16925_ net3379 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19644_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__buf_2
X_16856_ net3910 _09919_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15807_ _08880_ _08881_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_172_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19575_ _02998_ _03304_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__or2_1
X_16787_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09857_ sky130_fd_sc_hd__xnor2_1
X_13999_ _07111_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nor2_1
X_18526_ net4478 _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15738_ _08556_ net4954 vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__or2_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18457_ _02481_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__clkbuf_1
X_15669_ _08742_ _08743_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17408_ _09103_ _10406_ _09861_ _10407_ vssd1 vssd1 vccd1 vccd1 _10408_ sky130_fd_sc_hd__or4_1
X_18388_ _02414_ net3235 _02419_ _02420_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17339_ _10232_ _10233_ _10230_ vssd1 vssd1 vccd1 vccd1 _10339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19009_ net3885 net3904 _02973_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4004 net3494 vssd1 vssd1 vccd1 vccd1 net4528 sky130_fd_sc_hd__buf_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20281_ net3383 _03675_ _03769_ _03761_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4015 net7541 vssd1 vssd1 vccd1 vccd1 net4539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4026 _02761_ vssd1 vssd1 vccd1 vccd1 net4550 sky130_fd_sc_hd__dlygate4sd3_1
X_22020_ clknet_leaf_81_i_clk net3391 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4037 rbzero.debug_overlay.facingX\[0\] vssd1 vssd1 vccd1 vccd1 net4561 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold4048 net7490 vssd1 vssd1 vccd1 vccd1 net4572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3303 _03669_ vssd1 vssd1 vccd1 vccd1 net3827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3314 _05406_ vssd1 vssd1 vccd1 vccd1 net3838 sky130_fd_sc_hd__clkbuf_4
Xhold4059 _00426_ vssd1 vssd1 vccd1 vccd1 net4583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3325 _03590_ vssd1 vssd1 vccd1 vccd1 net3849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3336 _01005_ vssd1 vssd1 vccd1 vccd1 net3860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2602 _00811_ vssd1 vssd1 vccd1 vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3347 _00473_ vssd1 vssd1 vccd1 vccd1 net3871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2613 _00612_ vssd1 vssd1 vccd1 vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3358 _02733_ vssd1 vssd1 vccd1 vccd1 net3882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3369 net6212 vssd1 vssd1 vccd1 vccd1 net3893 sky130_fd_sc_hd__clkbuf_4
Xhold2624 net4392 vssd1 vssd1 vccd1 vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 _03528_ vssd1 vssd1 vccd1 vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1901 _04413_ vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2646 net4416 vssd1 vssd1 vccd1 vccd1 net3170 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1912 net7019 vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2657 _03245_ vssd1 vssd1 vccd1 vccd1 net3181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 _01491_ vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 _01180_ vssd1 vssd1 vccd1 vccd1 net3192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 net7084 vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2679 rbzero.row_render.size\[7\] vssd1 vssd1 vccd1 vccd1 net3551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1945 net6905 vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1956 _01403_ vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
X_20938__349 clknet_1_1__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__inv_2
Xhold1967 _04357_ vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 net7122 vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1989 _01127_ vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21804_ clknet_leaf_89_i_clk net2924 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21735_ clknet_leaf_23_i_clk net1870 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21666_ clknet_leaf_35_i_clk net5362 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20617_ net3965 net3979 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21597_ clknet_leaf_1_i_clk net4229 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11350_ net6840 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20548_ net3570 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ net5892 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20683__119 clknet_1_0__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__inv_2
X_20479_ net721 net3665 _03845_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5250 _00700_ vssd1 vssd1 vccd1 vccd1 net5774 sky130_fd_sc_hd__dlygate4sd3_1
X_13020_ _06138_ _06146_ _06151_ _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__and4bb_1
X_22218_ net350 net1528 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
Xhold5261 _00819_ vssd1 vssd1 vccd1 vccd1 net5785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5272 _03411_ vssd1 vssd1 vccd1 vccd1 net5796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5283 rbzero.map_overlay.i_otherx\[3\] vssd1 vssd1 vccd1 vccd1 net5807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5294 _04534_ vssd1 vssd1 vccd1 vccd1 net5818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4560 _00744_ vssd1 vssd1 vccd1 vccd1 net5084 sky130_fd_sc_hd__dlygate4sd3_1
X_22149_ net281 net2435 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
Xhold4571 net833 vssd1 vssd1 vccd1 vccd1 net5095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4582 net811 vssd1 vssd1 vccd1 vccd1 net5106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4593 net826 vssd1 vssd1 vccd1 vccd1 net5117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3870 rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 net4394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3881 net3161 vssd1 vssd1 vccd1 vccd1 net4405 sky130_fd_sc_hd__buf_1
X_14971_ _08092_ _08112_ _08113_ _08114_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__a31oi_2
Xhold3892 net7811 vssd1 vssd1 vccd1 vccd1 net4416 sky130_fd_sc_hd__dlygate4sd3_1
X_16710_ _09653_ _09767_ vssd1 vssd1 vccd1 vccd1 _09780_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__03997_ clknet_0__03997_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03997_
+ sky130_fd_sc_hd__clkbuf_16
X_13922_ net556 _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__xnor2_2
X_17690_ _10465_ _10466_ _10565_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16641_ _09693_ _09694_ _09710_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__nand3_1
X_13853_ _06998_ _06999_ _07002_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__nor3_1
XFILLER_0_187_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19360_ net4268 _03185_ _03190_ _03181_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__o211a_1
X_12804_ _05207_ _05957_ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16572_ _09642_ net3009 vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__and2_1
X_10996_ net2478 net7022 _04366_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__mux2_1
X_13784_ _06932_ _06934_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18311_ _02346_ _02347_ _02348_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15523_ net3046 _08312_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__and2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nor2_2
X_19291_ net5342 _03146_ _03151_ _03142_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__o211a_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18242_ _02216_ _02230_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__or2b_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _08373_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__clkbuf_4
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12666_ net6220 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14405_ _07554_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__nor2_1
X_11617_ _04768_ _04775_ _04777_ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a211o_1
X_18173_ _09231_ _09249_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__nor2_1
X_12597_ _05760_ _05761_ _04993_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__mux2_1
X_15385_ _08447_ _08459_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17124_ _09843_ _09844_ vssd1 vssd1 vccd1 vccd1 _10126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14336_ _07443_ _07486_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__xor2_1
X_11548_ _04718_ net3869 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold508 net6352 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
X_17055_ net3795 net3419 vssd1 vssd1 vccd1 vccd1 _10060_ sky130_fd_sc_hd__nand2_1
X_14267_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__or2_1
Xhold519 net5434 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ rbzero.spi_registers.texadd3\[10\] rbzero.spi_registers.texadd1\[10\] rbzero.spi_registers.texadd0\[10\]
+ rbzero.spi_registers.texadd2\[10\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__mux4_1
XFILLER_0_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16006_ _09070_ _09062_ _09069_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13218_ _06219_ net4897 net3804 net3984 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14198_ _07296_ _07298_ _07300_ _07258_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__a22o_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ net4433 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__inv_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 net6713 vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17957_ _02004_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__xnor2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1219 _01407_ vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_16908_ net4130 _09939_ _09940_ net6278 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__a22o_1
X_17888_ _09108_ _10406_ _01711_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__or3_1
X_19627_ net5140 net799 _03350_ _03343_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__o211a_1
X_16839_ net4288 net4105 net4088 vssd1 vssd1 vccd1 vccd1 _09909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19558_ net3100 _03305_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18509_ net628 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ net1608 _03265_ net5755 _03260_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__o211a_1
X_21520_ clknet_leaf_34_i_clk net5119 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21451_ clknet_leaf_46_i_clk net3267 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20402_ net2833 net3660 _03801_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21382_ clknet_leaf_58_i_clk _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20333_ clknet_1_1__leaf__03773_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20989__16 clknet_1_1__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
X_20264_ _08275_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3100 _08287_ vssd1 vssd1 vccd1 vccd1 net3624 sky130_fd_sc_hd__dlygate4sd3_1
X_22003_ net228 net1931 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold3111 _00432_ vssd1 vssd1 vccd1 vccd1 net3635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3122 net1322 vssd1 vssd1 vccd1 vccd1 net3646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3133 _03608_ vssd1 vssd1 vccd1 vccd1 net3657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3144 _01211_ vssd1 vssd1 vccd1 vccd1 net3668 sky130_fd_sc_hd__dlygate4sd3_1
X_20195_ _03440_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__clkbuf_4
Xhold2410 net5464 vssd1 vssd1 vccd1 vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3155 net1199 vssd1 vssd1 vccd1 vccd1 net3679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3166 net4698 vssd1 vssd1 vccd1 vccd1 net3690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2421 _03494_ vssd1 vssd1 vccd1 vccd1 net2945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3177 _03647_ vssd1 vssd1 vccd1 vccd1 net3701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2432 rbzero.pov.ready_buffer\[50\] vssd1 vssd1 vccd1 vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2443 _00690_ vssd1 vssd1 vccd1 vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3188 _01207_ vssd1 vssd1 vccd1 vccd1 net3712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2454 _02524_ vssd1 vssd1 vccd1 vccd1 net2978 sky130_fd_sc_hd__buf_2
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1720 _04458_ vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3199 _08194_ vssd1 vssd1 vccd1 vccd1 net3723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2465 net6026 vssd1 vssd1 vccd1 vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1731 _01443_ vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2476 _03499_ vssd1 vssd1 vccd1 vccd1 net3000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1742 _04409_ vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2487 net618 vssd1 vssd1 vccd1 vccd1 net3011 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_99_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1753 net6803 vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2498 net612 vssd1 vssd1 vccd1 vccd1 net3022 sky130_fd_sc_hd__buf_2
Xhold1764 rbzero.tex_b0\[57\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1775 _04195_ vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1786 net7100 vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1797 _01275_ vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10850_ net6702 net6437 _04288_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ net7233 net7203 _04255_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _05680_ _05682_ _05685_ _05061_ net81 vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21718_ clknet_leaf_8_i_clk net3013 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _05062_ _05004_ _05097_ _05104_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21649_ clknet_leaf_33_i_clk net2592 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11402_ net6598 net2215 _04584_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15170_ _08263_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__clkbuf_1
X_12382_ _05461_ _05548_ _05023_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_90 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _07270_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__xor2_1
X_11333_ net6728 net6592 _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20295__32 clknet_1_1__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
XFILLER_0_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ net552 _06918_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__or2_1
X_11264_ net2858 net7187 _04514_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13003_ _06098_ _06101_ _06103_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a21o_1
Xhold5080 rbzero.spi_registers.texadd3\[7\] vssd1 vssd1 vccd1 vccd1 net5604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5091 _00743_ vssd1 vssd1 vccd1 vccd1 net5615 sky130_fd_sc_hd__dlygate4sd3_1
X_18860_ net3700 net4799 _02846_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__o21ai_1
X_11195_ net2189 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
X_17811_ _01859_ _01860_ _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a21o_2
Xhold4390 _06347_ vssd1 vssd1 vccd1 vccd1 net4914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _04632_ _02777_ _02778_ _02783_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _01791_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__nor2_1
X_14954_ _06664_ _08054_ _08090_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _07053_ _07055_ _07051_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__a21o_1
X_17673_ _10529_ _10552_ _10550_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ _07991_ _07997_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19412_ _03141_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__clkbuf_4
X_16624_ _08351_ _08352_ vssd1 vssd1 vccd1 vccd1 _09695_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ _06866_ _06886_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19343_ _03141_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__clkbuf_4
X_16555_ _09581_ _09626_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_175_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10979_ _04332_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__clkbuf_4
X_13767_ _06914_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ net3162 _08328_ _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__a22oi_4
X_12718_ net14 _05875_ _05878_ _05869_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__a22o_1
X_19274_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__buf_2
XFILLER_0_210_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16486_ _09535_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13698_ _06833_ _06848_ _06678_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18225_ _02246_ _02247_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__nor2_1
X_15437_ _08317_ _08326_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ net53 _05786_ _05796_ net40 vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6709 net2499 vssd1 vssd1 vccd1 vccd1 net7233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _02086_ _02110_ _02201_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__nand3_1
X_15368_ net3008 _08381_ _08442_ _06209_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ _09251_ _08962_ vssd1 vssd1 vccd1 vccd1 _10109_ sky130_fd_sc_hd__or2b_1
Xhold305 net6344 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ _07268_ _07467_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__nand2_2
Xhold316 net7514 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ _01675_ _09310_ _02133_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15299_ _08347_ _08353_ _08367_ _08373_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold327 net4735 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold338 net5141 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _10041_ _10044_ vssd1 vssd1 vccd1 vccd1 _10045_ sky130_fd_sc_hd__nor2_1
Xhold349 net5335 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03776_ _03776_ vssd1 vssd1 vccd1 vccd1 clknet_0__03776_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_180_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ net6140 _02963_ _09999_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__mux2_1
Xhold1005 net5720 vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 net6523 vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1027 net6577 vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1038 rbzero.spi_registers.buf_texadd2\[14\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 net5730 vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21503_ clknet_leaf_14_i_clk net2803 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21434_ clknet_leaf_82_i_clk net4629 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21365_ clknet_leaf_54_i_clk _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold850 _01311_ vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
X_21296_ clknet_leaf_74_i_clk net4089 vssd1 vssd1 vccd1 vccd1 rbzero.side_hot sky130_fd_sc_hd__dfxtp_1
Xhold861 _01292_ vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold872 net5694 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
X_20247_ net5665 _03744_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or2_1
Xhold883 _03197_ vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 net6478 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ net5544 _03705_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__or2_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2240 _01445_ vssd1 vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2251 net5967 vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2262 _01277_ vssd1 vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2273 _04505_ vssd1 vssd1 vccd1 vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2284 net4878 vssd1 vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 net6747 vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2295 rbzero.tex_r1\[56\] vssd1 vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1561 rbzero.tex_r1\[14\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ net3144 net915 _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1572 _00914_ vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 net6823 vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1594 _01340_ vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_107 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_107/HI o_rgb[21]
+ sky130_fd_sc_hd__conb_1
X_10902_ net2453 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_118 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_118/HI zeros[10]
+ sky130_fd_sc_hd__conb_1
X_11882_ _05030_ _05036_ _05041_ _05049_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__o311a_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _07776_ _07773_ _07775_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__nand3_1
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_129 vssd1 vssd1 vccd1 vccd1 ones[5] top_ew_algofoogle_129/LO sky130_fd_sc_hd__conb_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10833_ net6405 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__clkbuf_1
X_13621_ _06768_ _06771_ _06743_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _09398_ _09400_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10764_ net7282 net7243 _04244_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__mux2_1
X_13552_ _06612_ _06552_ _06695_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _05279_ _05666_ _05668_ _05461_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__o211a_1
X_16271_ _09325_ _09326_ _09344_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__a21o_1
X_13483_ _06591_ _06609_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__nor2_1
X_10695_ net2374 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20689__125 clknet_1_1__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__inv_2
X_18010_ _01909_ _01952_ _01950_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a21oi_2
X_12434_ _05030_ _05588_ _05592_ _05051_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__o311a_1
X_15222_ net3535 _06207_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15153_ _08254_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12365_ _05532_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11316_ net6399 net2346 _04540_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__mux2_1
X_14104_ _07153_ _07151_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__or2b_1
X_19961_ _03502_ net3083 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__nor2_1
X_15084_ net4556 net4511 _08191_ vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__mux2_1
X_12296_ _05229_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ _07111_ _07149_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__xor2_1
X_18912_ _02893_ _02894_ _02895_ _02896_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a22o_1
X_11247_ net1880 net6708 _04503_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__mux2_1
X_19892_ net6210 _03479_ net726 _03519_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__a211o_1
X_18843_ _02529_ net4710 _02823_ net3862 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a31o_1
X_11178_ net2249 net6814 _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__mux2_1
X_18774_ _02760_ net4550 _02762_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__o21a_1
X_15986_ _09054_ _09059_ _09060_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17725_ _01774_ _01775_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_171_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ net7759 _08083_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__and2_1
XFILLER_0_171_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17656_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868_ _07918_ _08018_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16607_ _09547_ _09675_ _09677_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__o21a_1
X_13819_ _06885_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__buf_2
X_17587_ _10528_ _10506_ vssd1 vssd1 vccd1 vccd1 _10585_ sky130_fd_sc_hd__or2b_1
XFILLER_0_175_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14799_ _07935_ _07946_ _07949_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__a21oi_1
X_19326_ net4672 _03160_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16538_ net3185 _08628_ vssd1 vssd1 vccd1 vccd1 _09610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19257_ net4127 _03119_ net607 _03128_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__o211a_1
Xhold7207 rbzero.debug_overlay.playerX\[-6\] vssd1 vssd1 vccd1 vccd1 net7731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16469_ _09421_ _09540_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7218 net4432 vssd1 vssd1 vccd1 vccd1 net7742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_183_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7229 rbzero.texu_hot\[4\] vssd1 vssd1 vccd1 vccd1 net7753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18208_ _02252_ _02253_ _09999_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a21oi_2
Xhold6506 net2399 vssd1 vssd1 vccd1 vccd1 net7030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6517 rbzero.tex_b1\[50\] vssd1 vssd1 vccd1 vccd1 net7041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19188_ net5068 _03078_ _03091_ _03074_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6528 net2357 vssd1 vssd1 vccd1 vccd1 net7052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6539 rbzero.tex_g0\[58\] vssd1 vssd1 vccd1 vccd1 net7063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _02184_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5805 gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 net6329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5816 gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5827 net1031 vssd1 vssd1 vccd1 vccd1 net6351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _00954_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5838 rbzero.spi_registers.sclk_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _03059_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5849 net1041 vssd1 vssd1 vccd1 vccd1 net6373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _03444_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 net4952 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ net6168 net3535 _08200_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold146 net4388 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 net4137 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ net3328 net4865 net4797 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and3_1
Xhold168 rbzero.wall_tracer.visualWallDist\[-3\] vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold179 net5029 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
X_21081_ net4179 net4542 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20032_ net3878 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__clkbuf_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21983_ net208 net2532 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22466_ clknet_leaf_69_i_clk net1129 vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21417_ clknet_leaf_78_i_clk net3372 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22397_ net149 net2226 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12150_ _04880_ _04904_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__nand2_1
X_21348_ clknet_leaf_39_i_clk net4178 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11101_ net2129 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_13_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12081_ rbzero.tex_r1\[47\] rbzero.tex_r1\[46\] _05070_ vssd1 vssd1 vccd1 vccd1 _05250_
+ sky130_fd_sc_hd__mux2_1
X_21279_ clknet_leaf_59_i_clk _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold680 net5550 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold691 _03196_ vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net6543 net2659 _04392_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
X_20803__227 clknet_1_0__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__inv_2
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _08846_ _08848_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2070 _03380_ vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2081 net6809 vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 net7092 vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _08373_ _08625_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__nor2_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _06125_ _06127_ _06131_ _06129_ _06128_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__o2111a_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _08329_ _10380_ vssd1 vssd1 vccd1 vccd1 _10509_ sky130_fd_sc_hd__nor2_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1380 _03431_ vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1391 net5801 vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_19_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14722_ _07852_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11934_ net3014 _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or2_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ net3747 _02504_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nand2_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _10439_ _10440_ vssd1 vssd1 vccd1 vccd1 _10441_ sky130_fd_sc_hd__and2b_1
XFILLER_0_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _07367_ _07590_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__or2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__clkbuf_8
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _06638_ _06687_ _06718_ _06691_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__a211o_1
X_17372_ _10276_ _10344_ _10371_ vssd1 vssd1 vccd1 vccd1 _10372_ sky130_fd_sc_hd__a21o_1
X_10816_ net7151 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11796_ _04918_ _04920_ _04964_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a21oi_1
X_14584_ _07733_ _07718_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19111_ net5459 _03040_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__or2_1
X_16323_ _09395_ _09396_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ _06681_ _06683_ _06624_ _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__04800_ _04800_ vssd1 vssd1 vccd1 vccd1 clknet_0__04800_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19042_ net1727 _02988_ net3942 _02993_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__o211a_1
X_16254_ _08409_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ net6762 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__clkbuf_1
X_13466_ _06433_ _06415_ _06419_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__a21o_2
XFILLER_0_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _06382_ _06359_ _06267_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__o21bai_1
X_12417_ _05578_ _05580_ _05583_ _05062_ _04979_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a221o_1
X_16185_ _08799_ _09258_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__or2_1
X_13397_ net6123 _06431_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ _06386_ net3692 net4780 _08239_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _05493_ vssd1 vssd1 vccd1 vccd1 _05516_
+ sky130_fd_sc_hd__mux2_1
X_12279_ _05447_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
X_19944_ net4675 _03553_ _03558_ _03529_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__a22o_1
X_15067_ _08195_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__clkbuf_4
X_14018_ net552 _06922_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__nor2_1
X_19875_ net744 _03485_ _03474_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__o211a_1
X_20743__174 clknet_1_0__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__inv_2
X_18826_ rbzero.wall_tracer.rayAddendY\[0\] _02816_ _02714_ vssd1 vssd1 vccd1 vccd1
+ _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18757_ net4438 net723 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__nand2_1
X_15969_ _08432_ _09021_ _08625_ _09022_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__or4b_1
XFILLER_0_175_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17708_ _10594_ _10595_ _10592_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18688_ _02647_ _05401_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17639_ _01688_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20650_ net6557 _03026_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19309_ net1625 _03160_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20581_ net744 net3514 net3250 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__mux2_1
Xhold7004 rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 net7528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7015 rbzero.wall_tracer.trackDistY\[-6\] vssd1 vssd1 vccd1 vccd1 net7539 sky130_fd_sc_hd__dlygate4sd3_1
X_22320_ net452 net2670 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7026 rbzero.wall_tracer.trackDistX\[-5\] vssd1 vssd1 vccd1 vccd1 net7550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7037 rbzero.wall_tracer.trackDistY\[-9\] vssd1 vssd1 vccd1 vccd1 net7561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6303 rbzero.tex_r0\[37\] vssd1 vssd1 vccd1 vccd1 net6827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7048 _02675_ vssd1 vssd1 vccd1 vccd1 net7572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6314 net2331 vssd1 vssd1 vccd1 vccd1 net6838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7059 _00001_ vssd1 vssd1 vccd1 vccd1 net7583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6325 rbzero.tex_g1\[29\] vssd1 vssd1 vccd1 vccd1 net6849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22251_ net383 net1867 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold6336 net2319 vssd1 vssd1 vccd1 vccd1 net6860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6347 rbzero.tex_b0\[33\] vssd1 vssd1 vccd1 vccd1 net6871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5602 rbzero.debug_overlay.playerY\[-4\] vssd1 vssd1 vccd1 vccd1 net6126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6358 net2086 vssd1 vssd1 vccd1 vccd1 net6882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6369 rbzero.tex_g1\[22\] vssd1 vssd1 vccd1 vccd1 net6893 sky130_fd_sc_hd__dlygate4sd3_1
X_21202_ net941 _02528_ _02579_ net4802 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a22o_1
Xhold5624 net3627 vssd1 vssd1 vccd1 vccd1 net6148 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22182_ net314 net2742 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5646 net2090 vssd1 vssd1 vccd1 vccd1 net6170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4901 _01594_ vssd1 vssd1 vccd1 vccd1 net5425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5657 rbzero.debug_overlay.playerX\[2\] vssd1 vssd1 vccd1 vccd1 net6181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4912 _00781_ vssd1 vssd1 vccd1 vccd1 net5436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5668 _00976_ vssd1 vssd1 vccd1 vccd1 net6192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4923 net1008 vssd1 vssd1 vccd1 vccd1 net5447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4934 rbzero.spi_registers.buf_othery\[0\] vssd1 vssd1 vccd1 vccd1 net5458 sky130_fd_sc_hd__dlygate4sd3_1
X_21133_ net4136 net4679 vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__nand2_2
Xhold4945 net1071 vssd1 vssd1 vccd1 vccd1 net5469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4956 net5484 vssd1 vssd1 vccd1 vccd1 net5480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4967 net2907 vssd1 vssd1 vccd1 vccd1 net5491 sky130_fd_sc_hd__buf_1
Xhold4978 net1106 vssd1 vssd1 vccd1 vccd1 net5502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4989 net1113 vssd1 vssd1 vccd1 vccd1 net5513 sky130_fd_sc_hd__dlygate4sd3_1
X_21064_ _04058_ _04059_ _04060_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nand3_1
X_20015_ rbzero.debug_overlay.facingY\[-4\] _03582_ vssd1 vssd1 vccd1 vccd1 _03609_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_193_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ net191 net1444 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ clknet_leaf_95_i_clk net1382 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _04818_ net3535 net2 vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__o21a_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10601_ _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11581_ _04160_ _04672_ _04750_ _04752_ _04718_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a311o_1
XFILLER_0_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ _06432_ _06434_ _06470_ net4947 vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13251_ _06401_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xor2_1
X_22449_ clknet_leaf_66_i_clk _01618_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _05347_ _05351_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13182_ _06327_ _06334_ _06337_ _06322_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__o2bb2a_1
Xhold6881 _08381_ vssd1 vssd1 vccd1 vccd1 net7405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ net4059 _04759_ _05301_ _04606_ net4014 vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a32o_1
X_17990_ _09231_ _08705_ _02037_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12064_ _05034_ _05226_ _05228_ _05232_ _05022_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a221o_1
X_16941_ _09947_ _09948_ _09957_ net4875 vssd1 vssd1 vccd1 vccd1 _09959_ sky130_fd_sc_hd__a31o_1
XFILLER_0_198_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11015_ net6481 net2442 _04377_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__mux2_1
X_19660_ _03294_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__clkbuf_4
X_16872_ _04622_ _09930_ vssd1 vssd1 vccd1 vccd1 _09931_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18611_ _02620_ _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__nand2_1
X_15823_ _08860_ _08896_ _08897_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__nand3_2
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19591_ net3957 _03327_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__or2_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ net6243 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__clkbuf_1
X_15754_ _08807_ _08826_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__nor2_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ net4600 net3090 vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__nand2_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _07828_ _07827_ _07820_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11917_ _05085_ _05086_ _04992_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__mux2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ net3150 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__clkbuf_1
X_15685_ _08752_ _08759_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ net54 net55 net57 net56 _06046_ _06052_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _10297_ _10302_ _10301_ vssd1 vssd1 vccd1 vccd1 _10424_ sky130_fd_sc_hd__a21bo_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14636_ _07764_ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__xor2_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _04994_ vssd1 vssd1 vccd1 vccd1 _05018_
+ sky130_fd_sc_hd__mux2_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _10353_ _10354_ vssd1 vssd1 vccd1 vccd1 _10355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14567_ _07670_ _07679_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__xor2_2
Xclkbuf_1_1__f__03993_ clknet_0__03993_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03993_
+ sky130_fd_sc_hd__clkbuf_16
X_11779_ net924 net1364 net1456 net1072 vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a22o_1
X_16306_ _09230_ _09232_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ _06619_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__inv_2
X_17286_ _08684_ _09595_ vssd1 vssd1 vccd1 vccd1 _10287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ _07647_ _07648_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__or2_2
X_19025_ _08274_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__clkbuf_8
X_16237_ _08313_ _09310_ vssd1 vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__or2_2
X_13449_ _06598_ _06599_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_207_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16168_ _08655_ _08696_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4208 net3121 vssd1 vssd1 vccd1 vccd1 net4732 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4219 rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 net4743 sky130_fd_sc_hd__dlygate4sd3_1
X_15119_ net6098 _08223_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__or2_1
Xhold3507 _01611_ vssd1 vssd1 vccd1 vccd1 net4031 sky130_fd_sc_hd__dlygate4sd3_1
X_16099_ _08997_ _09078_ _09171_ _09173_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__o22a_2
XFILLER_0_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3518 _05199_ vssd1 vssd1 vccd1 vccd1 net4042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3529 _04164_ vssd1 vssd1 vccd1 vccd1 net4053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2806 _03666_ vssd1 vssd1 vccd1 vccd1 net3330 sky130_fd_sc_hd__dlygate4sd3_1
X_19927_ _08436_ _03476_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2817 rbzero.pov.spi_buffer\[50\] vssd1 vssd1 vccd1 vccd1 net3341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2828 net1226 vssd1 vssd1 vccd1 vccd1 net3352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2839 _01228_ vssd1 vssd1 vccd1 vccd1 net3363 sky130_fd_sc_hd__dlygate4sd3_1
X_19858_ net2935 _03475_ net6010 _03454_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__o211a_1
X_18809_ net7576 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__inv_2
X_19789_ net3038 _03442_ net1990 _03441_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__o211a_1
X_21820_ clknet_leaf_87_i_clk net3875 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21751_ clknet_leaf_0_i_clk net1640 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20702_ clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__buf_1
XFILLER_0_153_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21682_ clknet_leaf_35_i_clk net5245 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdyw\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20633_ net4061 _08275_ net4100 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__and3b_1
XFILLER_0_188_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20564_ net3707 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6100 net1903 vssd1 vssd1 vccd1 vccd1 net6624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6111 rbzero.tex_g1\[15\] vssd1 vssd1 vccd1 vccd1 net6635 sky130_fd_sc_hd__dlygate4sd3_1
X_22303_ net435 net1260 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6122 net1771 vssd1 vssd1 vccd1 vccd1 net6646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6133 _04447_ vssd1 vssd1 vccd1 vccd1 net6657 sky130_fd_sc_hd__dlygate4sd3_1
X_20495_ net3305 net1318 _03867_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6144 net1945 vssd1 vssd1 vccd1 vccd1 net6668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6155 _04412_ vssd1 vssd1 vccd1 vccd1 net6679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5410 rbzero.tex_g0\[0\] vssd1 vssd1 vccd1 vccd1 net5934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22234_ net366 net2480 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold6166 net1854 vssd1 vssd1 vccd1 vccd1 net6690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5421 _00656_ vssd1 vssd1 vccd1 vccd1 net5945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5432 gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 net5956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6177 rbzero.tex_r0\[15\] vssd1 vssd1 vccd1 vccd1 net6701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6188 net2054 vssd1 vssd1 vccd1 vccd1 net6712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5443 _00666_ vssd1 vssd1 vccd1 vccd1 net5967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6199 rbzero.tex_b0\[45\] vssd1 vssd1 vccd1 vccd1 net6723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5454 net2789 vssd1 vssd1 vccd1 vccd1 net5978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5465 net1554 vssd1 vssd1 vccd1 vccd1 net5989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4720 _00851_ vssd1 vssd1 vccd1 vccd1 net5244 sky130_fd_sc_hd__dlygate4sd3_1
X_22165_ net297 net2351 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold5476 _00667_ vssd1 vssd1 vccd1 vccd1 net6000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4731 net937 vssd1 vssd1 vccd1 vccd1 net5255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5487 _00959_ vssd1 vssd1 vccd1 vccd1 net6011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4742 rbzero.spi_registers.texadd1\[2\] vssd1 vssd1 vccd1 vccd1 net5266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4753 net944 vssd1 vssd1 vccd1 vccd1 net5277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5498 rbzero.row_render.size\[4\] vssd1 vssd1 vccd1 vccd1 net6022 sky130_fd_sc_hd__dlygate4sd3_1
X_21116_ net4160 net4653 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__and2_1
Xhold4764 _00797_ vssd1 vssd1 vccd1 vccd1 net5288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4775 _00730_ vssd1 vssd1 vccd1 vccd1 net5299 sky130_fd_sc_hd__dlygate4sd3_1
X_22096_ clknet_leaf_6_i_clk net1174 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4786 net884 vssd1 vssd1 vccd1 vccd1 net5310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4797 rbzero.spi_registers.buf_mapdxw\[0\] vssd1 vssd1 vccd1 vccd1 net5321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21047_ _04043_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ _05976_ _05978_ net25 vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915__328 clknet_1_1__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__inv_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ net19 _05908_ _05910_ net18 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21949_ net174 net1622 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ net2839 _04164_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _08300_ _06482_ _08320_ _08544_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__a211o_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ net13 net12 vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14421_ _07562_ _07571_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__and2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ net4020 net3897 net3964 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _08717_ _08574_ vssd1 vssd1 vccd1 vccd1 _10142_ sky130_fd_sc_hd__nor2_1
X_14352_ _07495_ _07501_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11564_ _04690_ _04689_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17071_ _10074_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14283_ _07432_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__and2_2
X_11495_ rbzero.texu_hot\[3\] _04653_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__or2_1
X_16022_ _09051_ _08755_ _09094_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7390 rbzero.wall_tracer.stepDistX\[10\] vssd1 vssd1 vccd1 vccd1 net7914 sky130_fd_sc_hd__dlygate4sd3_1
X_13234_ net3507 net4910 vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__nor2_1
X_20809__233 clknet_1_0__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__inv_2
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ _06319_ net3209 _06320_ net3554 vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ rbzero.tex_r1\[25\] rbzero.tex_r1\[24\] _05230_ vssd1 vssd1 vccd1 vccd1 _05285_
+ sky130_fd_sc_hd__mux2_1
X_17973_ _09582_ _02021_ _01940_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_2
X_13096_ net3772 net3718 net3627 net3222 vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or4_1
XFILLER_0_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12047_ _05002_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__or2_1
X_16924_ _04693_ net3378 _09943_ vssd1 vssd1 vccd1 vccd1 _09944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19712_ _03000_ _03393_ net2114 _03400_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__o211a_1
X_16855_ net3989 _09921_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__nor2_1
X_19643_ _02491_ _02514_ _02498_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__and3_2
X_15806_ _08512_ _08522_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__xnor2_1
X_19574_ net5322 _03302_ _03319_ _03314_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16786_ _09103_ _09595_ vssd1 vssd1 vccd1 vccd1 _09856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _07119_ _07147_ _07148_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__a21boi_2
X_18525_ _02541_ _02542_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__or2b_1
X_15737_ _08353_ _08625_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__nor2_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12949_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20855__275 clknet_1_0__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__inv_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _02480_ net3742 net4920 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_2
X_15668_ _08691_ _08723_ _08741_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__nand3_1
XFILLER_0_146_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _10152_ vssd1 vssd1 vccd1 vccd1 _10407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14619_ _07747_ _07748_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__or2_1
X_18387_ net4536 net4372 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _08564_ _08387_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17338_ _10252_ _10220_ vssd1 vssd1 vccd1 vccd1 _10338_ sky130_fd_sc_hd__or2b_1
XFILLER_0_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _10139_ _10140_ vssd1 vssd1 vccd1 vccd1 _10270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008_ net3906 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20280_ net3496 _03678_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4005 net7814 vssd1 vssd1 vccd1 vccd1 net4529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4016 net3460 vssd1 vssd1 vccd1 vccd1 net4540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4027 _02763_ vssd1 vssd1 vccd1 vccd1 net4551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4038 _03597_ vssd1 vssd1 vccd1 vccd1 net4562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4049 net3501 vssd1 vssd1 vccd1 vccd1 net4573 sky130_fd_sc_hd__buf_1
Xhold3304 _01033_ vssd1 vssd1 vccd1 vccd1 net3828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3315 _03626_ vssd1 vssd1 vccd1 vccd1 net3839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3326 _00990_ vssd1 vssd1 vccd1 vccd1 net3850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2603 net4379 vssd1 vssd1 vccd1 vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2614 net7781 vssd1 vssd1 vccd1 vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3359 _02734_ vssd1 vssd1 vccd1 vccd1 net3883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2625 net7595 vssd1 vssd1 vccd1 vccd1 net3149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2636 _00969_ vssd1 vssd1 vccd1 vccd1 net3160 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1902 _01370_ vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2647 net4713 vssd1 vssd1 vccd1 vccd1 net3171 sky130_fd_sc_hd__clkbuf_2
Xhold1913 _04522_ vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 _03246_ vssd1 vssd1 vccd1 vccd1 net3182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 rbzero.tex_b1\[63\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2669 net7826 vssd1 vssd1 vccd1 vccd1 net3193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1935 _04302_ vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1946 net6907 vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1957 net6805 vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 _01421_ vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1979 _04545_ vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21803_ clknet_leaf_89_i_clk net4895 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21734_ clknet_leaf_22_i_clk net1789 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21665_ clknet_leaf_35_i_clk net5304 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20616_ _09929_ net4017 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21596_ clknet_leaf_1_i_clk net4246 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20547_ _03902_ net3569 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ net5841 net5890 _04514_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20478_ net3414 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
Xhold5240 _00924_ vssd1 vssd1 vccd1 vccd1 net5764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5251 rbzero.tex_r0\[1\] vssd1 vssd1 vccd1 vccd1 net5775 sky130_fd_sc_hd__dlygate4sd3_1
X_22217_ net349 net2661 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5262 net1728 vssd1 vssd1 vccd1 vccd1 net5786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5273 _00913_ vssd1 vssd1 vccd1 vccd1 net5797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5284 net2043 vssd1 vssd1 vccd1 vccd1 net5808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5295 net1968 vssd1 vssd1 vccd1 vccd1 net5819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4550 net770 vssd1 vssd1 vccd1 vccd1 net5074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22148_ net280 net2251 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
Xhold4561 net879 vssd1 vssd1 vccd1 vccd1 net5085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4572 _00875_ vssd1 vssd1 vccd1 vccd1 net5096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4583 _00798_ vssd1 vssd1 vccd1 vccd1 net5107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4594 _00689_ vssd1 vssd1 vccd1 vccd1 net5118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3860 net1393 vssd1 vssd1 vccd1 vccd1 net4384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3871 net711 vssd1 vssd1 vccd1 vccd1 net4395 sky130_fd_sc_hd__dlygate4sd3_1
X_22079_ clknet_leaf_13_i_clk net3253 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_14970_ net7458 _08071_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__and2_1
Xhold3882 rbzero.debug_overlay.facingX\[10\] vssd1 vssd1 vccd1 vccd1 net4406 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3893 net3170 vssd1 vssd1 vccd1 vccd1 net4417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03996_ clknet_0__03996_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03996_
+ sky130_fd_sc_hd__clkbuf_16
X_13921_ _07032_ _07035_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16640_ _09693_ _09694_ _09710_ vssd1 vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _06998_ _06999_ _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ net40 _05956_ _05958_ net41 vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a22o_1
X_16571_ net4063 net3008 _08293_ vssd1 vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__mux2_1
X_13783_ _06880_ _06886_ _06933_ _06931_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__o2bb2a_1
X_10995_ net2877 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__clkbuf_1
X_18310_ _02352_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__clkbuf_1
X_15522_ net3169 _08298_ _06209_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__o21a_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12734_ net19 net18 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__nor2_1
X_19290_ net1829 _03147_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _02285_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__xnor2_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _08527_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__inv_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12665_ net6041 vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _07551_ _07552_ _07553_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18172_ _02096_ _02097_ _02218_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ _04727_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ _08448_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__nand2_1
X_12596_ rbzero.tex_b1\[11\] rbzero.tex_b1\[10\] _04988_ vssd1 vssd1 vccd1 vccd1 _05761_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17123_ _10093_ _10124_ vssd1 vssd1 vccd1 vccd1 _10125_ sky130_fd_sc_hd__xnor2_1
X_14335_ _07465_ _07469_ _07476_ _07485_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11547_ net3868 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__inv_2
Xhold509 _01129_ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ net3795 net3419 vssd1 vssd1 vccd1 vccd1 _10059_ sky130_fd_sc_hd__nor2_1
X_14266_ _07376_ _07379_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__or2b_1
X_11478_ rbzero.texu_hot\[5\] _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16005_ _09070_ _09062_ _09069_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__and3_1
XFILLER_0_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13217_ _06213_ _06190_ _06183_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__a21o_1
X_14197_ _07346_ _07347_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__xnor2_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _06300_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__and2_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17956_ _10380_ _09310_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__nor2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ net4387 _06190_ net4912 _04822_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a2bb2o_1
Xhold1209 _04265_ vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16907_ net4146 _09939_ _09940_ net6253 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22o_1
X_17887_ _09582_ _10539_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__or2_1
X_19626_ net3109 _03340_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__or2_1
X_16838_ _09781_ _09907_ vssd1 vssd1 vccd1 vccd1 _09908_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ _08873_ _08574_ vssd1 vssd1 vccd1 vccd1 _09839_ sky130_fd_sc_hd__or2_1
X_19557_ net930 _03303_ _03310_ _03295_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18508_ net6328 _02488_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__and2_2
X_19488_ net5754 _03266_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18439_ net7790 _02465_ _02070_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21450_ clknet_leaf_46_i_clk net3856 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ net3608 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21381_ clknet_leaf_58_i_clk _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20263_ net4850 net4839 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__or2_1
X_22002_ net227 net2417 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
Xhold3101 _08288_ vssd1 vssd1 vccd1 vccd1 net3625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3112 rbzero.pov.ready_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net3636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20194_ net1278 _03718_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or2_1
Xhold3123 _03907_ vssd1 vssd1 vccd1 vccd1 net3647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3134 _01000_ vssd1 vssd1 vccd1 vccd1 net3658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2400 _00973_ vssd1 vssd1 vccd1 vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3145 rbzero.pov.spi_buffer\[66\] vssd1 vssd1 vccd1 vccd1 net3669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3156 _03931_ vssd1 vssd1 vccd1 vccd1 net3680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2411 net7904 vssd1 vssd1 vccd1 vccd1 net2935 sky130_fd_sc_hd__buf_2
Xhold2422 _03495_ vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3167 net3779 vssd1 vssd1 vccd1 vccd1 net3691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3178 _03648_ vssd1 vssd1 vccd1 vccd1 net3702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2433 _03547_ vssd1 vssd1 vccd1 vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2444 net4704 vssd1 vssd1 vccd1 vccd1 net2968 sky130_fd_sc_hd__buf_1
Xhold3189 rbzero.pov.ready_buffer\[46\] vssd1 vssd1 vccd1 vccd1 net3713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1710 net2001 vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2455 _02989_ vssd1 vssd1 vccd1 vccd1 net2979 sky130_fd_sc_hd__clkbuf_2
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1721 _01329_ vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2466 rbzero.pov.ready_buffer\[48\] vssd1 vssd1 vccd1 vccd1 net2990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2477 _03500_ vssd1 vssd1 vccd1 vccd1 net3001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1732 net6179 vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1743 _01374_ vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03781_ clknet_0__03781_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03781_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2488 _03376_ vssd1 vssd1 vccd1 vccd1 net3012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1754 _04568_ vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2499 _00639_ vssd1 vssd1 vccd1 vccd1 net3023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1765 net1967 vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1776 _01564_ vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1787 net7102 vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1798 net7041 vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20359__89 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__inv_2
XFILLER_0_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ net6491 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ clknet_leaf_17_i_clk net1914 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _05616_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
X_21648_ clknet_leaf_33_i_clk net1737 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ net6335 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12381_ _05546_ _05547_ _05248_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__mux2_1
XANTENNA_80 _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21579_ clknet_leaf_2_i_clk net5009 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_91 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14120_ _06889_ _06931_ _06846_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__a21oi_1
X_11332_ _04403_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__clkbuf_4
X_14051_ _06861_ _06885_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or2_1
X_11263_ net2882 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5070 net1308 vssd1 vssd1 vccd1 vccd1 net5594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _06140_ _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__and2_1
Xhold5081 net1255 vssd1 vssd1 vccd1 vccd1 net5605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11194_ net5904 net6750 _04470_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__mux2_1
Xhold5092 net1378 vssd1 vssd1 vccd1 vccd1 net5616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4380 rbzero.wall_tracer.rayAddendY\[-7\] vssd1 vssd1 vccd1 vccd1 net4904 sky130_fd_sc_hd__dlygate4sd3_1
X_17810_ _01859_ _01860_ _06205_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o21ai_1
Xhold4391 _06348_ vssd1 vssd1 vccd1 vccd1 net4915 sky130_fd_sc_hd__dlygate4sd3_1
X_18790_ _02779_ _02782_ _08246_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17741_ _01789_ _01790_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__and2_1
Xhold3690 net4222 vssd1 vssd1 vccd1 vccd1 net4214 sky130_fd_sc_hd__dlygate4sd3_1
X_14953_ _08006_ _07990_ _07994_ _08050_ vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__a31o_1
X_13904_ _07029_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__and2_4
X_17672_ _01698_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__xnor2_1
X_14884_ _07991_ _08007_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16623_ _09583_ _09591_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__or2b_1
X_19411_ net1744 _03212_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _06965_ _06979_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap82 _06481_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
X_16554_ _09624_ _09625_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__and2b_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19342_ net1868 _03173_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__or2_1
X_13766_ net79 _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ net2358 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15505_ net3114 _08299_ _06210_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19273_ _08274_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__buf_4
X_12717_ _05876_ _05877_ net13 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__mux2_1
X_16485_ _09542_ _09556_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ _06584_ _06586_ _06722_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18224_ _02166_ _02169_ _02252_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a31o_1
X_15436_ _08461_ _08510_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__xnor2_2
X_12648_ net44 _05785_ _05795_ _05808_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a311o_1
XFILLER_0_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ _02086_ _02110_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15367_ _08381_ _08441_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__nor2_1
X_12579_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _05476_ vssd1 vssd1 vccd1 vccd1 _05744_
+ sky130_fd_sc_hd__mux2_1
X_20967__376 clknet_1_0__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__inv_2
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ _09833_ _09836_ _09834_ vssd1 vssd1 vccd1 vccd1 _10108_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14318_ net3246 _07467_ _07468_ net586 vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ _01675_ _09310_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__or3_1
X_20666__104 clknet_1_1__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__inv_2
Xhold306 _01402_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ net3172 _06209_ _08372_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold317 net5215 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold328 net4737 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ _10042_ _10043_ vssd1 vssd1 vccd1 vccd1 _10044_ sky130_fd_sc_hd__or2b_1
Xhold339 net4904 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03775_ _03775_ vssd1 vssd1 vccd1 vccd1 clknet_0__03775_ sky130_fd_sc_hd__clkbuf_16
X_14249_ _07399_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _09947_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__xnor2_1
Xhold1006 net5722 vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994__20 clknet_1_0__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
Xhold1017 net6525 vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1028 net6579 vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ _01934_ _01910_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__or2b_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1039 net594 vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19609_ net614 _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21502_ clknet_leaf_14_i_clk net1186 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_22482_ clknet_leaf_67_i_clk net1049 vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21433_ clknet_leaf_82_i_clk net3459 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21364_ clknet_leaf_54_i_clk _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21295_ clknet_leaf_27_i_clk net3512 vssd1 vssd1 vccd1 vccd1 rbzero.wall_hot\[1\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold840 net4700 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold851 net5204 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold862 net6468 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 net6492 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20246_ net5665 _03743_ _03750_ _03748_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__o211a_1
Xhold884 net4206 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 _01139_ vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ net5544 _03704_ _03711_ _03709_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__o211a_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2230 _04239_ vssd1 vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 net7132 vssd1 vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2252 net4648 vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__buf_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2263 net5745 vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__buf_1
Xhold2274 _01287_ vssd1 vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2285 net7275 vssd1 vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1540 net6699 vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1551 _01146_ vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2296 net2574 vssd1 vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1562 net6881 vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _04161_ _04608_ net3992 vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_192_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1573 net5878 vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1584 net6825 vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1595 net2196 vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
X_10901_ net6904 net7157 _04321_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_108 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_108/HI zeros[0] sky130_fd_sc_hd__conb_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_119 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_119/HI zeros[11]
+ sky130_fd_sc_hd__conb_1
X_11881_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__clkbuf_8
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _06691_ _06769_ _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ net6403 net1777 _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _06663_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__nand2_1
X_10763_ net7062 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _05229_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or2_1
X_16270_ _09333_ _09343_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13482_ _06631_ _06632_ _06629_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__and3_1
X_10694_ net6642 net6942 _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15221_ _08295_ vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__buf_4
X_12433_ _05000_ _05595_ _05599_ _04978_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ net4370 _08086_ _08249_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__mux2_1
X_12364_ reg_rgb\[14\] _05531_ _05204_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14103_ _07154_ _07187_ _07251_ _07253_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a22o_4
X_11315_ net1816 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19960_ _03569_ net3082 _03571_ _04827_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15083_ _08190_ _08205_ net3207 _01622_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12295_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _05262_ vssd1 vssd1 vccd1 vccd1 _05463_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ _07183_ _07184_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__and2b_1
X_18911_ _02863_ net3700 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nand2_1
X_11246_ net2167 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19891_ _04597_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18842_ _02830_ _02831_ rbzero.wall_tracer.rayAddendY\[1\] _09932_ vssd1 vssd1 vccd1
+ vccd1 _02832_ sky130_fd_sc_hd__a2bb2o_1
X_11177_ _04332_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_175_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15985_ _09047_ _09053_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__nor2_1
X_18773_ _05393_ net4438 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17724_ _09447_ _09784_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__nor2_1
X_14936_ _08020_ _08082_ _08069_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__mux2_1
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__04012_ clknet_0__04012_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04012_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17655_ _10541_ _01700_ _01705_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__nand3_1
X_14867_ _07881_ _07961_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__nor2_1
X_16606_ _09091_ _08795_ _09676_ vssd1 vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__or3_1
X_13818_ _06881_ _06953_ _06935_ _06932_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__a31o_1
XFILLER_0_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17586_ _10485_ _10500_ _10498_ vssd1 vssd1 vccd1 vccd1 _10584_ sky130_fd_sc_hd__a21o_1
X_14798_ _07943_ _07944_ _07946_ _07935_ _07948_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__o221a_1
XFILLER_0_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ net3722 _09304_ _09486_ _09608_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19325_ net5275 _03159_ _03170_ _03168_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__o211a_1
X_13749_ _06897_ _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16468_ _08310_ _09537_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__or2_1
X_19256_ net606 _03120_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__05994_ _05994_ vssd1 vssd1 vccd1 vccd1 clknet_0__05994_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7208 net4338 vssd1 vssd1 vccd1 vccd1 net7732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7219 rbzero.wall_tracer.stepDistY\[2\] vssd1 vssd1 vccd1 vccd1 net7743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15419_ net6259 _08299_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__nand2_1
X_18207_ _02252_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__or2_1
X_19187_ net1531 _03079_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__or2_1
X_16399_ _09466_ _09471_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6507 rbzero.tex_g0\[27\] vssd1 vssd1 vccd1 vccd1 net7031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6518 net2322 vssd1 vssd1 vccd1 vccd1 net7042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6529 rbzero.tex_b1\[30\] vssd1 vssd1 vccd1 vccd1 net7053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18138_ _08705_ _09602_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__nor2_1
Xhold5806 net4013 vssd1 vssd1 vccd1 vccd1 net6330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5817 net1047 vssd1 vssd1 vccd1 vccd1 net6341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 net6327 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5828 _04576_ vssd1 vssd1 vccd1 vccd1 net6352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5839 net1172 vssd1 vssd1 vccd1 vccd1 net6363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 net5700 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18069_ _08643_ _09420_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__or2_1
Xhold125 net5839 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold136 net4955 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 rbzero.wall_tracer.visualWallDist\[6\] vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold158 rbzero.wall_tracer.visualWallDist\[8\] vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_1
X_20100_ net4865 net4797 _03663_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__o21a_1
X_21080_ _04018_ _04072_ _04074_ _04017_ net4503 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a32o_1
Xhold169 net4147 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20031_ _03616_ net3877 vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__or2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720__153 clknet_1_0__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__inv_2
X_21982_ net207 net2392 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20337__70 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
XFILLER_0_14_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22465_ clknet_leaf_69_i_clk net659 vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20352__84 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__inv_2
X_21416_ clknet_leaf_78_i_clk net4756 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22396_ net148 net1855 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
X_21347_ clknet_leaf_39_i_clk net4162 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ net7083 net6844 _04426_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
X_12080_ rbzero.tex_r1\[45\] rbzero.tex_r1\[44\] _05230_ vssd1 vssd1 vccd1 vccd1 _05249_
+ sky130_fd_sc_hd__mux2_1
X_21278_ clknet_leaf_59_i_clk _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold670 net5535 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 net5552 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 net4209 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net2440 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__clkbuf_1
X_20229_ net5219 _03730_ _03740_ _03735_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__o211a_1
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 net6937 vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 _00891_ vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2082 net6811 vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
X_15770_ _08812_ _08815_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__xor2_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2093 _04451_ vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _06135_ _06137_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__nand2_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1370 net6821 vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _07854_ _07870_ _07871_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__a21oi_1
Xhold1381 _00926_ vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
X_20695__130 clknet_1_1__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__inv_2
X_11933_ _05098_ _05102_ net4239 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a21oi_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 net5803 vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _10437_ _10438_ vssd1 vssd1 vccd1 vccd1 _10440_ sky130_fd_sc_hd__nand2_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _07799_ _07801_ _07802_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__nand3_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11864_ _04999_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _06608_ _06687_ _06753_ _06676_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__a211o_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _10355_ _10370_ vssd1 vssd1 vccd1 vccd1 _10371_ sky130_fd_sc_hd__xnor2_1
X_10815_ net7149 net2668 _04277_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _07718_ _07733_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11795_ _04964_ _04918_ _04920_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16322_ _09393_ _09394_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19110_ net5973 _03037_ _03045_ _03022_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__o211a_1
X_13534_ _06613_ _06596_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__or3_4
X_10746_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19041_ net3941 _02990_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__or2_1
X_16253_ _08409_ _09091_ _09187_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _06423_ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_168_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10677_ net2635 net6760 _04203_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__mux2_1
X_15204_ net4079 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
X_12416_ _05581_ _05582_ _05235_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ _08799_ _09258_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ _06545_ _06546_ _06540_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_140_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15135_ net4779 _08223_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__or2_1
X_12347_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _05493_ vssd1 vssd1 vccd1 vccd1 _05515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19943_ net4675 _03553_ _03485_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__o21ai_1
X_15066_ _04624_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__clkbuf_8
X_12278_ reg_rgb\[7\] _05446_ _05204_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__mux2_4
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14017_ _07123_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__xnor2_1
X_11229_ net5867 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19874_ net3821 _08479_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a21o_1
X_18825_ _02810_ _02815_ _04623_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20778__205 clknet_1_0__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__inv_2
X_20661__99 clknet_1_0__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__inv_2
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18756_ _05393_ net738 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__nand2_1
X_15968_ _09017_ _09018_ _09024_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__a21oi_1
X_17707_ _01670_ _10584_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__or2b_1
XFILLER_0_175_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14919_ net7891 _08063_ _08064_ _08066_ net7566 vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__a311o_1
X_15899_ _08968_ _08972_ _08973_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__a21bo_1
X_18687_ _02646_ _05401_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__or2_1
XFILLER_0_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _01684_ _09484_ _10515_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__o31a_1
XFILLER_0_188_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _10566_ _10567_ vssd1 vssd1 vccd1 vccd1 _10568_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19308_ net5259 _03159_ _03161_ _03155_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20580_ net3681 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_1
Xhold7005 rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 net7529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7016 net4510 vssd1 vssd1 vccd1 vccd1 net7540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7027 rbzero.wall_tracer.trackDistX\[2\] vssd1 vssd1 vccd1 vccd1 net7551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19239_ net809 _03120_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__or2_1
Xhold7038 rbzero.wall_tracer.trackDistX\[-9\] vssd1 vssd1 vccd1 vccd1 net7562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6304 net1818 vssd1 vssd1 vccd1 vccd1 net6828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7049 rbzero.traced_texa\[8\] vssd1 vssd1 vccd1 vccd1 net7573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6315 _04560_ vssd1 vssd1 vccd1 vccd1 net6839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22250_ net382 net1823 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold6326 net1697 vssd1 vssd1 vccd1 vccd1 net6850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6337 rbzero.tex_b1\[13\] vssd1 vssd1 vccd1 vccd1 net6861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6348 net2027 vssd1 vssd1 vccd1 vccd1 net6872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5603 net3003 vssd1 vssd1 vccd1 vccd1 net6127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6359 rbzero.tex_b1\[59\] vssd1 vssd1 vccd1 vccd1 net6883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5614 _08202_ vssd1 vssd1 vccd1 vccd1 net6138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21201_ _02758_ net4801 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__xnor2_1
Xhold5625 _08234_ vssd1 vssd1 vccd1 vccd1 net6149 sky130_fd_sc_hd__dlygate4sd3_1
X_22181_ net313 net1919 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4902 net999 vssd1 vssd1 vccd1 vccd1 net5426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5647 rbzero.spi_registers.spi_buffer\[8\] vssd1 vssd1 vccd1 vccd1 net6171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5658 net4090 vssd1 vssd1 vccd1 vccd1 net6182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4913 net1044 vssd1 vssd1 vccd1 vccd1 net5437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5669 net2958 vssd1 vssd1 vccd1 vccd1 net6193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4924 _00679_ vssd1 vssd1 vccd1 vccd1 net5448 sky130_fd_sc_hd__dlygate4sd3_1
X_21132_ _04113_ _04114_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nor2_1
Xhold4935 net1058 vssd1 vssd1 vccd1 vccd1 net5459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4946 rbzero.traced_texa\[-6\] vssd1 vssd1 vccd1 vccd1 net5470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4957 net1335 vssd1 vssd1 vccd1 vccd1 net5481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4968 _00389_ vssd1 vssd1 vccd1 vccd1 net5492 sky130_fd_sc_hd__dlygate4sd3_1
X_21063_ net4130 net4395 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nand2_1
Xhold4979 rbzero.spi_registers.texadd2\[17\] vssd1 vssd1 vccd1 vccd1 net5503 sky130_fd_sc_hd__dlygate4sd3_1
X_20014_ net3657 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ net190 net2806 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21896_ clknet_leaf_95_i_clk net1471 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ net4004 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__buf_4
X_11580_ _04724_ _04675_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and3_1
XFILLER_0_193_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13250_ net4822 _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22448_ clknet_leaf_66_i_clk _01617_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _05353_ _05366_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _06325_ _06336_ _06321_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__a21oi_1
X_22379_ net511 net2857 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6882 _09296_ vssd1 vssd1 vccd1 vccd1 net7406 sky130_fd_sc_hd__dlygate4sd3_1
X_12132_ _04806_ _05192_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20727__159 clknet_1_1__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__inv_2
XFILLER_0_103_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ _05229_ _05231_ net80 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o21a_1
X_16940_ net4874 net3265 _09294_ vssd1 vssd1 vccd1 vccd1 _09958_ sky130_fd_sc_hd__o21a_1
X_11014_ net5833 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16871_ _04818_ net3535 _09929_ vssd1 vssd1 vccd1 vccd1 _09930_ sky130_fd_sc_hd__or3_4
XFILLER_0_99_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18610_ net87 _02613_ _02619_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15822_ _08857_ _08859_ _08858_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__a21o_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ net5072 _03325_ _03329_ _03330_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__o211a_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _08524_ _08511_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__xnor2_2
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18541_ net2919 net6241 _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _06112_ _06118_ _06120_ _06109_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__o211a_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _05077_ vssd1 vssd1 vccd1 vccd1 _05086_
+ sky130_fd_sc_hd__mux2_1
X_14704_ _07828_ _07820_ _07827_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__nand3_1
X_15684_ _08753_ _08758_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ net3074 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ net39 _06051_ _06052_ net36 vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and4b_1
XFILLER_0_185_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _10420_ _10421_ _10302_ vssd1 vssd1 vccd1 vccd1 _10423_ sky130_fd_sc_hd__a21o_1
X_14635_ _07766_ _07784_ _07785_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__a21oi_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11847_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _04994_ vssd1 vssd1 vccd1 vccd1 _05017_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _08724_ net7378 vssd1 vssd1 vccd1 vccd1 _10354_ sky130_fd_sc_hd__and2_1
X_14566_ _07714_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__nor2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ net1072 net1456 net1166 net700 vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03992_ clknet_0__03992_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03992_
+ sky130_fd_sc_hd__clkbuf_16
X_20316__51 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
X_16305_ _09362_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__xnor2_2
X_13517_ net84 _06588_ _06597_ _06610_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__and4_4
X_10729_ net2382 net6898 _04225_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__mux2_1
X_17285_ _10284_ _10285_ vssd1 vssd1 vccd1 vccd1 _10286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14497_ _07587_ _07591_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__xnor2_1
X_16236_ net6150 _08314_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19024_ net6307 _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__or2_1
X_13448_ _06515_ _06503_ _06560_ _06593_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_113_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20331__65 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
X_16167_ _09206_ _09241_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ _06527_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__xor2_2
Xhold4209 net7583 vssd1 vssd1 vccd1 vccd1 net4733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15118_ net4403 net4458 _08219_ vssd1 vssd1 vccd1 vccd1 _08231_ sky130_fd_sc_hd__mux2_1
X_16098_ _08997_ _09172_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__xnor2_1
Xhold3508 gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 net4032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3519 net4005 vssd1 vssd1 vccd1 vccd1 net4043 sky130_fd_sc_hd__buf_4
XFILLER_0_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15049_ net4431 _08181_ _08138_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__mux2_1
X_19926_ net6127 _03530_ net2890 _03496_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__o211a_1
Xhold2807 _01032_ vssd1 vssd1 vccd1 vccd1 net3331 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_74_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2818 net1343 vssd1 vssd1 vccd1 vccd1 net3342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 _03828_ vssd1 vssd1 vccd1 vccd1 net3353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19857_ _03479_ net6009 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__or2_1
X_18808_ _02792_ _02797_ net7575 net4626 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19788_ net1989 _03443_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
XFILLER_0_207_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_89_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18739_ net3805 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21750_ clknet_leaf_102_i_clk net2022 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21681_ clknet_leaf_35_i_clk net5285 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdxw\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04009_ _04009_ vssd1 vssd1 vccd1 vccd1 clknet_0__04009_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20832__254 clknet_1_1__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__inv_2
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20632_ _05816_ _03032_ net4060 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20563_ _03902_ net3706 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6101 rbzero.tex_r1\[35\] vssd1 vssd1 vccd1 vccd1 net6625 sky130_fd_sc_hd__dlygate4sd3_1
X_22302_ net434 net2065 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold6112 net1706 vssd1 vssd1 vccd1 vccd1 net6636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold6123 _04368_ vssd1 vssd1 vccd1 vccd1 net6647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6134 net1716 vssd1 vssd1 vccd1 vccd1 net6658 sky130_fd_sc_hd__dlygate4sd3_1
X_20494_ net3339 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
Xhold5400 net2650 vssd1 vssd1 vccd1 vccd1 net5924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6145 rbzero.tex_g0\[17\] vssd1 vssd1 vccd1 vccd1 net6669 sky130_fd_sc_hd__dlygate4sd3_1
X_22233_ net365 net830 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold6156 net1766 vssd1 vssd1 vccd1 vccd1 net6680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5411 net2191 vssd1 vssd1 vccd1 vccd1 net5935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6167 rbzero.tex_b0\[61\] vssd1 vssd1 vccd1 vccd1 net6691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5422 rbzero.map_overlay.i_mapdy\[3\] vssd1 vssd1 vccd1 vccd1 net5946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6178 net1973 vssd1 vssd1 vccd1 vccd1 net6702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5433 net4001 vssd1 vssd1 vccd1 vccd1 net5957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6189 rbzero.tex_r0\[45\] vssd1 vssd1 vccd1 vccd1 net6713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5444 rbzero.wall_tracer.mapX\[7\] vssd1 vssd1 vccd1 vccd1 net5968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4710 _01069_ vssd1 vssd1 vccd1 vccd1 net5234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5455 _00674_ vssd1 vssd1 vccd1 vccd1 net5979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4721 net844 vssd1 vssd1 vccd1 vccd1 net5245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5466 _04327_ vssd1 vssd1 vccd1 vccd1 net5990 sky130_fd_sc_hd__dlygate4sd3_1
X_22164_ net296 net1612 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5477 rbzero.map_overlay.i_mapdy\[1\] vssd1 vssd1 vccd1 vccd1 net6001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4732 _00820_ vssd1 vssd1 vccd1 vccd1 net5256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5488 net2936 vssd1 vssd1 vccd1 vccd1 net6012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4743 net971 vssd1 vssd1 vccd1 vccd1 net5267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4754 rbzero.spi_registers.buf_mapdyw\[1\] vssd1 vssd1 vccd1 vccd1 net5278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5499 net2993 vssd1 vssd1 vccd1 vccd1 net6023 sky130_fd_sc_hd__dlygate4sd3_1
X_21115_ net4160 net4653 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__nor2_1
Xhold4765 net1003 vssd1 vssd1 vccd1 vccd1 net5289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4776 net957 vssd1 vssd1 vccd1 vccd1 net5300 sky130_fd_sc_hd__dlygate4sd3_1
X_22095_ clknet_leaf_6_i_clk _01264_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4787 _00505_ vssd1 vssd1 vccd1 vccd1 net5311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4798 net904 vssd1 vssd1 vccd1 vccd1 net5322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21046_ _04044_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _05207_ _05904_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a21oi_1
X_21948_ net173 net2217 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ _04863_ _04599_ net4010 net2917 _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ net14 net15 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21879_ clknet_leaf_99_i_clk net1231 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _07568_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__xor2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ net4972 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14351_ _07495_ _07501_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ _04691_ _04694_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17070_ _10073_ net3417 net4903 vssd1 vssd1 vccd1 vccd1 _10074_ sky130_fd_sc_hd__mux2_1
X_14282_ _07386_ _07408_ _07431_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__nand3_1
X_11494_ _04658_ _04663_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21o_1
X_16021_ _08626_ vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7380 rbzero.debug_overlay.playerX\[-5\] vssd1 vssd1 vccd1 vccd1 net7904 sky130_fd_sc_hd__dlygate4sd3_1
X_13233_ net4917 vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__inv_2
Xhold7391 rbzero.wall_tracer.stepDistY\[5\] vssd1 vssd1 vccd1 vccd1 net7915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6690 rbzero.tex_b1\[48\] vssd1 vssd1 vccd1 vccd1 net7214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13164_ net3432 vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__inv_2
X_12115_ rbzero.tex_r1\[27\] rbzero.tex_r1\[26\] _05230_ vssd1 vssd1 vccd1 vccd1 _05284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17972_ _09582_ _01711_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__nor2_1
X_13095_ _06243_ _06247_ _06249_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__or4b_1
X_19711_ net6662 _03395_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__or2_1
X_12046_ rbzero.tex_r1\[53\] rbzero.tex_r1\[52\] _05071_ vssd1 vssd1 vccd1 vccd1 _05215_
+ sky130_fd_sc_hd__mux2_1
X_16923_ _08246_ _09930_ vssd1 vssd1 vccd1 vccd1 _09943_ sky130_fd_sc_hd__or2_4
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19642_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__clkbuf_4
X_16854_ _04727_ _04725_ _09920_ vssd1 vssd1 vccd1 vccd1 _09921_ sky130_fd_sc_hd__o21ai_1
X_15805_ _08865_ _08867_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19573_ _02996_ _03304_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__or2_1
X_16785_ _08587_ _09483_ vssd1 vssd1 vccd1 vccd1 _09855_ sky130_fd_sc_hd__or2_2
X_13997_ net3163 _07146_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__or2b_1
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18524_ net3838 net1076 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__nand2_1
X_15736_ _08556_ net7444 vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__nor2_2
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ _06098_ _06101_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18455_ _02254_ _02255_ _02479_ _02261_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a22o_1
X_15667_ _08691_ _08723_ _08741_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__a21o_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ net31 net30 vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2b_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17406_ _09064_ vssd1 vssd1 vccd1 vccd1 _10406_ sky130_fd_sc_hd__buf_2
XFILLER_0_158_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _07727_ _07729_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15598_ _08671_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__xor2_1
X_18386_ net4536 net4372 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17337_ _10209_ _10335_ _10333_ _10334_ vssd1 vssd1 vccd1 vccd1 _10337_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14549_ _07697_ _07698_ _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__nand3_1
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17268_ _10267_ _10268_ vssd1 vssd1 vccd1 vccd1 _10269_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19007_ net7357 _02967_ net3905 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__and3b_1
XFILLER_0_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ net7405 vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17199_ _10087_ _10200_ vssd1 vssd1 vccd1 vccd1 _10201_ sky130_fd_sc_hd__xor2_4
XFILLER_0_109_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4006 net3420 vssd1 vssd1 vccd1 vccd1 net4530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4017 rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 net4541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4028 _02764_ vssd1 vssd1 vccd1 vccd1 net4552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4039 _00994_ vssd1 vssd1 vccd1 vccd1 net4563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3316 _03627_ vssd1 vssd1 vccd1 vccd1 net3840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3327 net4688 vssd1 vssd1 vccd1 vccd1 net3851 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3338 _02832_ vssd1 vssd1 vccd1 vccd1 net3862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3349 net7349 vssd1 vssd1 vccd1 vccd1 net3873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2604 rbzero.color_floor\[5\] vssd1 vssd1 vccd1 vccd1 net3128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 rbzero.pov.ready_buffer\[39\] vssd1 vssd1 vccd1 vccd1 net3139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2626 net7338 vssd1 vssd1 vccd1 vccd1 net3150 sky130_fd_sc_hd__clkbuf_2
X_19909_ net3365 _03477_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a211o_1
XFILLER_0_209_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2637 net4404 vssd1 vssd1 vccd1 vccd1 net3161 sky130_fd_sc_hd__buf_1
Xhold1903 rbzero.tex_r1\[59\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 net4715 vssd1 vssd1 vccd1 vccd1 net3172 sky130_fd_sc_hd__clkbuf_2
Xhold1914 _01271_ vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2659 _00804_ vssd1 vssd1 vccd1 vccd1 net3183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1925 net2243 vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1936 _01470_ vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1947 _01570_ vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1958 net6807 vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1969 net5980 vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21802_ clknet_leaf_89_i_clk net2838 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21733_ clknet_leaf_22_i_clk net1911 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21664_ clknet_leaf_35_i_clk net5180 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20615_ net4016 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21595_ clknet_leaf_21_i_clk net4270 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20546_ net3081 net3568 _03889_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20477_ _03858_ net3413 vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__and2_1
Xhold5230 net1141 vssd1 vssd1 vccd1 vccd1 net5754 sky130_fd_sc_hd__dlygate4sd3_1
X_20310__46 clknet_1_0__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
X_22216_ net348 net1799 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
Xhold5241 net1614 vssd1 vssd1 vccd1 vccd1 net5765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5252 _04314_ vssd1 vssd1 vccd1 vccd1 net5776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5263 rbzero.spi_registers.texadd0\[1\] vssd1 vssd1 vccd1 vccd1 net5787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5274 rbzero.tex_r1\[38\] vssd1 vssd1 vccd1 vccd1 net5798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4540 rbzero.spi_registers.buf_mapdy\[0\] vssd1 vssd1 vccd1 vccd1 net5064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5285 _00658_ vssd1 vssd1 vccd1 vccd1 net5809 sky130_fd_sc_hd__dlygate4sd3_1
X_22147_ net279 net2324 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
Xhold5296 rbzero.tex_r1\[40\] vssd1 vssd1 vccd1 vccd1 net5820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4551 rbzero.spi_registers.texadd0\[21\] vssd1 vssd1 vccd1 vccd1 net5075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4562 rbzero.spi_registers.buf_texadd0\[0\] vssd1 vssd1 vccd1 vccd1 net5086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4573 net834 vssd1 vssd1 vccd1 vccd1 net5097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4584 net812 vssd1 vssd1 vccd1 vccd1 net5108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4595 net827 vssd1 vssd1 vccd1 vccd1 net5119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3850 net3115 vssd1 vssd1 vccd1 vccd1 net4374 sky130_fd_sc_hd__buf_1
Xhold3861 net7787 vssd1 vssd1 vccd1 vccd1 net4385 sky130_fd_sc_hd__dlygate4sd3_1
X_22078_ clknet_leaf_13_i_clk net3313 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3872 _01598_ vssd1 vssd1 vccd1 vccd1 net4396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3883 _03598_ vssd1 vssd1 vccd1 vccd1 net4407 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03995_ clknet_0__03995_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03995_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21029_ _04028_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13920_ _07024_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ _06880_ _06889_ _07000_ _07001_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_97_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ net53 _05946_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__nand2_1
X_16570_ _09641_ vssd1 vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__inv_2
X_13782_ _06882_ _06883_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__and2_4
X_10994_ net7022 net7286 _04366_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__nor2_1
X_15521_ _08320_ _08593_ _08595_ _08379_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__a211o_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15452_ _08332_ _08526_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__or2_1
X_18240_ _08705_ _09732_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__nor2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ net3965 _05795_ _05799_ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a22o_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _07551_ _07552_ _07553_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__and3_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ _04714_ _04781_ _04783_ _04721_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a221o_1
XFILLER_0_182_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15383_ _08448_ _08450_ _08457_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__nand3_1
X_18171_ _01802_ _09602_ _02094_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__or3_1
X_12595_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04988_ vssd1 vssd1 vccd1 vccd1 _05760_
+ sky130_fd_sc_hd__mux2_1
X_17122_ _10122_ _10123_ vssd1 vssd1 vccd1 vccd1 _10124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _07478_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11546_ net4891 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17053_ _10050_ _10051_ _10052_ vssd1 vssd1 vccd1 vccd1 _10058_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ _07414_ _07415_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ rbzero.spi_registers.texadd3\[11\] rbzero.spi_registers.texadd1\[11\] rbzero.spi_registers.texadd0\[11\]
+ rbzero.spi_registers.texadd2\[11\] _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04649_
+ sky130_fd_sc_hd__mux4_1
X_16004_ _09036_ _09037_ _09039_ _09077_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__a22o_1
X_13216_ _06217_ _06216_ net3984 net4874 vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__or4_1
X_14196_ _07297_ _07296_ _07294_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ net3555 _06299_ net3472 _06301_ _06302_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a221oi_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20861__280 clknet_1_0__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__inv_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17955_ _02002_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__and2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ net3881 _06186_ _06196_ net3279 _06233_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12029_ net4041 net4004 net3992 vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16906_ net4152 _09939_ _09940_ net645 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
X_17886_ _01826_ _01829_ _01827_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a21bo_1
X_19625_ net4991 net799 _03349_ _03343_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__o211a_1
X_16837_ _09782_ _09906_ vssd1 vssd1 vccd1 vccd1 _09907_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_164_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19556_ net3070 _03305_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__or2_1
X_16768_ _09833_ _09837_ vssd1 vssd1 vccd1 vccd1 _09838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18507_ _02526_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__clkbuf_1
X_15719_ _08312_ _08793_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__or2_1
X_19487_ net1572 _03265_ net2542 _03260_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__o211a_1
X_16699_ net7446 net3028 _08293_ vssd1 vssd1 vccd1 vccd1 _09770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18438_ _02462_ _02463_ _01870_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18369_ _02404_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__clkbuf_1
X_20400_ _03791_ net3607 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21380_ clknet_leaf_64_i_clk _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03989_ _03989_ vssd1 vssd1 vccd1 vccd1 clknet_0__03989_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20944__355 clknet_1_0__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__inv_2
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20262_ net4850 _03756_ _03759_ _03748_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22001_ net226 net1908 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
Xhold3102 _00463_ vssd1 vssd1 vccd1 vccd1 net3626 sky130_fd_sc_hd__dlygate4sd3_1
X_20193_ net5114 _03717_ _03720_ _03709_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__o211a_1
Xhold3113 _03798_ vssd1 vssd1 vccd1 vccd1 net3637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3124 _03908_ vssd1 vssd1 vccd1 vccd1 net3648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3135 net5600 vssd1 vssd1 vccd1 vccd1 net3659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2401 net6016 vssd1 vssd1 vccd1 vccd1 net2925 sky130_fd_sc_hd__buf_1
Xhold3146 net1241 vssd1 vssd1 vccd1 vccd1 net3670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2412 net6011 vssd1 vssd1 vccd1 vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3157 _03932_ vssd1 vssd1 vccd1 vccd1 net3681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2423 net4301 vssd1 vssd1 vccd1 vccd1 net2947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3168 _08242_ vssd1 vssd1 vccd1 vccd1 net3692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3179 _01025_ vssd1 vssd1 vccd1 vccd1 net3703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2434 net6192 vssd1 vssd1 vccd1 vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1700 net6781 vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2445 net4706 vssd1 vssd1 vccd1 vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1711 _04352_ vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2456 _03024_ vssd1 vssd1 vccd1 vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1722 net7074 vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2467 _03543_ vssd1 vssd1 vccd1 vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 net6200 vssd1 vssd1 vccd1 vccd1 net3002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _03372_ vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1744 net6951 vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03780_ clknet_0__03780_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03780_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2489 _00887_ vssd1 vssd1 vccd1 vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1755 _01136_ vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1766 _04535_ vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1777 net6997 vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1788 _01434_ vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1799 _04473_ vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21716_ clknet_leaf_26_i_clk net2258 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21647_ clknet_leaf_34_i_clk net2555 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11400_ net6333 net1620 _04584_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12380_ rbzero.tex_g1\[63\] rbzero.tex_g1\[62\] _05483_ vssd1 vssd1 vccd1 vccd1 _05547_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_70 rbzero.wall_tracer.visualWallDist\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21578_ clknet_leaf_2_i_clk net5316 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_81 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11331_ net2531 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_92 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20529_ net3437 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
X_14050_ _07199_ _07200_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or2_1
X_11262_ net7187 net7298 _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5060 rbzero.pov.spi_buffer\[15\] vssd1 vssd1 vccd1 vccd1 net5584 sky130_fd_sc_hd__dlygate4sd3_1
X_13001_ _06124_ _06117_ _06121_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__nand3_1
XFILLER_0_123_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5071 _00755_ vssd1 vssd1 vccd1 vccd1 net5595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5082 _00785_ vssd1 vssd1 vccd1 vccd1 net5606 sky130_fd_sc_hd__dlygate4sd3_1
X_11193_ net6427 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5093 rbzero.pov.spi_buffer\[28\] vssd1 vssd1 vccd1 vccd1 net5617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4370 _00972_ vssd1 vssd1 vccd1 vccd1 net4894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4381 net863 vssd1 vssd1 vccd1 vccd1 net4905 sky130_fd_sc_hd__buf_1
XFILLER_0_98_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4392 _06359_ vssd1 vssd1 vccd1 vccd1 net4916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3680 net891 vssd1 vssd1 vccd1 vccd1 net4204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17740_ _01789_ _01790_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nor2_1
Xhold3691 _03166_ vssd1 vssd1 vccd1 vccd1 net4215 sky130_fd_sc_hd__dlygate4sd3_1
X_14952_ _08097_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__clkbuf_1
X_13903_ _07026_ _07028_ _07027_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__a21bo_1
Xhold2990 net1360 vssd1 vssd1 vccd1 vccd1 net3514 sky130_fd_sc_hd__clkdlybuf4s25_1
X_17671_ _01721_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nor2_1
X_14883_ _06664_ _08030_ _08032_ net7457 vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__a31o_1
X_19410_ net5690 _03211_ _03218_ _03207_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__o211a_1
X_16622_ _09585_ _09590_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ _06981_ _06983_ _06984_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19341_ net5642 _03172_ _03179_ _03168_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__o211a_1
X_16553_ _09621_ _09623_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__nand2_1
X_13765_ net561 _06796_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__xnor2_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap83 _04816_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
X_10977_ net6415 net7052 _04355_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15504_ _08320_ _08576_ _08578_ _08305_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__a211o_2
X_19272_ net5034 _03133_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__or2_1
X_12716_ _04159_ _04718_ _04726_ _04777_ net10 net11 vssd1 vssd1 vccd1 vccd1 _05877_
+ sky130_fd_sc_hd__mux4_1
X_16484_ _09553_ _09555_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13696_ _06660_ _06751_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__nor2_1
X_18223_ _02164_ _02268_ _02251_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a21oi_1
X_15435_ _08463_ _08509_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__xor2_2
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12647_ net4043 _05785_ _05799_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__and3_1
XFILLER_0_210_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18154_ _02178_ _02200_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__xnor2_1
X_15366_ _08439_ _08440_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__nand2_1
X_12578_ _05062_ _05738_ _05740_ _05742_ _05030_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _09676_ _09815_ _09814_ vssd1 vssd1 vccd1 vccd1 _10107_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14317_ _07311_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__nor2_2
X_11529_ _04699_ _04700_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand2_1
X_18085_ _02131_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__xnor2_1
X_15297_ _08298_ _08370_ _08371_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold307 net5078 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 net5217 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03774_ _03774_ vssd1 vssd1 vccd1 vccd1 clknet_0__03774_ sky130_fd_sc_hd__clkbuf_16
X_17036_ net4560 net4399 vssd1 vssd1 vccd1 vccd1 _10043_ sky130_fd_sc_hd__nand2_1
X_14248_ _07351_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__xnor2_2
Xhold329 net5154 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ _07328_ _07329_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ net4874 _09968_ _09974_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a21oi_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 net6228 vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _01889_ _01904_ _01902_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a21o_1
Xhold1018 _00812_ vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1029 _01497_ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17869_ _01916_ _01917_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or2_1
X_19608_ _03326_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__buf_2
X_20880_ clknet_1_1__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__buf_1
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19539_ _02491_ _02497_ net3076 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21501_ clknet_leaf_14_i_clk net638 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22481_ clknet_leaf_66_i_clk net663 vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21432_ clknet_leaf_80_i_clk net3248 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21363_ clknet_leaf_56_i_clk _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold830 _01502_ vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21294_ clknet_leaf_27_i_clk net3626 vssd1 vssd1 vccd1 vccd1 rbzero.wall_hot\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold841 net4702 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold852 net5206 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold863 net6470 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_20245_ net5623 _03744_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or2_1
Xhold874 net6494 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 net3556 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 net5638 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ net5520 _03705_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__or2_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2220 _04469_ vssd1 vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2231 _01524_ vssd1 vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2242 _04361_ vssd1 vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2253 net4650 vssd1 vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2264 net5747 vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1530 net6711 vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2275 net7269 vssd1 vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2286 _04585_ vssd1 vssd1 vccd1 vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1541 _01471_ vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2297 _04179_ vssd1 vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 net6853 vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 _01536_ vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1574 net5880 vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10900_ net7159 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1585 _01467_ vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1596 net5866 vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
X_11880_ _04971_ _05026_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__nor2_2
Xtop_ew_algofoogle_109 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_109/HI zeros[1] sky130_fd_sc_hd__conb_1
XFILLER_0_212_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10831_ _04243_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13550_ _06692_ _06696_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ net7060 net2756 _04244_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _05262_ vssd1 vssd1 vccd1 vccd1 _05667_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13481_ _06549_ _06553_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__xor2_2
XFILLER_0_109_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10693_ _04169_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ _08294_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__clkbuf_4
X_12432_ _05003_ _05596_ _05598_ _05009_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15151_ _08253_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12363_ _04816_ _05530_ net4044 vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14102_ _07154_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__xor2_2
XFILLER_0_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11314_ net6742 net6399 _04540_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15082_ net3206 _08201_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__or2_1
X_12294_ _05279_ _05458_ _05460_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14033_ net537 _07143_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__xor2_1
X_18910_ _02863_ net3700 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or2_1
X_11245_ net6708 net6926 _04503_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
X_19890_ net3524 _03485_ _03516_ _03517_ _03474_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18841_ _02828_ _02829_ _04624_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a21o_1
X_11176_ net2744 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18772_ _05393_ net4438 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__nand2_1
X_15984_ _09055_ _09058_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17723_ _01772_ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14935_ net7908 _08011_ _08081_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__04011_ clknet_0__04011_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04011_
+ sky130_fd_sc_hd__clkbuf_16
X_17654_ _10541_ _01700_ _01705_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a21o_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ net527 _07965_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__xor2_4
XFILLER_0_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16605_ _08409_ _09250_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__or2_1
X_20973__381 clknet_1_1__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__inv_2
X_13817_ _06897_ _06899_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__a21bo_1
X_17585_ _10581_ _10582_ vssd1 vssd1 vccd1 vccd1 _10583_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14797_ _07938_ _07940_ _07945_ _07947_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19324_ net1768 _03160_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__or2_1
X_16536_ _09606_ _09607_ _08609_ vssd1 vssd1 vccd1 vccd1 _09608_ sky130_fd_sc_hd__o21ai_4
X_13748_ net3370 _06898_ _06885_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19255_ net4248 _03119_ _03130_ _03128_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__o211a_1
X_16467_ _08310_ _09420_ _09538_ _08326_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__o22a_1
X_13679_ _06725_ _06828_ _06829_ _06716_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7209 _09277_ vssd1 vssd1 vccd1 vccd1 net7733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _02166_ _02169_ _02164_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a21bo_1
X_15418_ _08492_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19186_ net2966 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
X_16398_ _09469_ _09470_ vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__xnor2_1
Xhold6508 net2527 vssd1 vssd1 vccd1 vccd1 net7032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6519 rbzero.tex_r1\[42\] vssd1 vssd1 vccd1 vccd1 net7043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _02182_ _02183_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15349_ _08422_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5807 _01257_ vssd1 vssd1 vccd1 vccd1 net6331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5818 rbzero.tex_g1\[8\] vssd1 vssd1 vccd1 vccd1 net6342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5829 net1032 vssd1 vssd1 vccd1 vccd1 net6353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _02527_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold115 net3285 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ _02051_ _02032_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__or2b_1
Xhold126 net4961 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold137 net4957 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net4161 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold159 net4134 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _10026_ _10024_ _10025_ _06205_ vssd1 vssd1 vccd1 vccd1 _10028_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20030_ net3876 net3709 _03594_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21981_ net206 net1826 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22464_ clknet_leaf_57_i_clk _01633_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21415_ clknet_leaf_78_i_clk net3798 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22395_ net147 net2300 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
X_21346_ clknet_leaf_39_i_clk net4145 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21277_ clknet_leaf_59_i_clk _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold660 _01647_ vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 net5537 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 net6432 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net7064 net6543 _04392_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__mux2_1
X_20228_ net5205 _03731_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or2_1
Xhold693 net5791 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ net5500 _03692_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__or2_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2050 net2819 vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2061 _04512_ vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 net7096 vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2083 _01274_ vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _06134_ _06136_ _06130_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2094 _01336_ vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _03402_ vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 _04564_ vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _07855_ _07856_ _07869_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__and3_1
Xhold1382 net6691 vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ net4254 net4280 _04977_ _05099_ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__o41a_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 net6715 vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11863_ _05003_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__or2_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _07755_ _07757_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ net6946 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__clkbuf_1
X_13602_ _06697_ _06698_ _06603_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__a21oi_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17370_ _10368_ _10369_ vssd1 vssd1 vccd1 vccd1 _10370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ net2931 _04963_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__xor2_1
X_14582_ _07719_ _07731_ _07732_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_138_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16321_ _09393_ _09394_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13533_ _06606_ _06627_ _06600_ _06603_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__or4_1
X_10745_ _04241_ _04160_ _04166_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__or3b_4
XFILLER_0_193_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19040_ net6225 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__clkbuf_1
X_16252_ _09214_ _09207_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13464_ _06614_ _06541_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__or2_2
X_10676_ net2344 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12415_ rbzero.tex_g1\[7\] rbzero.tex_g1\[6\] _05457_ vssd1 vssd1 vccd1 vccd1 _05582_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15203_ _08279_ net4078 vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16183_ _09256_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__nor2_1
X_13395_ net6098 _06431_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12346_ _05510_ _05513_ net80 vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15134_ net3691 net3058 _06344_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ net3722 _06386_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__nand2_1
X_19942_ net3286 _03485_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12277_ net4007 vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _07125_ _07124_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__or2b_1
X_11228_ net2197 net5865 _04492_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__mux2_1
X_19873_ _03485_ _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18824_ _02811_ _02814_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__xnor2_1
X_20704__138 clknet_1_1__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__inv_2
X_11159_ net5814 net5848 _04459_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18755_ net4640 net4905 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__nor2_1
X_15967_ _09017_ _09018_ _09024_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_1__f__06092_ clknet_0__06092_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__06092_
+ sky130_fd_sc_hd__clkbuf_16
X_17706_ _10469_ _01735_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14918_ _07995_ _08036_ _08037_ _08065_ net7843 vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__o311a_1
X_18686_ _02686_ _02687_ net4811 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__nand3_2
XFILLER_0_78_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _08970_ _08971_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__nand2_1
X_17637_ _10517_ _10518_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__or2_1
X_14849_ _07995_ _07999_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17568_ _10465_ _10466_ _10565_ vssd1 vssd1 vccd1 vccd1 _10567_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19307_ net1647 _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16519_ _09585_ _09590_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _10496_ _10497_ vssd1 vssd1 vccd1 vccd1 _10498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7006 net4488 vssd1 vssd1 vccd1 vccd1 net7530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7017 rbzero.wall_tracer.trackDistX\[1\] vssd1 vssd1 vccd1 vccd1 net7541 sky130_fd_sc_hd__dlygate4sd3_1
X_19238_ net5639 _03119_ _03121_ _03115_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7028 net4783 vssd1 vssd1 vccd1 vccd1 net7552 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6305 _04274_ vssd1 vssd1 vccd1 vccd1 net6829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6316 net2332 vssd1 vssd1 vccd1 vccd1 net6840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6327 rbzero.tex_r1\[21\] vssd1 vssd1 vccd1 vccd1 net6851 sky130_fd_sc_hd__dlygate4sd3_1
X_19169_ _03039_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__clkbuf_4
Xhold6338 net2340 vssd1 vssd1 vccd1 vccd1 net6862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5604 _00975_ vssd1 vssd1 vccd1 vccd1 net6128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6349 _04561_ vssd1 vssd1 vccd1 vccd1 net6873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21200_ _02750_ net4800 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5615 net3791 vssd1 vssd1 vccd1 vccd1 net6139 sky130_fd_sc_hd__dlygate4sd3_1
X_22180_ net312 net2719 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold5626 net3718 vssd1 vssd1 vccd1 vccd1 net6150 sky130_fd_sc_hd__clkbuf_4
Xhold4903 rbzero.spi_registers.buf_vshift\[1\] vssd1 vssd1 vccd1 vccd1 net5427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5648 net3093 vssd1 vssd1 vccd1 vccd1 net6172 sky130_fd_sc_hd__buf_2
XFILLER_0_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4914 rbzero.pov.spi_buffer\[40\] vssd1 vssd1 vccd1 vccd1 net5438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5659 _00966_ vssd1 vssd1 vccd1 vccd1 net6183 sky130_fd_sc_hd__dlygate4sd3_1
X_21131_ net4740 _04017_ _04014_ _04117_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4925 rbzero.pov.spi_buffer\[48\] vssd1 vssd1 vccd1 vccd1 net5449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4936 _00825_ vssd1 vssd1 vccd1 vccd1 net5460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4947 net985 vssd1 vssd1 vccd1 vccd1 net5471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4958 _03714_ vssd1 vssd1 vccd1 vccd1 net5482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4969 net2908 vssd1 vssd1 vccd1 vccd1 net5493 sky130_fd_sc_hd__dlygate4sd3_1
X_21062_ net4130 net4395 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__or2_1
X_20013_ _03261_ net3656 vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21964_ net189 net2483 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ clknet_leaf_95_i_clk net1439 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ clknet_1_1__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__buf_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22447_ clknet_leaf_69_i_clk _01616_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12200_ _05341_ _05348_ _05357_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__and3b_1
XFILLER_0_161_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ _06317_ _06335_ _06326_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__o21ai_1
Xhold6850 _10574_ vssd1 vssd1 vccd1 vccd1 net7374 sky130_fd_sc_hd__dlygate4sd3_1
X_22378_ net510 net2486 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6883 _09297_ vssd1 vssd1 vccd1 vccd1 net7407 sky130_fd_sc_hd__buf_2
X_12131_ net4058 _04602_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__xnor2_1
X_21329_ clknet_leaf_36_i_clk net4256 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12062_ rbzero.tex_r1\[63\] rbzero.tex_r1\[62\] _05230_ vssd1 vssd1 vccd1 vccd1 _05231_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold490 _03501_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ net2442 net5831 _04377_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__mux2_1
X_16870_ net3979 vssd1 vssd1 vccd1 vccd1 _09929_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15821_ _08891_ _08894_ _08895_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__a21o_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18540_ _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__buf_4
X_15752_ _08807_ _08826_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__xor2_2
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _06119_ _06110_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__or2b_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 net6064 vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _07851_ _07853_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__nor2_1
X_11915_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _05077_ vssd1 vssd1 vccd1 vccd1 _05085_
+ sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _02491_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15683_ _08753_ _08756_ _08757_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__nand3_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ net35 vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__buf_2
XFILLER_0_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _10302_ _10420_ _10421_ vssd1 vssd1 vccd1 vccd1 _10422_ sky130_fd_sc_hd__nand3_1
XFILLER_0_158_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14634_ _07767_ _07783_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__nor2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ _05003_ _05015_ _04999_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _10351_ _10352_ vssd1 vssd1 vccd1 vccd1 _10353_ sky130_fd_sc_hd__nor2_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ net1886 _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14565_ _07702_ _07711_ _07713_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_1__f__03991_ clknet_0__03991_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03991_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16304_ _09373_ _09377_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10728_ net2222 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__clkbuf_1
X_13516_ _06665_ _06619_ _06666_ _06628_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__a31o_4
XFILLER_0_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17284_ _09064_ _09484_ _09603_ _09103_ vssd1 vssd1 vccd1 vccd1 _10285_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ _07644_ _07646_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19023_ net2979 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__clkbuf_2
X_16235_ _09307_ _09308_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ net2083 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ net4947 _06497_ _06499_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_8_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20784__210 clknet_1_0__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__inv_2
XFILLER_0_152_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16166_ _09238_ _09240_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__xor2_1
X_13378_ _06478_ net82 _06517_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ _08218_ _08229_ net3631 _08215_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__o211a_1
X_12329_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _05493_ vssd1 vssd1 vccd1 vccd1 _05497_
+ sky130_fd_sc_hd__mux2_1
X_16097_ _09036_ _09078_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3509 _04805_ vssd1 vssd1 vccd1 vccd1 net4033 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_167_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19925_ net3580 _03477_ _03532_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a211o_1
X_15048_ _08180_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2808 net4726 vssd1 vssd1 vccd1 vccd1 net3332 sky130_fd_sc_hd__clkbuf_2
Xhold2819 _03894_ vssd1 vssd1 vccd1 vccd1 net3343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19856_ net6008 _08402_ _03484_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18807_ net4625 rbzero.wall_tracer.rayAddendY\[-1\] vssd1 vssd1 vccd1 vccd1 _02799_
+ sky130_fd_sc_hd__or2_1
X_19787_ net3022 _03442_ net2015 _03441_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__o211a_1
X_16999_ _06205_ vssd1 vssd1 vccd1 vccd1 _10010_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18738_ net6188 net3804 _06394_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18669_ _02646_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__inv_2
XFILLER_0_176_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21680_ clknet_leaf_35_i_clk net5324 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdxw\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__04008_ _04008_ vssd1 vssd1 vccd1 vccd1 clknet_0__04008_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20631_ net4060 _05816_ _03032_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20562_ net3030 net3705 _03911_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22301_ net433 net2460 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6102 net1891 vssd1 vssd1 vccd1 vccd1 net6626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6113 _04370_ vssd1 vssd1 vccd1 vccd1 net6637 sky130_fd_sc_hd__dlygate4sd3_1
X_20493_ _03858_ net3338 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__and2_1
Xhold6124 net1772 vssd1 vssd1 vccd1 vccd1 net6648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6135 rbzero.spi_registers.buf_texadd3\[6\] vssd1 vssd1 vccd1 vccd1 net6659 sky130_fd_sc_hd__dlygate4sd3_1
X_22232_ net364 net2516 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold5401 _04595_ vssd1 vssd1 vccd1 vccd1 net5925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6146 net1850 vssd1 vssd1 vccd1 vccd1 net6670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5412 _04456_ vssd1 vssd1 vccd1 vccd1 net5936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6157 rbzero.spi_registers.buf_texadd2\[2\] vssd1 vssd1 vccd1 vccd1 net6681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5423 net2791 vssd1 vssd1 vccd1 vccd1 net5947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6168 net1906 vssd1 vssd1 vccd1 vccd1 net6692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6179 rbzero.tex_r0\[41\] vssd1 vssd1 vccd1 vccd1 net6703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5434 rbzero.map_overlay.i_othery\[2\] vssd1 vssd1 vccd1 vccd1 net5958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4700 net850 vssd1 vssd1 vccd1 vccd1 net5224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5445 net2611 vssd1 vssd1 vccd1 vccd1 net5969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5456 rbzero.tex_r1\[29\] vssd1 vssd1 vccd1 vccd1 net5980 sky130_fd_sc_hd__dlygate4sd3_1
X_22163_ net295 net752 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold4711 rbzero.spi_registers.buf_texadd0\[3\] vssd1 vssd1 vccd1 vccd1 net5235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5467 net1555 vssd1 vssd1 vccd1 vccd1 net5991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4722 rbzero.spi_registers.buf_vshift\[0\] vssd1 vssd1 vccd1 vccd1 net5246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5478 net2879 vssd1 vssd1 vccd1 vccd1 net6002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4733 net938 vssd1 vssd1 vccd1 vccd1 net5257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4744 _00732_ vssd1 vssd1 vccd1 vccd1 net5268 sky130_fd_sc_hd__dlygate4sd3_1
X_21114_ _04098_ _04099_ _04100_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5489 rbzero.map_overlay.i_otherx\[2\] vssd1 vssd1 vccd1 vccd1 net6013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4755 net973 vssd1 vssd1 vccd1 vccd1 net5279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4766 rbzero.spi_registers.texadd3\[22\] vssd1 vssd1 vccd1 vccd1 net5290 sky130_fd_sc_hd__dlygate4sd3_1
X_22094_ clknet_leaf_49_i_clk net3938 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold4777 rbzero.spi_registers.buf_vshift\[4\] vssd1 vssd1 vccd1 vccd1 net5301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4788 net885 vssd1 vssd1 vccd1 vccd1 net5312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21045_ net5310 net5455 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nand2_1
Xhold4799 _00849_ vssd1 vssd1 vccd1 vccd1 net5323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21947_ net172 net2410 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _04864_ _04865_ _04866_ _04867_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a221o_1
X_12680_ _05841_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ clknet_leaf_98_i_clk net1287 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ net4971 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__buf_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14350_ _07450_ _07496_ _07499_ _07500_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__o31a_1
X_11562_ _04691_ _04694_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13301_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14281_ _07386_ _07408_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11493_ _04656_ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16020_ _09090_ _08664_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__or3b_2
XFILLER_0_126_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13232_ net4911 net4900 _06387_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7392 net4367 vssd1 vssd1 vccd1 vccd1 net7916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6680 rbzero.spi_registers.ss_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net7204 sky130_fd_sc_hd__dlygate4sd3_1
X_13163_ net3155 vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__inv_2
Xhold6691 net2544 vssd1 vssd1 vccd1 vccd1 net7215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _05279_ _05280_ _05282_ _05061_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5990 net1428 vssd1 vssd1 vccd1 vccd1 net6514 sky130_fd_sc_hd__dlygate4sd3_1
X_17971_ _01937_ _01940_ _01938_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__o21ai_1
X_13094_ _04837_ _06217_ _06248_ rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1
+ vccd1 _06250_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19710_ _02998_ _03393_ net1869 _03400_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__o211a_1
X_12045_ rbzero.tex_r1\[55\] rbzero.tex_r1\[54\] _05072_ vssd1 vssd1 vccd1 vccd1 _05214_
+ sky130_fd_sc_hd__mux2_1
X_16922_ net4155 _09941_ _09942_ net7554 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19641_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__clkbuf_4
X_16853_ _04241_ net3979 vssd1 vssd1 vccd1 vccd1 _09920_ sky130_fd_sc_hd__nor2_4
X_15804_ _08875_ _08878_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19572_ net5079 _03302_ _03318_ _03314_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__o211a_1
X_16784_ _09064_ _09477_ vssd1 vssd1 vccd1 vccd1 _09854_ sky130_fd_sc_hd__or2_1
X_13996_ _07145_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18523_ net3837 net1076 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15735_ _08548_ net4954 vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _06096_ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__or2b_1
XFILLER_0_198_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20816__239 clknet_1_1__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__inv_2
X_18454_ _02477_ _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__xnor2_1
X_15666_ _08730_ _08740_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__xnor2_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ net57 _06008_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17405_ _10293_ _10296_ _10404_ vssd1 vssd1 vccd1 vccd1 _10405_ sky130_fd_sc_hd__a21bo_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07753_ _07759_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__xor2_2
X_11829_ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__clkbuf_8
X_18385_ _02418_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15597_ _08548_ _08549_ _08347_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__a21oi_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _10333_ _10334_ _10209_ _10335_ vssd1 vssd1 vccd1 vccd1 _10336_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14548_ _06990_ _07354_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17267_ _08717_ _08582_ vssd1 vssd1 vccd1 vccd1 _10268_ sky130_fd_sc_hd__nor2_1
X_14479_ _07617_ _07628_ _07629_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ net3904 _02973_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16218_ _09280_ _09291_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17198_ _10198_ _10199_ vssd1 vssd1 vccd1 vccd1 _10200_ sky130_fd_sc_hd__xor2_4
XFILLER_0_102_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4007 rbzero.row_render.side vssd1 vssd1 vccd1 vccd1 net4531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4018 net1456 vssd1 vssd1 vccd1 vccd1 net4542 sky130_fd_sc_hd__dlygate4sd3_1
X_16149_ _08615_ _08607_ _08173_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__o21ai_1
Xhold4029 _00599_ vssd1 vssd1 vccd1 vccd1 net4553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3306 net7337 vssd1 vssd1 vccd1 vccd1 net3830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3317 _01011_ vssd1 vssd1 vccd1 vccd1 net3841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3328 net4686 vssd1 vssd1 vccd1 vccd1 net3852 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3339 net4711 vssd1 vssd1 vccd1 vccd1 net3863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2605 _03103_ vssd1 vssd1 vccd1 vccd1 net3129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2616 net7351 vssd1 vssd1 vccd1 vccd1 net3140 sky130_fd_sc_hd__dlygate4sd3_1
X_19908_ net4355 _03480_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nor2_1
Xhold2627 _02494_ vssd1 vssd1 vccd1 vccd1 net3151 sky130_fd_sc_hd__buf_2
Xhold2638 net7494 vssd1 vssd1 vccd1 vccd1 net3162 sky130_fd_sc_hd__buf_1
Xhold1904 net5825 vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 net7742 vssd1 vssd1 vccd1 vccd1 net3173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1915 net7063 vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1926 _04457_ vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
X_19839_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__buf_2
Xhold1937 net7126 vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1948 net5827 vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1959 _01133_ vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21801_ clknet_leaf_89_i_clk net4357 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21732_ clknet_leaf_22_i_clk net5731 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20756__186 clknet_1_1__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__inv_2
XFILLER_0_8_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21663_ clknet_leaf_35_i_clk net5549 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20614_ net4002 _04802_ net4015 _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21594_ clknet_leaf_23_i_clk net5752 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20545_ net3648 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ net951 net3412 _03845_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5220 _00709_ vssd1 vssd1 vccd1 vccd1 net5744 sky130_fd_sc_hd__dlygate4sd3_1
X_22215_ net347 net2899 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
Xhold5231 _03268_ vssd1 vssd1 vccd1 vccd1 net5755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5242 rbzero.pov.spi_buffer\[55\] vssd1 vssd1 vccd1 vccd1 net5766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5253 net1489 vssd1 vssd1 vccd1 vccd1 net5777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5264 net1721 vssd1 vssd1 vccd1 vccd1 net5788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5275 _04198_ vssd1 vssd1 vccd1 vccd1 net5799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4530 _00745_ vssd1 vssd1 vccd1 vccd1 net5054 sky130_fd_sc_hd__dlygate4sd3_1
X_22146_ net278 net2287 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
Xhold5286 rbzero.tex_r1\[37\] vssd1 vssd1 vccd1 vccd1 net5810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4541 net807 vssd1 vssd1 vccd1 vccd1 net5065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5297 net588 vssd1 vssd1 vccd1 vccd1 net5821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4552 net819 vssd1 vssd1 vccd1 vccd1 net5076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4563 net837 vssd1 vssd1 vccd1 vccd1 net5087 sky130_fd_sc_hd__dlygate4sd3_1
X_20921__334 clknet_1_0__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__inv_2
Xhold4574 rbzero.spi_registers.buf_mapdx\[5\] vssd1 vssd1 vccd1 vccd1 net5098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3840 _03584_ vssd1 vssd1 vccd1 vccd1 net4364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4585 rbzero.spi_registers.buf_otherx\[3\] vssd1 vssd1 vccd1 vccd1 net5109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3851 net7900 vssd1 vssd1 vccd1 vccd1 net4375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4596 rbzero.spi_registers.buf_texadd0\[11\] vssd1 vssd1 vccd1 vccd1 net5120 sky130_fd_sc_hd__dlygate4sd3_1
X_22077_ clknet_leaf_9_i_clk net3527 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3862 net3143 vssd1 vssd1 vccd1 vccd1 net4386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3873 net712 vssd1 vssd1 vccd1 vccd1 net4397 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03994_ clknet_0__03994_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03994_
+ sky130_fd_sc_hd__clkbuf_16
X_21028_ _04029_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__and2b_1
Xhold3884 _00995_ vssd1 vssd1 vccd1 vccd1 net4408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3895 _03610_ vssd1 vssd1 vccd1 vccd1 net4419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13850_ _06880_ _06889_ net529 _06895_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ _05201_ _05946_ _05956_ net73 _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ net6529 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__clkbuf_1
X_13781_ _06931_ _06884_ _06886_ _06880_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__and4b_1
XFILLER_0_167_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _04646_ _06138_ _08295_ _08594_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__o211a_2
X_12732_ _05892_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _08461_ _08510_ _08525_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__a21boi_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ net6265 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__buf_4
XFILLER_0_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _07507_ _07506_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18170_ _02131_ _02132_ _02134_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a21bo_1
X_11614_ _04784_ _04785_ _04725_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__o21a_1
X_15382_ _08444_ _08456_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__nor2_1
X_12594_ _05177_ _05756_ _05758_ _05010_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o211a_1
X_17121_ _09847_ _10094_ _10121_ vssd1 vssd1 vccd1 vccd1 _10123_ sky130_fd_sc_hd__nand3_1
XFILLER_0_154_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ _07479_ _07480_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ _04701_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nand2_1
X_17052_ _10057_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14264_ _07369_ _07410_ _07413_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__nand3_1
X_11476_ _04646_ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16003_ _09036_ _09037_ _09039_ _09077_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__nand4_2
X_13215_ _06219_ net4897 _06370_ _06216_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _07345_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ net3381 _06298_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__and2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _01778_ _08793_ _02000_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__o21ai_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ net3952 _06181_ _06221_ net3995 vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20896__311 clknet_1_1__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__inv_2
XFILLER_0_100_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12028_ _04806_ _05192_ _05195_ _05196_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__a41o_1
X_16905_ net5310 _09939_ _09940_ net3262 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__a22o_1
X_17885_ _01910_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16836_ _09904_ _09905_ vssd1 vssd1 vccd1 vccd1 _09906_ sky130_fd_sc_hd__or2_2
X_19624_ net3072 _03340_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__or2_1
XFILLER_0_206_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19555_ net824 _03303_ _03309_ _03295_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__o211a_1
X_16767_ _09835_ _09836_ vssd1 vssd1 vccd1 vccd1 _09837_ sky130_fd_sc_hd__nor2_1
X_13979_ _06876_ _06970_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ net44 _02488_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__and2_1
X_15718_ net6098 _08299_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__nand2_4
XFILLER_0_38_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19486_ net2541 _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__or2_1
X_16698_ _09652_ _09768_ vssd1 vssd1 vccd1 vccd1 _09769_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _02462_ net7789 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _08454_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ _02403_ net4489 _02338_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17319_ _10219_ _10319_ vssd1 vssd1 vccd1 vccd1 _10320_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18299_ _02334_ _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03988_ _03988_ vssd1 vssd1 vccd1 vccd1 clknet_0__03988_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20261_ net3476 net4839 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22000_ net225 net1463 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold3103 net652 vssd1 vssd1 vccd1 vccd1 net3627 sky130_fd_sc_hd__clkbuf_2
X_20192_ net3782 _03718_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3114 _03799_ vssd1 vssd1 vccd1 vccd1 net3638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3125 _01231_ vssd1 vssd1 vccd1 vccd1 net3649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3136 net1230 vssd1 vssd1 vccd1 vccd1 net3660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3147 _03929_ vssd1 vssd1 vccd1 vccd1 net3671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2402 net6018 vssd1 vssd1 vccd1 vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2413 net7329 vssd1 vssd1 vccd1 vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3158 _01242_ vssd1 vssd1 vccd1 vccd1 net3682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 net6046 vssd1 vssd1 vccd1 vccd1 net2948 sky130_fd_sc_hd__buf_1
Xhold3169 net4781 vssd1 vssd1 vccd1 vccd1 net3693 sky130_fd_sc_hd__dlygate4sd3_1
X_20762__190 clknet_1_0__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__inv_2
Xhold2435 net7736 vssd1 vssd1 vccd1 vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1701 _04193_ vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2446 net3108 vssd1 vssd1 vccd1 vccd1 net2970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1712 _01425_ vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2457 _00650_ vssd1 vssd1 vccd1 vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1723 net7076 vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2468 net4295 vssd1 vssd1 vccd1 vccd1 net2992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _00885_ vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2479 net6126 vssd1 vssd1 vccd1 vccd1 net3003 sky130_fd_sc_hd__clkbuf_2
Xhold1745 net6953 vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1756 net4267 vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1767 _01166_ vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1778 net6999 vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1789 net6923 vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21715_ clknet_leaf_17_i_clk net2092 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21646_ clknet_leaf_33_i_clk net1609 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21577_ clknet_leaf_4_i_clk net4217 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_60 _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_71 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ net7014 net6728 _04540_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__mux2_1
XANTENNA_93 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20528_ _03880_ net3436 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11261_ _04168_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__clkbuf_4
X_20459_ net3835 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5050 rbzero.pov.spi_buffer\[19\] vssd1 vssd1 vccd1 vccd1 net5574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5061 net1162 vssd1 vssd1 vccd1 vccd1 net5585 sky130_fd_sc_hd__dlygate4sd3_1
X_13000_ _06154_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11192_ net2188 net6425 _04470_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__mux2_1
Xhold5072 net1309 vssd1 vssd1 vccd1 vccd1 net5596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5083 net1256 vssd1 vssd1 vccd1 vccd1 net5607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5094 rbzero.spi_registers.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 net5618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4360 net2122 vssd1 vssd1 vccd1 vccd1 net4884 sky130_fd_sc_hd__dlygate4sd3_1
X_22129_ net261 net1399 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold4371 net2941 vssd1 vssd1 vccd1 vccd1 net4895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4382 _01642_ vssd1 vssd1 vccd1 vccd1 net4906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4393 _06383_ vssd1 vssd1 vccd1 vccd1 net4917 sky130_fd_sc_hd__buf_1
Xhold3670 net7649 vssd1 vssd1 vccd1 vccd1 net4194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3681 net7654 vssd1 vssd1 vccd1 vccd1 net4205 sky130_fd_sc_hd__dlygate4sd3_1
X_14951_ net4374 _08096_ _08027_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3692 _00746_ vssd1 vssd1 vccd1 vccd1 net4216 sky130_fd_sc_hd__dlygate4sd3_1
X_13902_ _07051_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nor2_1
X_17670_ _01718_ _01720_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__and2_1
Xhold2980 net7467 vssd1 vssd1 vccd1 vccd1 net3504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2991 _03933_ vssd1 vssd1 vccd1 vccd1 net3515 sky130_fd_sc_hd__dlygate4sd3_1
X_14882_ _07991_ _07989_ _08031_ _06707_ vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__a211o_1
X_16621_ _09569_ _09578_ _09576_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13833_ _06980_ _06951_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19340_ net1787 _03173_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__or2_1
X_16552_ _09621_ _09623_ vssd1 vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20739__170 clknet_1_1__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__inv_2
X_13764_ _06736_ _06860_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__or3_4
X_10976_ net6858 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap84 _06429_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlymetal6s2s_1
X_15503_ _04646_ net8126 _08295_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__o211a_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19271_ net5042 _03132_ _03139_ _03128_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__o211a_1
X_12715_ _04162_ net3993 net10 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__mux2_1
X_16483_ _09423_ _09432_ _09554_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__o21a_1
X_13695_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__buf_6
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18222_ _02174_ _02175_ _02249_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a21o_1
X_15434_ _08507_ _08508_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__and2b_1
X_12646_ net46 _05785_ _05796_ _05787_ net43 vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18153_ _02180_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__xor2_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15365_ net3008 _08418_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__nand2_1
X_12577_ _04984_ _05741_ _05000_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__o21a_1
X_17104_ _10104_ _10105_ vssd1 vssd1 vccd1 vccd1 _10106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _07466_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18084_ _09231_ _08793_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ rbzero.spi_registers.texadd3\[21\] rbzero.spi_registers.texadd1\[21\] rbzero.spi_registers.texadd0\[21\]
+ rbzero.spi_registers.texadd2\[21\] _04692_ _04693_ vssd1 vssd1 vccd1 vccd1 _04700_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15296_ net3057 _08303_ _08306_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 net5080 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17035_ net4560 net4399 vssd1 vssd1 vccd1 vccd1 _10042_ sky130_fd_sc_hd__nor2_1
Xhold319 net5242 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03773_ _03773_ vssd1 vssd1 vccd1 vccd1 clknet_0__03773_ sky130_fd_sc_hd__clkbuf_16
X_14247_ _07362_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__xor2_4
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ net7582 net3403 _04631_ _04633_ _04628_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14178_ _06881_ _07082_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13129_ net3566 vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ net3855 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 net6230 vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ _01984_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nor2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 net6548 vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17868_ _01916_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19607_ net798 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16819_ _09747_ _09749_ vssd1 vssd1 vccd1 vccd1 _09889_ sky130_fd_sc_hd__nor2_1
X_17799_ _01724_ _01725_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__nor2_1
X_19538_ net5360 _03288_ _03297_ _03295_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19469_ _03088_ net3078 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20950__360 clknet_1_1__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__inv_2
X_21500_ clknet_leaf_14_i_clk net4347 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22480_ clknet_leaf_67_i_clk net1137 vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21431_ clknet_leaf_82_i_clk net2886 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21362_ clknet_leaf_55_i_clk _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 net5433 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
X_21293_ clknet_leaf_75_i_clk net4080 vssd1 vssd1 vccd1 vccd1 reg_rgb\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold831 net3751 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold842 net3448 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
X_20244_ net5623 _03743_ _03749_ _03748_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__o211a_1
Xhold853 net5613 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 _01155_ vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold875 _01298_ vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold886 net5483 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold897 net5640 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
X_20175_ net5520 _03704_ _03710_ _03709_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__o211a_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2210 net7136 vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2221 _01319_ vssd1 vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2232 net7281 vssd1 vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2243 _01417_ vssd1 vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2254 net2854 vssd1 vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2265 net5977 vssd1 vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__clkbuf_2
Xhold1520 net5809 vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2276 _04541_ vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1531 _04287_ vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2287 _01121_ vssd1 vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1542 net6817 vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1553 _03365_ vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2298 _01578_ vssd1 vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1564 net3111 vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 _01397_ vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1586 net6915 vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1597 _01294_ vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ net2055 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10761_ net2680 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _05457_ vssd1 vssd1 vccd1 vccd1 _05666_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ net2485 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__clkbuf_1
X_13480_ _06543_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12431_ _04982_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21629_ clknet_leaf_2_i_clk net5108 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15150_ net4727 _08074_ _08249_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net6168 _04817_ _04820_ _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__o22a_1
X_14101_ _07150_ _07187_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__or2_4
X_11313_ net2800 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12293_ _05009_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__buf_4
X_15081_ net4597 net4591 _08191_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11244_ net2797 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
X_14032_ _07163_ _07181_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net6814 net7239 _04459_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__mux2_1
X_18840_ _02828_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4190 net3171 vssd1 vssd1 vccd1 vccd1 net4714 sky130_fd_sc_hd__buf_1
XFILLER_0_140_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18771_ net1091 _02528_ _02529_ net4552 _02766_ vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ _09056_ _09057_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17722_ _01770_ _01771_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nand2_1
X_14934_ net7908 _08017_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__nand2_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04010_ clknet_0__04010_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04010_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__xor2_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _08006_ _08008_ _08010_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__o31a_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16604_ _08409_ _08795_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__nor2_1
X_13816_ _06876_ net529 net577 vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__or3_1
X_17584_ _10502_ _10579_ _10580_ vssd1 vssd1 vccd1 vccd1 _10582_ sky130_fd_sc_hd__and3_1
X_14796_ _07205_ _07305_ _07941_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ net5007 _03159_ _03169_ _03168_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16535_ _08180_ _09605_ net77 _08296_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__a31o_1
X_13747_ _06844_ _06881_ _06827_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__or3b_4
X_10959_ net2490 net6433 _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19254_ net4115 _03120_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__or2_1
X_16466_ _09537_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13678_ _06725_ _06794_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18205_ _02250_ _02251_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__nor2_1
X_15417_ _08490_ _08491_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__nand2_1
X_19185_ _03088_ net2965 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__or2_1
X_12629_ _05790_ net8 vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nor2_1
X_16397_ _08684_ _08588_ vssd1 vssd1 vccd1 vccd1 _09470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6509 rbzero.tex_g1\[36\] vssd1 vssd1 vccd1 vccd1 net7033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18136_ _01802_ _09732_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__nor2_1
X_15348_ _08393_ _08405_ _08411_ _08422_ vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__or4_1
Xhold5808 rbzero.tex_b0\[10\] vssd1 vssd1 vccd1 vccd1 net6332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5819 net828 vssd1 vssd1 vccd1 vccd1 net6343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18067_ _01999_ _02014_ _02012_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a21o_1
Xhold105 _00576_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ net4893 net3024 net4355 vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__or3_1
Xhold116 _03557_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold127 net4963 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net4958 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _10024_ _10025_ _10026_ vssd1 vssd1 vccd1 vccd1 _10027_ sky130_fd_sc_hd__a21oi_1
Xhold149 rbzero.wall_tracer.visualWallDist\[0\] vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_1
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18969_ net3996 _02261_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__nor2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21980_ net205 net1198 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20874__291 clknet_1_1__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__inv_2
XFILLER_0_37_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22463_ clknet_leaf_39_i_clk _01632_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21414_ clknet_leaf_84_i_clk net4670 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_22394_ net146 net2084 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21345_ clknet_leaf_40_i_clk net4188 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21276_ clknet_leaf_59_i_clk _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold650 _01265_ vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 net5558 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 net6428 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 net6434 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20227_ net5205 _03730_ _03739_ _03735_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__o211a_1
Xhold694 _03184_ vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20158_ net5500 _03691_ _03700_ _03696_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__o211a_1
Xhold2040 _01460_ vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2051 _04178_ vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2062 _01280_ vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2073 _04486_ vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_20089_ net3225 net4795 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__nand2_1
X_12980_ _06131_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__inv_2
Xhold2084 net6977 vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2095 net7222 vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1350 net5889 vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 _00906_ vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1372 _01140_ vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ net4303 net4271 _05022_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__or4_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 _04531_ vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 net6717 vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _07444_ _07523_ _07800_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__or3_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _04988_ vssd1 vssd1 vccd1 vccd1 _05032_
+ sky130_fd_sc_hd__mux2_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _06743_ _06656_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__nor2_1
X_10813_ net6944 net2641 _04277_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14581_ _07721_ _07730_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nor2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04915_ _04916_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__nand2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16320_ _09247_ _09264_ _09245_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ _06654_ _06682_ _06650_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__o21ai_2
X_10744_ _04167_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__clkinv_8
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16251_ _09208_ _09213_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13463_ _06421_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__inv_2
X_10675_ net6760 net7056 _04203_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ net4084 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12414_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _05457_ vssd1 vssd1 vccd1 vccd1 _05581_
+ sky130_fd_sc_hd__mux2_1
X_16182_ _08726_ _08728_ _09255_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13394_ net4947 _06479_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__nor2_4
XFILLER_0_180_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _08218_ _08240_ net6136 _08239_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__o211a_1
X_12345_ _05511_ _05512_ _04981_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15064_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1 vccd1 vccd1 _08193_
+ sky130_fd_sc_hd__inv_2
X_19941_ net6207 _03530_ net2893 _03550_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__o211a_1
X_12276_ net83 _05323_ net4006 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__o21ai_1
X_14015_ _07127_ _07128_ _07132_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__a21o_1
X_11227_ net5874 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19872_ net3821 _08479_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__or2_1
X_18823_ _02812_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__nand2_1
X_11158_ net1519 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15966_ _09014_ _09040_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__xnor2_1
X_11089_ net6914 net6770 _04415_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__mux2_1
X_18754_ net4799 net941 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17705_ _01732_ _01734_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or2_1
X_14917_ _07995_ _08041_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__nand2_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ _08970_ _08971_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__xor2_1
X_18685_ _02686_ _02687_ net4811 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17636_ _01686_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14848_ _07997_ _07998_ _06690_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17567_ _10465_ _10466_ _10565_ vssd1 vssd1 vccd1 vccd1 _10566_ sky130_fd_sc_hd__a21oi_1
X_14779_ _07923_ _07929_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16518_ _09588_ _09589_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__xor2_1
X_19306_ _03039_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__buf_2
X_17498_ _10356_ _10365_ _10363_ vssd1 vssd1 vccd1 vccd1 _10497_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7007 rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1 vccd1 net7531 sky130_fd_sc_hd__dlygate4sd3_1
X_16449_ net3003 net7428 _08293_ vssd1 vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__mux2_1
X_19237_ net5318 _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__or2_1
Xhold7018 rbzero.wall_tracer.trackDistY\[4\] vssd1 vssd1 vccd1 vccd1 net7542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7029 _00511_ vssd1 vssd1 vccd1 vccd1 net7553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6306 net1819 vssd1 vssd1 vccd1 vccd1 net6830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19168_ _03036_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6317 rbzero.tex_b1\[47\] vssd1 vssd1 vccd1 vccd1 net6841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6328 net2007 vssd1 vssd1 vccd1 vccd1 net6852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6339 _04513_ vssd1 vssd1 vccd1 vccd1 net6863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18119_ _01980_ _01981_ _02064_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5605 rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 net6129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5616 rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1 net6140 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5627 _08236_ vssd1 vssd1 vccd1 vccd1 net6151 sky130_fd_sc_hd__dlygate4sd3_1
X_19099_ _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__buf_4
Xhold5638 net7886 vssd1 vssd1 vccd1 vccd1 net6162 sky130_fd_sc_hd__clkbuf_4
X_21130_ _04113_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__xnor2_1
Xhold4904 net1006 vssd1 vssd1 vccd1 vccd1 net5428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5649 _00933_ vssd1 vssd1 vccd1 vccd1 net6173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4915 net1491 vssd1 vssd1 vccd1 vccd1 net5439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4926 _01084_ vssd1 vssd1 vccd1 vccd1 net5450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4937 net1059 vssd1 vssd1 vccd1 vccd1 net5461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4948 _00504_ vssd1 vssd1 vccd1 vccd1 net5472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4959 _01063_ vssd1 vssd1 vccd1 vccd1 net5483 sky130_fd_sc_hd__dlygate4sd3_1
X_21061_ _04053_ _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20012_ rbzero.debug_overlay.facingY\[-5\] net3547 _03594_ vssd1 vssd1 vccd1 vccd1
+ _03607_ sky130_fd_sc_hd__mux2_1
X_20679__116 clknet_1_0__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__inv_2
X_21963_ net188 net2032 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21894_ clknet_leaf_95_i_clk net1410 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22446_ clknet_leaf_70_i_clk _01615_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6840 gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 net7364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6851 _10576_ vssd1 vssd1 vccd1 vccd1 net7375 sky130_fd_sc_hd__dlygate4sd3_1
X_22377_ net509 net2375 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6884 rbzero.wall_tracer.trackDistX\[6\] vssd1 vssd1 vccd1 vccd1 net7408 sky130_fd_sc_hd__dlygate4sd3_1
X_12130_ _04831_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__buf_4
X_21328_ clknet_leaf_36_i_clk net4282 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12061_ _05070_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__clkbuf_8
X_21259_ clknet_leaf_52_i_clk net3224 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 net5352 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 net4220 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ net5881 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__clkbuf_1
X_15820_ _08892_ _08893_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__and2_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _08823_ _08824_ _08825_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__a21oi_2
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__nand2_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20890__306 clknet_1_0__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__inv_2
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 _03363_ vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1191 net6655 vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _07845_ _07849_ _07850_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__and3_1
XFILLER_0_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11914_ _05080_ _05083_ _05009_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__mux2_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ net4326 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__buf_2
X_15682_ _08557_ _08625_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ net38 _06047_ _06049_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a22o_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _10418_ _10419_ _10417_ vssd1 vssd1 vccd1 vccd1 _10421_ sky130_fd_sc_hd__a21o_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14633_ _07767_ _07783_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__xor2_2
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11845_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _05014_ vssd1 vssd1 vccd1 vccd1 _05015_
+ sky130_fd_sc_hd__mux2_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _10349_ _10350_ vssd1 vssd1 vccd1 vccd1 _10352_ sky130_fd_sc_hd__and2_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _07668_ _07682_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__xnor2_4
Xclkbuf_1_1__f__03990_ clknet_0__03990_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03990_
+ sky130_fd_sc_hd__clkbuf_16
X_11776_ _04942_ _04941_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__nand2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16303_ _08618_ _08665_ _09376_ _09229_ _09223_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__a32o_1
XFILLER_0_144_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13515_ _06428_ _06620_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__xor2_4
X_10727_ net6898 net7073 _04225_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
X_17283_ _09103_ _09064_ _09483_ _09603_ vssd1 vssd1 vccd1 vccd1 _10284_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14495_ _07645_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19022_ net3945 net88 net2978 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__or3b_1
X_16234_ _09133_ _09306_ _09252_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__a21boi_1
X_13446_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__inv_2
X_10658_ net5821 net6848 _04192_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16165_ _08573_ _08654_ _09239_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13377_ _06432_ _06434_ _06470_ net4947 _06485_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15116_ net6123 _08223_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__or2_1
X_12328_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _05070_ vssd1 vssd1 vccd1 vccd1 _05496_
+ sky130_fd_sc_hd__mux2_1
X_16096_ _09121_ _09169_ _09170_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19924_ _08414_ _03476_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nor2_1
X_15047_ net7433 _06715_ _08135_ _08179_ _06625_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__o311a_2
X_12259_ _04889_ _05196_ _05426_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__or4_1
X_19855_ net4338 _03475_ net3032 _03454_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__o211a_1
X_18806_ _05391_ rbzero.wall_tracer.rayAddendY\[-1\] vssd1 vssd1 vccd1 vccd1 _02798_
+ sky130_fd_sc_hd__nand2_1
X_19786_ net2014 _03443_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ _10005_ _10008_ vssd1 vssd1 vccd1 vccd1 _10009_ sky130_fd_sc_hd__xnor2_1
X_18737_ net4387 _10019_ net6187 _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
X_15949_ _09019_ _09023_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__xor2_1
XFILLER_0_211_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18668_ net4696 _02666_ net7571 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ _10584_ _01670_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18599_ _02609_ _02610_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__04007_ _04007_ vssd1 vssd1 vccd1 vccd1 clknet_0__04007_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20630_ _05816_ _03032_ _03966_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20561_ net3260 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22300_ net432 net2145 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6103 _04202_ vssd1 vssd1 vccd1 vccd1 net6627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20492_ net3337 net1491 _03867_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__mux2_1
Xhold6114 net1707 vssd1 vssd1 vccd1 vccd1 net6638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6125 rbzero.spi_registers.buf_texadd3\[13\] vssd1 vssd1 vccd1 vccd1 net6649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22231_ net363 net2601 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold6136 net1964 vssd1 vssd1 vccd1 vccd1 net6660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5402 net2651 vssd1 vssd1 vccd1 vccd1 net5926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6147 _04439_ vssd1 vssd1 vccd1 vccd1 net6671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5413 net2192 vssd1 vssd1 vccd1 vccd1 net5937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6158 net1787 vssd1 vssd1 vccd1 vccd1 net6682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6169 rbzero.spi_registers.buf_texadd3\[2\] vssd1 vssd1 vccd1 vccd1 net6693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5424 _00675_ vssd1 vssd1 vccd1 vccd1 net5948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5435 net2864 vssd1 vssd1 vccd1 vccd1 net5959 sky130_fd_sc_hd__dlygate4sd3_1
X_22162_ net294 net2193 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold4701 rbzero.spi_registers.buf_texadd0\[2\] vssd1 vssd1 vccd1 vccd1 net5225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5446 _00524_ vssd1 vssd1 vccd1 vccd1 net5970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4712 net894 vssd1 vssd1 vccd1 vccd1 net5236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5457 net2493 vssd1 vssd1 vccd1 vccd1 net5981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4723 net906 vssd1 vssd1 vccd1 vccd1 net5247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5468 rbzero.map_overlay.i_othery\[4\] vssd1 vssd1 vccd1 vccd1 net5992 sky130_fd_sc_hd__dlygate4sd3_1
X_21113_ _04018_ _04101_ _04102_ _03083_ net4649 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a32o_1
Xhold4734 rbzero.spi_registers.texadd1\[11\] vssd1 vssd1 vccd1 vccd1 net5258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5479 _00673_ vssd1 vssd1 vccd1 vccd1 net6003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4745 net972 vssd1 vssd1 vccd1 vccd1 net5269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4756 _00852_ vssd1 vssd1 vccd1 vccd1 net5280 sky130_fd_sc_hd__dlygate4sd3_1
X_22093_ clknet_leaf_49_i_clk net3931 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4767 net983 vssd1 vssd1 vccd1 vccd1 net5291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4778 net991 vssd1 vssd1 vccd1 vccd1 net5302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4789 rbzero.spi_registers.texadd1\[17\] vssd1 vssd1 vccd1 vccd1 net5313 sky130_fd_sc_hd__dlygate4sd3_1
X_21044_ net5310 net5455 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21946_ net171 net1359 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ clknet_leaf_98_i_clk net1225 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20733__165 clknet_1_0__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__inv_2
X_11561_ _04724_ _04729_ _04730_ _04731_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ _06448_ _06449_ _06450_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _07428_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11492_ rbzero.texu_hot\[2\] _04655_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13231_ _06344_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__or2_1
X_22429_ clknet_leaf_41_i_clk net4397 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7382 rbzero.wall_tracer.stepDistY\[10\] vssd1 vssd1 vccd1 vccd1 net7906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6670 rbzero.spi_registers.buf_texadd1\[15\] vssd1 vssd1 vccd1 vccd1 net7194 sky130_fd_sc_hd__dlygate4sd3_1
X_13162_ _06311_ _06313_ _06315_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6681 net1211 vssd1 vssd1 vccd1 vccd1 net7205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6692 rbzero.tex_g0\[18\] vssd1 vssd1 vccd1 vccd1 net7216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ _05068_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__or2_1
Xhold5980 net1383 vssd1 vssd1 vccd1 vccd1 net6504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5991 rbzero.tex_r1\[60\] vssd1 vssd1 vccd1 vccd1 net6515 sky130_fd_sc_hd__dlygate4sd3_1
X_17970_ _01987_ _02018_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ rbzero.debug_overlay.playerX\[5\] _06248_ net2611 net2807 vssd1 vssd1 vccd1
+ vccd1 _06249_ sky130_fd_sc_hd__a211o_1
X_12044_ _05207_ _05210_ _05212_ net4077 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a31o_1
X_16921_ net4136 _09941_ _09942_ net7440 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ net3075 net3151 net4327 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__or3_1
X_16852_ net3870 _04795_ _09919_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15803_ _08515_ _08877_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__xnor2_1
X_16783_ _09593_ _09595_ _09729_ _09727_ vssd1 vssd1 vccd1 vccd1 _09853_ sky130_fd_sc_hd__o31a_1
X_19571_ net3096 _03304_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or2_1
X_13995_ _07104_ _07106_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__xor2_2
XFILLER_0_204_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15734_ _08753_ _08756_ _08757_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__a21o_1
X_18522_ _02530_ _02538_ net4477 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15665_ _08738_ _08739_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__nor2_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _02468_ _02471_ _02469_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__a21bo_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ net54 _05998_ _06007_ net55 vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _09138_ _10174_ _10294_ vssd1 vssd1 vccd1 vccd1 _10404_ sky130_fd_sc_hd__or3_1
X_14616_ _07719_ _07731_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__xnor2_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _04957_ _04971_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__or3_1
X_18384_ _02417_ net4429 _02411_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15596_ _08367_ _08557_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__nor2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _10211_ vssd1 vssd1 vccd1 vccd1 _10335_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _07532_ _07400_ _07439_ _07534_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__o22ai_2
X_11759_ net923 net1569 vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ _10265_ _10266_ vssd1 vssd1 vccd1 vccd1 _10267_ sky130_fd_sc_hd__xor2_1
X_14478_ _07620_ _07627_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__nor2_1
X_16217_ _09280_ _09291_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__nand2_1
X_19005_ net3904 _02973_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13429_ _06572_ _06573_ _06576_ _06577_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__and4_1
X_17197_ _09792_ _09900_ _09899_ _09898_ vssd1 vssd1 vccd1 vccd1 _10199_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16148_ _08626_ _09222_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__nor2_1
Xhold4008 net3014 vssd1 vssd1 vccd1 vccd1 net4532 sky130_fd_sc_hd__buf_2
Xhold4019 _01601_ vssd1 vssd1 vccd1 vccd1 net4543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16079_ _09152_ _09153_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__nor2_1
Xhold3307 _03604_ vssd1 vssd1 vccd1 vccd1 net3831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3318 net5568 vssd1 vssd1 vccd1 vccd1 net3842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3329 net7346 vssd1 vssd1 vccd1 vccd1 net3853 sky130_fd_sc_hd__clkbuf_4
Xhold2606 _03104_ vssd1 vssd1 vccd1 vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
X_19907_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__clkbuf_4
Xhold2617 _03592_ vssd1 vssd1 vccd1 vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2628 _03460_ vssd1 vssd1 vccd1 vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2639 net7757 vssd1 vssd1 vccd1 vccd1 net3538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1905 _01581_ vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1916 _04393_ vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
X_19838_ net40 _03473_ _03035_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__o21ai_2
Xhold1927 _01330_ vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 _04338_ vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1949 net5829 vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 i_debug_map_overlay vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_19769_ _03000_ _03427_ net1872 _03424_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21800_ clknet_leaf_12_i_clk net3160 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21731_ clknet_leaf_21_i_clk net1550 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21662_ clknet_leaf_35_i_clk net5430 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20613_ net3930 _05196_ net3937 vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__or3b_1
XFILLER_0_188_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21593_ clknet_leaf_24_i_clk net5760 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20544_ _03902_ net3647 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20475_ net3424 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5210 _00677_ vssd1 vssd1 vccd1 vccd1 net5734 sky130_fd_sc_hd__dlygate4sd3_1
X_22214_ net346 net1899 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5221 rbzero.wall_tracer.mapX\[9\] vssd1 vssd1 vccd1 vccd1 net5745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5232 _00815_ vssd1 vssd1 vccd1 vccd1 net5756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5243 rbzero.tex_b0\[1\] vssd1 vssd1 vccd1 vccd1 net5767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5254 rbzero.pov.spi_buffer\[56\] vssd1 vssd1 vccd1 vccd1 net5778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4520 rbzero.spi_registers.buf_othery\[3\] vssd1 vssd1 vccd1 vccd1 net5044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5265 _00707_ vssd1 vssd1 vccd1 vccd1 net5789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4531 net778 vssd1 vssd1 vccd1 vccd1 net5055 sky130_fd_sc_hd__dlygate4sd3_1
X_22145_ net277 net2546 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
Xhold5276 net1763 vssd1 vssd1 vccd1 vccd1 net5800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5287 net1992 vssd1 vssd1 vccd1 vccd1 net5811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4542 _00843_ vssd1 vssd1 vccd1 vccd1 net5066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5298 _04197_ vssd1 vssd1 vccd1 vccd1 net5822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4553 _00727_ vssd1 vssd1 vccd1 vccd1 net5077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4564 _00853_ vssd1 vssd1 vccd1 vccd1 net5088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4575 net817 vssd1 vssd1 vccd1 vccd1 net5099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3830 _08118_ vssd1 vssd1 vccd1 vccd1 net4354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3841 _00986_ vssd1 vssd1 vccd1 vccd1 net4365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4586 net821 vssd1 vssd1 vccd1 vccd1 net5110 sky130_fd_sc_hd__dlygate4sd3_1
X_22076_ clknet_leaf_9_i_clk net3386 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3852 net1422 vssd1 vssd1 vccd1 vccd1 net4376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4597 net603 vssd1 vssd1 vccd1 vccd1 net5121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3863 rbzero.debug_overlay.playerY\[2\] vssd1 vssd1 vccd1 vccd1 net4387 sky130_fd_sc_hd__buf_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03993_ clknet_0__03993_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03993_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3874 net7594 vssd1 vssd1 vccd1 vccd1 net4398 sky130_fd_sc_hd__dlygate4sd3_1
X_21027_ net890 net5334 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nand2_1
Xhold3885 net928 vssd1 vssd1 vccd1 vccd1 net4409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3896 _01002_ vssd1 vssd1 vccd1 vccd1 net4420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ net52 _05957_ _05958_ net51 vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a22o_1
X_13780_ net79 vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__buf_2
X_10992_ net2876 net6527 _04366_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ reg_gpout\[1\] clknet_1_1__leaf__05891_ _05204_ vssd1 vssd1 vccd1 vccd1 _05892_
+ sky130_fd_sc_hd__mux2_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21929_ clknet_leaf_8_i_clk net1254 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15450_ _08511_ _08524_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__or2b_1
XFILLER_0_210_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ net6287 vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__buf_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ _07531_ _07540_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__xor2_2
XFILLER_0_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ rbzero.spi_registers.texadd3\[4\] _04640_ _04642_ rbzero.spi_registers.texadd2\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a22o_1
X_15381_ _08455_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__clkbuf_4
X_12593_ _04983_ _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17120_ _09847_ _10094_ _10121_ vssd1 vssd1 vccd1 vccd1 _10122_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ _07481_ _07482_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__and2_1
X_11544_ _04699_ _04700_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17051_ _10056_ net3462 net4903 vssd1 vssd1 vccd1 vccd1 _10057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14263_ _07369_ _07410_ _07413_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__a21o_1
X_11475_ rbzero.spi_registers.texadd3\[12\] rbzero.spi_registers.texadd1\[12\] rbzero.spi_registers.texadd0\[12\]
+ rbzero.spi_registers.texadd2\[12\] _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04647_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _09076_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__inv_2
X_13214_ net4896 _06186_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__xnor2_1
X_20301__37 clknet_1_1__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
X_14194_ _07343_ _07344_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ net3501 vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _01778_ _08793_ _02000_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__or3_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ net3880 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12027_ net3989 _04803_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__or2b_1
X_16904_ net5471 _09939_ _09940_ net3356 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17884_ _01932_ _01933_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19623_ net5061 net799 _03348_ _03343_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__o211a_1
X_16835_ _09901_ _09903_ vssd1 vssd1 vccd1 vccd1 _09905_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19554_ net3088 _03305_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__or2_1
X_16766_ _08717_ _08588_ _08556_ _08317_ vssd1 vssd1 vccd1 vccd1 _09836_ sky130_fd_sc_hd__o22a_1
X_13978_ _06876_ _06970_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ net3214 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__clkbuf_1
X_15717_ _08778_ _08784_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__or2b_1
X_12929_ _06085_ _06052_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__or2b_1
X_16697_ _09653_ _09767_ vssd1 vssd1 vccd1 vccd1 _09768_ sky130_fd_sc_hd__xor2_4
X_19485_ _02491_ _02500_ _03238_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__and3_2
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18436_ _02452_ _02455_ _02453_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__o21a_1
X_15648_ _08687_ _08693_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__nand2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15579_ _08639_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__xnor2_2
X_18367_ _02401_ _02402_ _10072_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17318_ _10316_ _10318_ vssd1 vssd1 vccd1 vccd1 _10319_ sky130_fd_sc_hd__xor2_2
XFILLER_0_161_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _02340_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17249_ _10221_ _10222_ _10249_ vssd1 vssd1 vccd1 vccd1 _10250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03987_ _03987_ vssd1 vssd1 vccd1 vccd1 clknet_0__03987_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20260_ net3476 _03756_ _03758_ _03748_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20905__319 clknet_1_0__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__inv_2
XFILLER_0_122_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20191_ net3782 _03717_ _03719_ _03709_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3104 net6149 vssd1 vssd1 vccd1 vccd1 net3628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3115 _01182_ vssd1 vssd1 vccd1 vccd1 net3639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3126 net5617 vssd1 vssd1 vccd1 vccd1 net3650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3137 _03810_ vssd1 vssd1 vccd1 vccd1 net3661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3148 _03930_ vssd1 vssd1 vccd1 vccd1 net3672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2403 rbzero.pov.ready_buffer\[65\] vssd1 vssd1 vccd1 vccd1 net2927 sky130_fd_sc_hd__buf_1
Xhold3159 net5530 vssd1 vssd1 vccd1 vccd1 net3683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2414 _03660_ vssd1 vssd1 vccd1 vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2425 _03025_ vssd1 vssd1 vccd1 vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2436 _08244_ vssd1 vssd1 vccd1 vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1702 _01566_ vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2447 _03020_ vssd1 vssd1 vccd1 vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1713 net7027 vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2458 net6167 vssd1 vssd1 vccd1 vccd1 net2982 sky130_fd_sc_hd__clkbuf_2
Xhold1724 _01444_ vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2469 net6022 vssd1 vssd1 vccd1 vccd1 net2993 sky130_fd_sc_hd__clkbuf_2
Xhold1735 net2698 vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1746 _01126_ vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1757 net4269 vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1768 net7114 vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1779 _01389_ vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ clknet_leaf_25_i_clk net2276 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21645_ clknet_leaf_34_i_clk net6273 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21576_ clknet_leaf_4_i_clk net5055 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_50 net3772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_72 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_83 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20527_ net2914 net3435 _03889_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_94 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ net6864 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20458_ _03836_ net3834 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__and2_1
Xhold5040 net1124 vssd1 vssd1 vccd1 vccd1 net5564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5051 net1389 vssd1 vssd1 vccd1 vccd1 net5575 sky130_fd_sc_hd__dlygate4sd3_1
X_20845__266 clknet_1_0__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__inv_2
Xhold5062 _01051_ vssd1 vssd1 vccd1 vccd1 net5586 sky130_fd_sc_hd__dlygate4sd3_1
X_11191_ net6389 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5073 rbzero.pov.mosi vssd1 vssd1 vccd1 vccd1 net5597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20389_ net3250 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__buf_4
Xhold5084 rbzero.spi_registers.texadd0\[4\] vssd1 vssd1 vccd1 vccd1 net5608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4350 net6158 vssd1 vssd1 vccd1 vccd1 net4874 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5095 net1296 vssd1 vssd1 vccd1 vccd1 net5619 sky130_fd_sc_hd__dlygate4sd3_1
X_22128_ net260 net2510 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold4361 _01106_ vssd1 vssd1 vccd1 vccd1 net4885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4372 net6288 vssd1 vssd1 vccd1 vccd1 net4896 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_207_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4383 net864 vssd1 vssd1 vccd1 vccd1 net4907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4394 _06389_ vssd1 vssd1 vccd1 vccd1 net4918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3660 net7448 vssd1 vssd1 vccd1 vccd1 net4184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3671 _00777_ vssd1 vssd1 vccd1 vccd1 net4195 sky130_fd_sc_hd__dlygate4sd3_1
X_14950_ _08088_ _08091_ _08095_ _08068_ net6162 vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__a221o_2
X_22059_ clknet_leaf_10_i_clk net3363 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3682 _00770_ vssd1 vssd1 vccd1 vccd1 net4206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3693 net795 vssd1 vssd1 vccd1 vccd1 net4217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2970 net4527 vssd1 vssd1 vccd1 vccd1 net3494 sky130_fd_sc_hd__dlygate4sd3_1
X_13901_ _07045_ _07046_ _07050_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a21oi_1
X_14881_ net7908 _07986_ _07988_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__and3_2
Xhold2981 net3392 vssd1 vssd1 vccd1 vccd1 net3505 sky130_fd_sc_hd__buf_1
Xhold2992 _03934_ vssd1 vssd1 vccd1 vccd1 net3516 sky130_fd_sc_hd__dlygate4sd3_1
X_16620_ _09658_ _09690_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__xnor2_4
X_13832_ _06873_ _06982_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ _09475_ _09501_ _09622_ vssd1 vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__a21boi_1
X_13763_ _06860_ _06864_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__xor2_1
X_10975_ net2357 net6856 _04355_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _04646_ _08336_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__nand2_1
X_12714_ _05872_ _05874_ net13 vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__mux2_1
X_16482_ _09327_ _09331_ _09431_ vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__a21o_1
X_19270_ net4607 _03133_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13694_ net3132 _06837_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__a21bo_1
X_15433_ _08500_ _08506_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__nand2_1
X_18221_ net4575 _02265_ _01870_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a21o_1
X_12645_ net51 _05795_ _05799_ net52 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18152_ _02197_ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__nand2_1
X_15364_ net3008 _08418_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ rbzero.tex_b1\[27\] rbzero.tex_b1\[26\] _04989_ vssd1 vssd1 vccd1 vccd1 _05741_
+ sky130_fd_sc_hd__mux2_1
X_17103_ _08310_ net7378 vssd1 vssd1 vccd1 vccd1 _10105_ sky130_fd_sc_hd__and2_1
X_14315_ _07405_ _07437_ _07462_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__a21oi_2
X_18083_ _01778_ _09249_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nor2_1
X_11527_ _04696_ _04697_ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15295_ _08117_ net7810 _08294_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17034_ _10032_ _10033_ _10034_ vssd1 vssd1 vccd1 vccd1 _10041_ sky130_fd_sc_hd__o21a_1
X_14246_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__and2_2
Xhold309 net5094 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14177_ _06895_ _06867_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__or2_1
X_11389_ net6978 net6732 _04573_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ net3327 _06283_ net3447 _06281_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__a2bb2o_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ net3854 net4874 net4902 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17936_ _01906_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__and3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ net3620 _04899_ net4874 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__a21o_1
Xhold1009 net6231 vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17867_ _01778_ _08705_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19606_ net5391 _03325_ _03338_ _03330_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16818_ _09885_ _09886_ _09860_ vssd1 vssd1 vccd1 vccd1 _09888_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _01798_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19537_ net1727 _03289_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__or2_1
X_16749_ _09817_ _09818_ vssd1 vssd1 vccd1 vccd1 _09819_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20349__81 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19468_ net1607 net2973 net3077 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ _02440_ _02441_ _02438_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19399_ net1686 _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21430_ clknet_leaf_81_i_clk net4554 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21361_ clknet_leaf_56_i_clk _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold810 _01358_ vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21292_ clknet_leaf_75_i_clk net4085 vssd1 vssd1 vccd1 vccd1 reg_rgb\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold821 net5641 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 net4841 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 net4774 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
X_20243_ net3800 _03744_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2_1
Xhold854 net5615 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 net5574 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 net5664 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 net3495 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_20982__9 clknet_1_0__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
Xhold898 net7901 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
X_20174_ net5517 _03705_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or2_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2200 _04238_ vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2211 net7138 vssd1 vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2222 rbzero.tex_g1\[63\] vssd1 vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2233 _04253_ vssd1 vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
X_20985__12 clknet_1_1__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_72_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 net5705 vssd1 vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__buf_1
Xhold1510 net1929 vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2255 _04211_ vssd1 vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1521 net7033 vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2266 net5979 vssd1 vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2277 _01161_ vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1532 _01483_ vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 net6819 vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2288 net7310 vssd1 vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1554 _00879_ vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2299 net5992 vssd1 vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_212_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1565 _00907_ vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1576 rbzero.tex_r0\[59\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1587 net6917 vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1598 net4883 vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ net7121 net7060 _04244_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10691_ net6942 net7209 _04203_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12430_ rbzero.tex_g1\[23\] rbzero.tex_g1\[22\] _04987_ vssd1 vssd1 vccd1 vccd1 _05597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21628_ clknet_leaf_2_i_clk net5289 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12361_ _04842_ _05528_ _04858_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21559_ clknet_leaf_19_i_clk net920 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14100_ _07231_ _07249_ _07250_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__o21bai_4
X_11312_ net7270 net6742 _04540_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__mux2_1
X_15080_ _08190_ _08203_ net6092 _01622_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12292_ _05229_ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14031_ _07179_ _07180_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__and2_1
X_11243_ net6926 net7251 _04503_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
X_11174_ net6766 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
Xhold4180 rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 net4704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4191 net7606 vssd1 vssd1 vccd1 vccd1 net4715 sky130_fd_sc_hd__dlygate4sd3_1
X_18770_ _02765_ _08195_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15982_ _08347_ _08367_ _08455_ _08492_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__or4_1
XFILLER_0_140_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3490 _04889_ vssd1 vssd1 vccd1 vccd1 net4014 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17721_ _01770_ _01771_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__or2_1
X_14933_ _08077_ _08079_ _06589_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17652_ _09582_ _10407_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14864_ _08006_ _08014_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__nand2_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16603_ _08454_ _09311_ vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__or2_1
X_13815_ _06893_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__buf_6
XFILLER_0_212_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17583_ _10502_ _10579_ _10580_ vssd1 vssd1 vccd1 vccd1 _10581_ sky130_fd_sc_hd__a21oi_2
X_14795_ _07936_ _07942_ _07945_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19322_ net1729 _03160_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ _06895_ net547 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__nor2_1
X_16534_ _08180_ net77 _09605_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__a21oi_2
X_10958_ _04332_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19253_ net4149 _03119_ net610 _03128_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16465_ _09304_ _09536_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__or2_2
X_13677_ _06606_ _06608_ _06727_ _06619_ _06692_ _06688_ vssd1 vssd1 vccd1 vccd1 _06828_
+ sky130_fd_sc_hd__mux4_1
X_10889_ net6990 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__05891_ clknet_0__05891_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05891_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18204_ _02174_ _02175_ _02249_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__and3_1
X_15416_ net3470 _06209_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12628_ net7 vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__inv_2
X_16396_ _09467_ _09468_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__xnor2_1
X_19184_ net2964 net7322 _03084_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18135_ _10259_ _09863_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15347_ _08307_ _08416_ _08417_ _08421_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__a2bb2o_4
X_12559_ _04983_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5809 net728 vssd1 vssd1 vccd1 vccd1 net6333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15278_ net3397 _06209_ _08351_ _08352_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__a2bb2o_4
X_18066_ _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__xor2_1
Xhold106 net823 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold117 net4676 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
X_20828__250 clknet_1_0__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__inv_2
Xhold128 rbzero.wall_tracer.visualWallDist\[5\] vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17017_ _10014_ _10015_ _10016_ vssd1 vssd1 vccd1 vccd1 _10026_ sky130_fd_sc_hd__o21ai_2
X_14229_ _07376_ _07379_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__xnor2_1
Xhold139 net4960 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _06217_ _09950_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__or2_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _01741_ _01744_ _01859_ _01968_ _01858_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__o311a_4
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _02854_ net4459 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22462_ clknet_leaf_39_i_clk _01631_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21413_ clknet_leaf_84_i_clk net3596 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22393_ net525 net590 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21344_ clknet_leaf_56_i_clk net4526 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold640 net5503 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21275_ clknet_leaf_72_i_clk _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold651 net3475 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 net5560 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 net6430 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
X_20226_ net1270 _03731_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__or2_1
Xhold684 _01422_ vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold695 net4212 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20157_ net1162 _03692_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2030 net6276 vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2041 net2577 vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2052 _01579_ vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2063 net7106 vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2074 _01304_ vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ net3225 _03653_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__or2_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2085 _04581_ vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1340 net4323 vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2096 _04563_ vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 net5891 vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net4254 net4280 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__nand2_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 net7655 vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_197_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1373 net6801 vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1384 _01170_ vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 _01350_ vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11861_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _04989_ vssd1 vssd1 vccd1 vccd1 _05031_
+ sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06662_ _06741_ _06750_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__o21a_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ net6409 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _07721_ _07730_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__xor2_2
XFILLER_0_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _04926_ _04960_ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ _06530_ _06543_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__nor2_1
X_20328__62 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
X_10743_ net6455 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16250_ _09192_ _09201_ _09199_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13462_ _06612_ _06557_ _06564_ _06587_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__or4bb_4
X_10674_ net2569 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15201_ _08279_ net4083 vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__and2_1
X_12413_ _05261_ _05579_ _05244_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__o21a_1
X_20343__76 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
X_16181_ _08726_ _08728_ _09255_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13393_ _06531_ _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__or2_4
XFILLER_0_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ net6134 _08223_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12344_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _04986_ vssd1 vssd1 vccd1 vccd1 _05512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15063_ net4568 net4475 _08191_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19940_ net3360 _03480_ _03532_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ _04816_ _05441_ _05443_ net4043 _05201_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a311oi_1
X_14014_ _07163_ _07164_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__nand2_1
X_11226_ net5865 net5872 _04492_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__mux2_1
X_19871_ net4219 _03479_ net1014 _03502_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__a211o_1
X_18822_ net4634 rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02813_
+ sky130_fd_sc_hd__nand2_1
X_11157_ net5848 net6547 _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18753_ net3035 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15965_ _09028_ _09027_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__and2b_1
X_11088_ net2314 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
X_17704_ _01753_ _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14916_ _06690_ _07993_ _08029_ _07995_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__a211o_1
X_18684_ _02662_ _02663_ _02688_ net4810 net4767 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a311o_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _08422_ _08501_ vssd1 vssd1 vccd1 vccd1 _08971_ sky130_fd_sc_hd__nor2_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ _08717_ _09595_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14847_ _07584_ _07978_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ _10340_ _10564_ vssd1 vssd1 vccd1 vccd1 _10565_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14778_ _07924_ _07927_ _07928_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_147_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ _03036_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__clkbuf_4
X_16517_ _08684_ _08574_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13729_ _06844_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17497_ _10486_ _10495_ vssd1 vssd1 vccd1 vccd1 _10496_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19236_ _03039_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__buf_2
X_16448_ _09518_ _09520_ vssd1 vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__xor2_4
Xhold7008 net4486 vssd1 vssd1 vccd1 vccd1 net7532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7019 rbzero.wall_tracer.trackDistY\[-5\] vssd1 vssd1 vccd1 vccd1 net7543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6307 rbzero.tex_b0\[29\] vssd1 vssd1 vccd1 vccd1 net6831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19167_ net5710 _03065_ _03077_ _03074_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6318 net2200 vssd1 vssd1 vccd1 vccd1 net6842 sky130_fd_sc_hd__dlygate4sd3_1
X_16379_ _08564_ _08471_ _08516_ _08565_ vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__or4_1
XFILLER_0_182_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6329 rbzero.spi_registers.buf_texadd1\[2\] vssd1 vssd1 vccd1 vccd1 net6853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18118_ _02164_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5606 net3008 vssd1 vssd1 vccd1 vccd1 net6130 sky130_fd_sc_hd__dlygate4sd3_1
X_19098_ _04881_ _05816_ _03032_ _03033_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__nand4_4
Xhold5617 _02964_ vssd1 vssd1 vccd1 vccd1 net6141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5639 rbzero.spi_registers.spi_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net6163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4905 _00831_ vssd1 vssd1 vccd1 vccd1 net5429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18049_ _08705_ _09375_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4916 _01076_ vssd1 vssd1 vccd1 vccd1 net5440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4927 rbzero.spi_registers.texadd0\[18\] vssd1 vssd1 vccd1 vccd1 net5451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4938 net8009 vssd1 vssd1 vccd1 vccd1 net5462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4949 net986 vssd1 vssd1 vccd1 vccd1 net5473 sky130_fd_sc_hd__dlygate4sd3_1
X_21060_ net4736 _03519_ _04014_ _04057_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20011_ net3745 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21962_ net187 net2713 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20913_ clknet_1_1__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__buf_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21893_ clknet_leaf_95_i_clk net1336 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22445_ clknet_leaf_51_i_clk net3982 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6830 rbzero.spi_registers.spi_counter\[1\] vssd1 vssd1 vccd1 vccd1 net7354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22376_ net508 net1749 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__04012_ clknet_0__04012_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04012_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6841 rbzero.color_floor\[3\] vssd1 vssd1 vccd1 vccd1 net7365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6852 _10578_ vssd1 vssd1 vccd1 vccd1 net7376 sky130_fd_sc_hd__dlygate4sd3_1
X_21327_ clknet_leaf_36_i_clk net4305 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ _04982_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__buf_4
Xhold470 net5372 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
X_21258_ clknet_leaf_71_i_clk net3632 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold481 net5354 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net5831 net5879 _04377_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__mux2_1
Xhold492 net5454 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
X_20209_ net5646 _03718_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__or2_1
X_21189_ net4806 _02528_ _02579_ _04146_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _08808_ _08822_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__nor2_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _06105_ _06114_ _06113_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 _00890_ vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _05081_ _05082_ _04992_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__mux2_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _07817_ _07830_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__xnor2_1
Xhold1181 _00877_ vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 net6657 vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _08754_ _08631_ _08755_ _08540_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__a22o_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ net4095 _05446_ _06046_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17420_ _10417_ _10418_ _10419_ vssd1 vssd1 vccd1 vccd1 _10420_ sky130_fd_sc_hd__nand3_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _04987_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__clkbuf_8
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _07768_ _07781_ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__a21boi_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _10349_ _10350_ vssd1 vssd1 vccd1 vccd1 _10351_ sky130_fd_sc_hd__nor2_1
X_14563_ _07702_ _07711_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__a21oi_4
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _04940_ _04943_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ net7444 _09375_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__nor2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ net6870 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__clkbuf_1
X_13514_ _06588_ _06597_ _06610_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__and3_1
X_17282_ _10162_ _10165_ _10282_ vssd1 vssd1 vccd1 vccd1 _10283_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14494_ _07356_ _07304_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19021_ net2842 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__buf_2
X_16233_ _09252_ _09133_ _09306_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__and3b_1
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13445_ _06591_ _06595_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ net2299 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20710__144 clknet_1_0__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__inv_2
XFILLER_0_181_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16164_ _08639_ _08653_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ net4947 _06523_ _06524_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__a31o_2
XFILLER_0_134_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ _05492_ _05494_ _04992_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15115_ net4501 net4613 _08219_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__mux2_1
X_16095_ _09078_ _09079_ _09120_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19923_ net4294 _03530_ net2991 _03496_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__o211a_1
X_15046_ _08157_ _08176_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12258_ rbzero.debug_overlay.playerY\[2\] _05369_ _05384_ rbzero.debug_overlay.playerY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a22o_1
X_11209_ net6421 net7107 _04481_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
X_19854_ _03479_ net3031 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__or2_1
X_12189_ _05339_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18805_ net3699 rbzero.wall_tracer.rayAddendY\[-2\] _02789_ vssd1 vssd1 vccd1 vccd1
+ _02797_ sky130_fd_sc_hd__o21a_1
X_19785_ net5838 _03442_ net648 _03441_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__o211a_1
X_16997_ _10006_ _10007_ vssd1 vssd1 vccd1 vccd1 _10008_ sky130_fd_sc_hd__or2b_1
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18736_ _01870_ _06192_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__nor2_1
X_15948_ _08432_ _08626_ _09021_ _09022_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__o31a_1
X_18667_ net4696 _02666_ _02673_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a21o_1
X_15879_ _08559_ _08411_ _08432_ _08367_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _01668_ _01669_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18598_ net6237 _05403_ _02607_ _02608_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__04006_ _04006_ vssd1 vssd1 vccd1 vccd1 clknet_0__04006_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17549_ _10538_ _10547_ vssd1 vssd1 vccd1 vccd1 _10548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20560_ _03902_ net3259 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__and2_1
X_20307__43 clknet_1_0__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_0_117_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19219_ net5852 _03106_ _03110_ _03096_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__o211a_1
Xhold6104 net1892 vssd1 vssd1 vccd1 vccd1 net6628 sky130_fd_sc_hd__dlygate4sd3_1
X_20491_ net3532 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__clkbuf_1
Xhold6115 rbzero.tex_g0\[13\] vssd1 vssd1 vccd1 vccd1 net6639 sky130_fd_sc_hd__dlygate4sd3_1
X_22230_ net362 net2327 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold6126 net1718 vssd1 vssd1 vccd1 vccd1 net6650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6137 rbzero.spi_registers.buf_texadd2\[4\] vssd1 vssd1 vccd1 vccd1 net6661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5403 net5975 vssd1 vssd1 vccd1 vccd1 net5927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6148 net1851 vssd1 vssd1 vccd1 vccd1 net6672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5414 rbzero.map_overlay.i_mapdy\[4\] vssd1 vssd1 vccd1 vccd1 net5938 sky130_fd_sc_hd__dlygate4sd3_1
X_20685__121 clknet_1_0__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__inv_2
Xhold6159 rbzero.tex_g0\[55\] vssd1 vssd1 vccd1 vccd1 net6683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5425 rbzero.map_overlay.i_mapdx\[2\] vssd1 vssd1 vccd1 vccd1 net5949 sky130_fd_sc_hd__dlygate4sd3_1
X_22161_ net293 net2451 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5436 _00662_ vssd1 vssd1 vccd1 vccd1 net5960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4702 net886 vssd1 vssd1 vccd1 vccd1 net5226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5447 net2612 vssd1 vssd1 vccd1 vccd1 net5971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5458 _04209_ vssd1 vssd1 vccd1 vccd1 net5982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4713 _00856_ vssd1 vssd1 vccd1 vccd1 net5237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4724 _00830_ vssd1 vssd1 vccd1 vccd1 net5248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5469 net2823 vssd1 vssd1 vccd1 vccd1 net5993 sky130_fd_sc_hd__dlygate4sd3_1
X_21112_ _04099_ _04100_ _04098_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__o21ai_1
Xhold4735 net900 vssd1 vssd1 vccd1 vccd1 net5259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4746 rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 net5270 sky130_fd_sc_hd__dlygate4sd3_1
X_22092_ clknet_leaf_49_i_clk net4003 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4757 net974 vssd1 vssd1 vccd1 vccd1 net5281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4768 _00800_ vssd1 vssd1 vccd1 vccd1 net5292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4779 _00834_ vssd1 vssd1 vccd1 vccd1 net5303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21043_ _04038_ _04039_ _04040_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o21a_1
XFILLER_0_201_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_199_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21945_ net170 net2795 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ clknet_leaf_98_i_clk net1246 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _04724_ _04696_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20758_ clknet_1_0__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__buf_1
XFILLER_0_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11491_ _04660_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13230_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22428_ clknet_leaf_46_i_clk net4738 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7383 net4331 vssd1 vssd1 vccd1 vccd1 net7907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7394 rbzero.wall_tracer.stepDistY\[7\] vssd1 vssd1 vccd1 vccd1 net7918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6660 rbzero.tex_b0\[16\] vssd1 vssd1 vccd1 vccd1 net7184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ _06314_ net3174 _06316_ net3460 vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a2bb2o_1
X_22359_ net491 net2384 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6671 net2487 vssd1 vssd1 vccd1 vccd1 net7195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6682 rbzero.tex_r0\[40\] vssd1 vssd1 vccd1 vccd1 net7206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6693 net2665 vssd1 vssd1 vccd1 vccd1 net7217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ rbzero.tex_r1\[23\] rbzero.tex_r1\[22\] _05218_ vssd1 vssd1 vccd1 vccd1 _05281_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5970 _04493_ vssd1 vssd1 vccd1 vccd1 net6494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13092_ net3265 vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__inv_2
Xhold5981 rbzero.tex_b0\[60\] vssd1 vssd1 vccd1 vccd1 net6505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5992 net1464 vssd1 vssd1 vccd1 vccd1 net6516 sky130_fd_sc_hd__dlygate4sd3_1
X_16920_ net4133 _09941_ _09942_ net7442 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a22o_1
X_12043_ net4254 _05051_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21o_1
X_16851_ _04160_ _09919_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ _08518_ _08876_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19570_ net5186 _03302_ _03317_ _03314_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__o211a_1
X_16782_ _08899_ _08599_ _09721_ _09851_ vssd1 vssd1 vccd1 vccd1 _09852_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13994_ _07141_ _07143_ _07144_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a21oi_2
X_18521_ net4476 net908 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__nand2_1
X_15733_ _08760_ _08765_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__xnor2_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _06099_
+ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__a31o_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ net3059 _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__nand2_1
X_15664_ _08735_ _08737_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__and2_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _06025_ _06033_ net30 vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _10285_ _10287_ _10284_ vssd1 vssd1 vccd1 vccd1 _10403_ sky130_fd_sc_hd__a21bo_1
X_14615_ _07763_ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__nor2_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11827_ _04956_ _04944_ _04953_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__nor3_1
X_18383_ _09987_ _02415_ net3235 _10206_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a31o_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _08657_ _08659_ _08669_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__a21o_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ net3474 net4349 vssd1 vssd1 vccd1 vccd1 _10334_ sky130_fd_sc_hd__or2_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _04925_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__nand2_1
X_14546_ _06957_ _06955_ _07399_ _07438_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__or4_4
XFILLER_0_154_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ net2703 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17265_ _08872_ _09477_ vssd1 vssd1 vccd1 vccd1 _10266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14477_ _07620_ _07627_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__xor2_4
X_11689_ _04842_ net4064 _04849_ _04851_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a41o_1
XFILLER_0_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19004_ net3915 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16216_ _09283_ _09289_ _09290_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13428_ _06569_ _06571_ _06578_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17196_ _10092_ _10197_ vssd1 vssd1 vccd1 vccd1 _10198_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ net3170 _08313_ _08630_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13359_ _06440_ _06509_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__xnor2_2
Xhold4009 _00482_ vssd1 vssd1 vccd1 vccd1 net4533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _09131_ _09151_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__xnor2_1
Xhold3308 _00998_ vssd1 vssd1 vccd1 vccd1 net3832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3319 net1339 vssd1 vssd1 vccd1 vccd1 net3843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19906_ net41 _03473_ _03035_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__o21ai_2
X_15029_ _08092_ _08164_ net7836 vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__a21oi_1
Xhold2607 _00699_ vssd1 vssd1 vccd1 vccd1 net3131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2618 _00991_ vssd1 vssd1 vccd1 vccd1 net3142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _03461_ vssd1 vssd1 vccd1 vccd1 net3153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1906 net6933 vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_19837_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__clkbuf_4
Xhold1917 _01388_ vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1928 net7156 vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 _01438_ vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xinput2 i_debug_trace_overlay vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
X_19768_ net6720 _03429_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18719_ net4787 _02557_ _09943_ _02720_ _02722_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19699_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21730_ clknet_leaf_21_i_clk net1672 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21661_ clknet_leaf_35_i_clk net5249 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20612_ _04777_ net2988 _03953_ _08276_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21592_ clknet_leaf_24_i_clk net5738 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20543_ net747 net3646 _03889_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20474_ _03858_ net3423 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5200 net1557 vssd1 vssd1 vccd1 vccd1 net5724 sky130_fd_sc_hd__dlygate4sd3_1
X_22213_ net345 net1112 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
Xhold5211 rbzero.spi_registers.texadd2\[7\] vssd1 vssd1 vccd1 vccd1 net5735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5222 net2787 vssd1 vssd1 vccd1 vccd1 net5746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5233 rbzero.spi_registers.texadd2\[8\] vssd1 vssd1 vccd1 vccd1 net5757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5244 _04596_ vssd1 vssd1 vccd1 vccd1 net5768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5255 rbzero.spi_registers.vshift\[2\] vssd1 vssd1 vccd1 vccd1 net5779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4510 net781 vssd1 vssd1 vccd1 vccd1 net5034 sky130_fd_sc_hd__dlygate4sd3_1
X_22144_ net276 net2202 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
Xhold5266 rbzero.pov.spi_buffer\[57\] vssd1 vssd1 vccd1 vccd1 net5790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4521 net786 vssd1 vssd1 vccd1 vccd1 net5045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5277 rbzero.spi_registers.vshift\[5\] vssd1 vssd1 vccd1 vccd1 net5801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4532 rbzero.spi_registers.buf_texadd0\[4\] vssd1 vssd1 vccd1 vccd1 net5056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5288 _04199_ vssd1 vssd1 vccd1 vccd1 net5812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4543 rbzero.color_sky\[3\] vssd1 vssd1 vccd1 vccd1 net5067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4554 rbzero.spi_registers.buf_mapdy\[5\] vssd1 vssd1 vccd1 vccd1 net5078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5299 net589 vssd1 vssd1 vccd1 vccd1 net5823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3820 net3040 vssd1 vssd1 vccd1 vccd1 net4344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4565 net838 vssd1 vssd1 vccd1 vccd1 net5089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3831 net7999 vssd1 vssd1 vccd1 vccd1 net4355 sky130_fd_sc_hd__buf_2
X_22075_ clknet_leaf_13_i_clk net3499 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4576 _00842_ vssd1 vssd1 vccd1 vccd1 net5100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3842 net706 vssd1 vssd1 vccd1 vccd1 net4366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4587 _00823_ vssd1 vssd1 vccd1 vccd1 net5111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3853 net7812 vssd1 vssd1 vccd1 vccd1 net4377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4598 _00864_ vssd1 vssd1 vccd1 vccd1 net5122 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03992_ clknet_0__03992_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03992_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3864 _00981_ vssd1 vssd1 vccd1 vccd1 net4388 sky130_fd_sc_hd__dlygate4sd3_1
X_21026_ net890 net5334 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__nor2_1
Xhold3875 net3149 vssd1 vssd1 vccd1 vccd1 net4399 sky130_fd_sc_hd__buf_1
Xhold3886 net7493 vssd1 vssd1 vccd1 vccd1 net4410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3897 net889 vssd1 vssd1 vccd1 vccd1 net4421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10991_ net1742 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ net4066 _05846_ _05851_ _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__o22a_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21928_ clknet_leaf_6_i_clk net1283 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12661_ net7 net8 _05819_ _05821_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a32o_1
XFILLER_0_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21859_ clknet_leaf_83_i_clk net2901 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _07465_ _07469_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__xor2_2
X_11612_ rbzero.spi_registers.texadd1\[4\] _04644_ _04709_ rbzero.spi_registers.texadd0\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a22o_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12592_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _04994_ vssd1 vssd1 vccd1 vccd1 _05757_
+ sky130_fd_sc_hd__mux2_1
X_15380_ net3332 _06210_ _08454_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_33_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14331_ _07470_ _07480_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__xnor2_1
X_11543_ _04705_ _04712_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17050_ _06206_ net7596 _10055_ vssd1 vssd1 vccd1 vccd1 _10056_ sky130_fd_sc_hd__o21ai_1
X_14262_ _07411_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11474_ net4086 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16001_ _09072_ _09074_ _09075_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13213_ net3984 _06222_ net4874 vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _07288_ _07308_ _07342_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__and3_1
Xhold6490 net2530 vssd1 vssd1 vccd1 vccd1 net7014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ net3381 _06298_ net3555 _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17952_ _01894_ _01895_ _02000_ _01780_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ net3853 _06229_ _06190_ net4387 _06230_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20822__245 clknet_1_0__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__inv_2
X_12026_ net4059 net4033 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__or2_1
X_16903_ net5379 _09939_ _09940_ net3206 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a22o_1
X_17883_ _01911_ _01912_ _01931_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__nand3_1
XFILLER_0_139_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19622_ net1591 _03340_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__or2_1
X_16834_ _09901_ _09903_ vssd1 vssd1 vccd1 vccd1 _09904_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19553_ net5155 _03303_ _03308_ _03295_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__o211a_1
X_16765_ _09834_ vssd1 vssd1 vccd1 vccd1 _09835_ sky130_fd_sc_hd__inv_2
X_13977_ _07121_ _07122_ _07126_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__a21o_1
X_18504_ _02492_ net3213 _02523_ net2978 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__and4bb_1
X_15716_ _08783_ _08781_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__or2b_1
X_19484_ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__clkbuf_2
X_12928_ _05194_ net4060 net3930 net3937 net34 net36 vssd1 vssd1 vccd1 vccd1 _06085_
+ sky130_fd_sc_hd__mux4_1
X_16696_ _09654_ _09766_ vssd1 vssd1 vccd1 vccd1 _09767_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ _02460_ _02461_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__or2b_1
X_15647_ _08710_ _08720_ _08721_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__a21o_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ net43 _05998_ _06007_ net46 vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18366_ net3394 _02398_ _02399_ _06205_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15578_ _08636_ _08640_ _08647_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__a31o_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ _10125_ _10191_ _10317_ vssd1 vssd1 vccd1 vccd1 _10318_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14529_ _07671_ _07678_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__nor2_1
X_18297_ net4467 net4310 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ _10234_ _10248_ vssd1 vssd1 vccd1 vccd1 _10249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03986_ _03986_ vssd1 vssd1 vccd1 vccd1 clknet_0__03986_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17179_ _09868_ _09880_ _09879_ vssd1 vssd1 vccd1 vccd1 _10181_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20190_ net5175 _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3105 _00429_ vssd1 vssd1 vccd1 vccd1 net3629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3116 rbzero.pov.spi_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net3640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3127 net1438 vssd1 vssd1 vccd1 vccd1 net3651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3138 _03811_ vssd1 vssd1 vccd1 vccd1 net3662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2404 _03497_ vssd1 vssd1 vccd1 vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3149 _01241_ vssd1 vssd1 vccd1 vccd1 net3673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 net6177 vssd1 vssd1 vccd1 vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2426 _00651_ vssd1 vssd1 vccd1 vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2437 net4830 vssd1 vssd1 vccd1 vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 net6911 vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _00647_ vssd1 vssd1 vccd1 vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _04418_ vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 _04131_ vssd1 vssd1 vccd1 vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 net7045 vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
X_20797__222 clknet_1_1__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__inv_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1736 _04228_ vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 net7049 vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 net6050 vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 net7116 vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21713_ clknet_leaf_26_i_clk net1606 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21644_ clknet_leaf_27_i_clk net3119 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_40 _10329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21575_ clknet_leaf_4_i_clk net5085 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_51 net4050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 _05177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20526_ net3344 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_73 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_95 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20457_ net3833 net1470 _03845_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5030 net1286 vssd1 vssd1 vccd1 vccd1 net5554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5041 rbzero.pov.spi_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net5565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5052 _01055_ vssd1 vssd1 vccd1 vccd1 net5576 sky130_fd_sc_hd__dlygate4sd3_1
X_11190_ net1372 net6387 _04470_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20388_ net3249 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__buf_1
Xhold5063 rbzero.pov.spi_buffer\[58\] vssd1 vssd1 vccd1 vccd1 net5587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5074 net953 vssd1 vssd1 vccd1 vccd1 net5598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4340 rbzero.pov.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 net4864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5085 net1310 vssd1 vssd1 vccd1 vccd1 net5609 sky130_fd_sc_hd__dlygate4sd3_1
X_22127_ net259 net2187 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold5096 _00627_ vssd1 vssd1 vccd1 vccd1 net5620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4351 _09958_ vssd1 vssd1 vccd1 vccd1 net4875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4362 rbzero.wall_tracer.mapY\[8\] vssd1 vssd1 vccd1 vccd1 net4886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4373 _06227_ vssd1 vssd1 vccd1 vccd1 net4897 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4384 net7353 vssd1 vssd1 vccd1 vccd1 net4908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4395 _06391_ vssd1 vssd1 vccd1 vccd1 net4919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3650 _00509_ vssd1 vssd1 vccd1 vccd1 net4174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3661 net1060 vssd1 vssd1 vccd1 vccd1 net4185 sky130_fd_sc_hd__dlygate4sd3_1
X_22058_ clknet_leaf_7_i_clk net3803 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3672 net1117 vssd1 vssd1 vccd1 vccd1 net4196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3683 net1408 vssd1 vssd1 vccd1 vccd1 net4207 sky130_fd_sc_hd__dlygate4sd3_1
X_21009_ net773 net4987 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__or2_1
X_13900_ _07045_ _07046_ _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__and3_1
Xhold3694 rbzero.debug_overlay.playerX\[-1\] vssd1 vssd1 vccd1 vccd1 net4218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2960 _03912_ vssd1 vssd1 vccd1 vccd1 net3484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2971 net4855 vssd1 vssd1 vccd1 vccd1 net3495 sky130_fd_sc_hd__dlygate4sd3_1
X_14880_ _06690_ _07993_ _08029_ _06678_ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__a211o_1
Xhold2982 net4929 vssd1 vssd1 vccd1 vccd1 net3506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2993 _01243_ vssd1 vssd1 vccd1 vccd1 net3517 sky130_fd_sc_hd__dlygate4sd3_1
X_13831_ _06912_ _06911_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__and2b_1
XFILLER_0_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _09498_ _09500_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__or2b_1
X_10974_ net2639 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__clkbuf_1
X_13762_ _06873_ _06911_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15501_ _08152_ _08575_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__xnor2_2
X_12713_ net3937 _05853_ _05854_ net3930 _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a221o_1
X_16481_ _09543_ _09552_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ _06788_ _06839_ _06843_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__a21o_4
XFILLER_0_183_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18220_ net4575 _02265_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__nor2_1
X_15432_ _08500_ _08506_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ _05790_ net6 _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18151_ _02181_ _02196_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12575_ _05177_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15363_ net6253 _08437_ _08305_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ _10102_ _10103_ vssd1 vssd1 vccd1 vccd1 _10104_ sky130_fd_sc_hd__nor2_1
X_14314_ _07444_ net558 vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__nor2_2
XFILLER_0_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18082_ _02035_ _02036_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ rbzero.spi_registers.texadd3\[20\] rbzero.spi_registers.texadd1\[20\] rbzero.spi_registers.texadd0\[20\]
+ rbzero.spi_registers.texadd2\[20\] _04692_ _04693_ vssd1 vssd1 vccd1 vccd1 _04698_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15294_ net7809 _06497_ net4086 vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _10040_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14245_ _07294_ _07346_ _07394_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__a21o_1
X_11457_ _04621_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ _07270_ _07271_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11388_ net2817 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ net3503 vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ net3853 _02959_ _09999_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17935_ _01906_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a21oi_4
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ net2825 _06213_ net4874 net3620 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12009_ _05177_ _05120_ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__or3b_1
X_17866_ _01914_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16817_ _09860_ _09885_ _09886_ vssd1 vssd1 vccd1 vccd1 _09887_ sky130_fd_sc_hd__nand3_1
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19605_ net3096 _03327_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__or2_1
X_17797_ _01846_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19536_ net5302 _03288_ _03296_ _03295_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__o211a_1
X_16748_ _09811_ _09816_ vssd1 vssd1 vccd1 vccd1 _09818_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19467_ net1572 net3077 net1535 _03233_ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__o211a_1
X_16679_ _09747_ _09749_ vssd1 vssd1 vccd1 vccd1 _09750_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18418_ _02445_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19398_ _03084_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18349_ _02383_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21360_ clknet_leaf_58_i_clk _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20311_ clknet_1_1__leaf__03773_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__buf_1
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold800 net5218 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
X_21291_ clknet_leaf_75_i_clk net4068 vssd1 vssd1 vccd1 vccd1 reg_rgb\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold811 net5480 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 net5643 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold833 net6460 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_20242_ net3800 _03743_ _03747_ _03748_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__o211a_1
Xhold844 net5632 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 net5680 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 net5576 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold877 net5666 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20292__29 clknet_1_1__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
X_20173_ net5517 _03704_ _03708_ _03709_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__o211a_1
Xhold888 _01105_ vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 net4240 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2201 _01525_ vssd1 vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2212 _01122_ vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2223 net2720 vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2234 _01514_ vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1500 net1956 vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 net5707 vssd1 vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 _04527_ vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2256 _01549_ vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1522 _04347_ vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2267 net5946 vssd1 vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__clkbuf_2
Xhold1533 net6987 vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2278 net5917 vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1544 _01571_ vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2289 _03508_ vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 net6897 vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1566 net6169 vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 net1472 vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1588 _01456_ vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1599 _03029_ vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ net2856 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20851__271 clknet_1_1__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__inv_2
XFILLER_0_192_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21627_ clknet_leaf_4_i_clk net5415 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ _05526_ _05527_ net4077 vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__mux2_2
X_21558_ clknet_leaf_20_i_clk net820 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11311_ _04403_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20509_ _03880_ net3574 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__and2_1
X_12291_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _05230_ vssd1 vssd1 vccd1 vccd1 _05459_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21489_ clknet_leaf_15_i_clk net2044 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14030_ _07179_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11242_ net6541 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ net2743 net6764 _04459_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4170 net3407 vssd1 vssd1 vccd1 vccd1 net4694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4181 net2968 vssd1 vssd1 vccd1 vccd1 net4705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4192 net3172 vssd1 vssd1 vccd1 vccd1 net4716 sky130_fd_sc_hd__clkdlybuf4s25_1
X_15981_ _08559_ _08456_ _08493_ _08560_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _10474_ _10586_ _10588_ _10589_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22oi_1
Xhold3480 net7361 vssd1 vssd1 vccd1 vccd1 net4004 sky130_fd_sc_hd__clkbuf_2
X_14932_ net7566 _08078_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__nand2_1
Xhold3491 _03950_ vssd1 vssd1 vccd1 vccd1 net4015 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17651_ _01701_ _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__nand2_1
Xhold2790 net7532 vssd1 vssd1 vccd1 vccd1 net3314 sky130_fd_sc_hd__buf_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _06690_ _08011_ _08013_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__o21ba_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _09564_ _09568_ _09565_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__a21o_1
X_13814_ _06963_ _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__or2_1
XFILLER_0_203_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17582_ _09051_ _09784_ _10483_ _10481_ vssd1 vssd1 vccd1 vccd1 _10580_ sky130_fd_sc_hd__o31a_1
X_14794_ _07943_ _07944_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__nand2_1
X_20934__346 clknet_1_1__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__inv_2
X_19321_ net5314 _03159_ _03167_ _03168_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__o211a_1
X_16533_ _08150_ _08142_ _08183_ _08176_ _08047_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__a221oi_4
X_13745_ net540 _06837_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ net1698 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19252_ net969 _03120_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or2_1
X_16464_ net7442 _08314_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__nand2_2
X_13676_ _06781_ _06796_ _06806_ net562 _06826_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__a2111o_1
X_10888_ net2781 net6988 _04236_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18203_ _02174_ _02175_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a21oi_1
X_15415_ _08299_ _08488_ _08489_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__a21o_4
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19183_ _04597_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__buf_2
X_12627_ net4045 net4066 net4083 net4078 net4 net7 vssd1 vssd1 vccd1 vccd1 _05789_
+ sky130_fd_sc_hd__mux4_1
X_16395_ _08449_ _08582_ vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18134_ _02023_ _02083_ _02091_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ net7404 _08420_ _08306_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__o21a_1
X_12558_ rbzero.tex_b1\[35\] rbzero.tex_b1\[34\] _04994_ vssd1 vssd1 vccd1 vccd1 _05723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18065_ _02031_ _02052_ _02029_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11509_ _04645_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ net3392 _08305_ _08307_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_124_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12489_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _05263_ vssd1 vssd1 vccd1 vccd1 _05655_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 _03058_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 net6103 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_1
XFILLER_0_106_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold129 net4144 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ net4597 net4370 vssd1 vssd1 vccd1 vccd1 _10025_ sky130_fd_sc_hd__nand2_1
X_14228_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14159_ _07266_ _07272_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ net3823 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__clkbuf_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _01756_ _01757_ _01856_ _01738_ _01736_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a311o_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18898_ _02851_ _02869_ _02844_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_206_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ _01897_ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19519_ net5045 _03274_ _03285_ _03280_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__o211a_1
X_20791_ clknet_1_0__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__buf_1
XFILLER_0_147_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22461_ clknet_leaf_38_i_clk _01630_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21412_ clknet_leaf_84_i_clk net4694 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22392_ net524 net1764 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21343_ clknet_leaf_56_i_clk net4287 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold630 net6408 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21274_ clknet_leaf_51_i_clk _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold641 net5505 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold652 net4854 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20225_ net5240 _03730_ _03738_ _03735_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__o211a_1
Xhold663 net4860 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _01149_ vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 net4832 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
X_20881__297 clknet_1_1__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__inv_2
XFILLER_0_200_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold696 net3382 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20156_ net5585 _03691_ _03699_ _03696_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__o211a_1
Xhold2020 net7214 vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 net6277 vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2042 _04464_ vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2053 rbzero.tex_b1\[57\] vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20087_ net4794 net2122 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__and2b_1
Xhold2064 _04487_ vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2075 net7128 vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 net6689 vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 net6981 vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2086 _01124_ vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2097 _01141_ vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 _01269_ vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1363 net4939 vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1374 _04398_ vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 net6567 vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1396 net6554 vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _05022_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__clkbuf_8
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ net6407 net2445 _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11791_ _04923_ _04925_ _04922_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a21oi_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _06588_ _06644_ _06630_ _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__a211o_1
X_10742_ net6453 net2753 _04236_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10673_ net7056 net7141 _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__mux2_1
X_13461_ _06561_ _06566_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ net4067 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
X_12412_ rbzero.tex_g1\[3\] rbzero.tex_g1\[2\] _05476_ vssd1 vssd1 vccd1 vccd1 _05579_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16180_ _09253_ _09254_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13392_ _06538_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15131_ net4497 net4437 _08219_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__mux2_1
X_12343_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _05493_ vssd1 vssd1 vccd1 vccd1 _05511_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12274_ _05342_ _05197_ _05333_ net85 vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__nand4_1
X_15062_ _06344_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11225_ net2186 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
X_14013_ _07162_ _07157_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19870_ _04597_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11156_ _04332_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__clkbuf_4
X_18821_ net4634 rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18752_ _02748_ net6309 _06392_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
X_15964_ _09009_ _09038_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__xnor2_2
X_11087_ net6924 net6914 _04415_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17703_ net7375 _10577_ net7374 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__o21a_1
X_14915_ _08006_ _08035_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18683_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] _02637_
+ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__o21a_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _08969_ _08490_ _08491_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__and3_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858__277 clknet_1_0__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__inv_2
X_17634_ _01683_ _01685_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__and2_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14846_ _07996_ _07976_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17565_ _10562_ _10563_ vssd1 vssd1 vccd1 vccd1 _10564_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _07774_ _07524_ _07925_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__or3_1
X_11989_ net3040 net2955 vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19304_ net4124 _03146_ net619 _03155_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ _09586_ _09587_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ _06874_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1__f__05942_ clknet_0__05942_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05942_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _10493_ _10494_ vssd1 vssd1 vccd1 vccd1 _10495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19235_ _03036_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16447_ _09184_ _09275_ _09402_ _09519_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ _06676_ _06759_ _06760_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__or3_1
XFILLER_0_184_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7009 rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 net7533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_71_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19166_ net2553 _03066_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16378_ _09449_ _09450_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6308 net2295 vssd1 vssd1 vccd1 vccd1 net6832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6319 rbzero.tex_g0\[24\] vssd1 vssd1 vccd1 vccd1 net6843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18117_ _02161_ _02163_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__nand2_1
X_15329_ _08307_ _08400_ _08401_ _08403_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5607 _00961_ vssd1 vssd1 vccd1 vccd1 net6131 sky130_fd_sc_hd__dlygate4sd3_1
X_19097_ _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5618 _02965_ vssd1 vssd1 vccd1 vccd1 net6142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5629 _08206_ vssd1 vssd1 vccd1 vccd1 net6153 sky130_fd_sc_hd__dlygate4sd3_1
X_18048_ _02094_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4906 net1007 vssd1 vssd1 vccd1 vccd1 net5430 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_86_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold4917 rbzero.mapdyw\[0\] vssd1 vssd1 vccd1 vccd1 net5441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4928 net1086 vssd1 vssd1 vccd1 vccd1 net5452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4939 net2933 vssd1 vssd1 vccd1 vccd1 net5463 sky130_fd_sc_hd__buf_1
XFILLER_0_2_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20010_ _03261_ net3744 vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or2_1
X_19999_ net3440 _03578_ net4407 _03550_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21961_ net186 net2205 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21892_ clknet_leaf_96_i_clk net1340 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_20917__330 clknet_1_1__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__inv_2
XFILLER_0_90_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_147_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22444_ clknet_leaf_72_i_clk net2984 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22375_ net507 net2330 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__04011_ clknet_0__04011_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04011_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6831 _02970_ vssd1 vssd1 vccd1 vccd1 net7355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6842 rbzero.spi_registers.buf_sky\[4\] vssd1 vssd1 vccd1 vccd1 net7366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6853 net4827 vssd1 vssd1 vccd1 vccd1 net7377 sky130_fd_sc_hd__clkbuf_1
X_21326_ clknet_leaf_36_i_clk net4273 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20963__372 clknet_1_0__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__inv_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold460 net5292 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
X_21257_ clknet_leaf_71_i_clk net4584 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20662__100 clknet_1_0__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__inv_2
Xhold471 net6358 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ net1980 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__clkbuf_1
Xhold482 net5427 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
X_20208_ net5646 _03717_ _03728_ _03722_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__o211a_1
Xhold493 net5456 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21188_ _02536_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20139_ net3585 _03676_ _03689_ _03683_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _06095_ _06104_ _06108_ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__or4_4
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 net5928 vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _07845_ _07849_ _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a21oi_2
Xhold1171 net5757 vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 net6635 vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _05077_ vssd1 vssd1 vccd1 vccd1 _05082_
+ sky130_fd_sc_hd__mux2_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _08327_ net7444 vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__nor2_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1193 _01339_ vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _06048_ net38 vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nor2_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _07780_ _07769_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__or2b_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _04983_ _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__or2_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _10225_ _10227_ _10224_ _09797_ vssd1 vssd1 vccd1 vccd1 _10350_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _07649_ _07712_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__nand2_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _04940_ _04943_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nor2_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16301_ _09374_ _09226_ _08328_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__a21o_2
XFILLER_0_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13513_ net7843 vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__buf_2
X_10725_ net2221 net6868 _04225_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
X_17281_ _09139_ _10152_ _10163_ vssd1 vssd1 vccd1 vccd1 _10282_ sky130_fd_sc_hd__or3_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _06859_ _07590_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19020_ net3945 net88 net2978 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__nor3b_1
X_16232_ _09305_ _08793_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13444_ _06592_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_181_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10656_ net6848 net7044 _04192_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ _09215_ _09237_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13375_ net7582 _06139_ _06145_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__o31a_1
XFILLER_0_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15114_ _08218_ net3167 net4582 _08215_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__o211a_1
X_12326_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _05493_ vssd1 vssd1 vccd1 vccd1 _05494_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16094_ _09039_ _09123_ _09168_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _08178_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19922_ net2990 _03477_ _03532_ _03542_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__a211o_1
X_12257_ net3003 _05383_ _05425_ net3952 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11208_ net2597 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
X_19853_ net3030 _08385_ _03484_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
X_12188_ net3762 _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18804_ net6109 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11139_ net6794 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
X_16996_ net4689 net4570 vssd1 vssd1 vccd1 vccd1 _10007_ sky130_fd_sc_hd__nand2_1
X_19784_ net647 _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ _08664_ _09020_ _08961_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__or3b_1
X_18735_ net6186 _06189_ _06191_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or3_1
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18666_ _02637_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _02673_
+ sky130_fd_sc_hd__xnor2_2
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _08347_ _08366_ _08410_ _08432_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17617_ _10526_ _10585_ _01667_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nand3_1
X_14829_ _07467_ _07575_ _07498_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18597_ net6237 _05403_ _02607_ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__nor4_1
XFILLER_0_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__04005_ _04005_ vssd1 vssd1 vccd1 vccd1 clknet_0__04005_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17548_ _10545_ _10546_ vssd1 vssd1 vccd1 vccd1 _10547_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17479_ _09328_ _09666_ vssd1 vssd1 vccd1 vccd1 _10478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19218_ net5178 _03107_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20490_ _03858_ net3531 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6105 rbzero.spi_registers.buf_texadd1\[4\] vssd1 vssd1 vccd1 vccd1 net6629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6116 net1888 vssd1 vssd1 vccd1 vccd1 net6640 sky130_fd_sc_hd__dlygate4sd3_1
X_19149_ net5186 _03066_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__or2_1
Xhold6127 rbzero.tex_r0\[53\] vssd1 vssd1 vccd1 vccd1 net6651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6138 net2113 vssd1 vssd1 vccd1 vccd1 net6662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5404 _04227_ vssd1 vssd1 vccd1 vccd1 net5928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6149 rbzero.tex_r0\[21\] vssd1 vssd1 vccd1 vccd1 net6673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5415 net2726 vssd1 vssd1 vccd1 vccd1 net5939 sky130_fd_sc_hd__dlygate4sd3_1
X_22160_ net292 net2245 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold5426 net2825 vssd1 vssd1 vccd1 vccd1 net5950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5437 rbzero.tex_b1\[25\] vssd1 vssd1 vccd1 vccd1 net5961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4703 _00855_ vssd1 vssd1 vccd1 vccd1 net5227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5448 rbzero.map_overlay.i_otherx\[4\] vssd1 vssd1 vccd1 vccd1 net5972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5459 net2494 vssd1 vssd1 vccd1 vccd1 net5983 sky130_fd_sc_hd__dlygate4sd3_1
X_21111_ _04098_ _04099_ _04100_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__or3_1
Xhold4714 net895 vssd1 vssd1 vccd1 vccd1 net5238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4725 net907 vssd1 vssd1 vccd1 vccd1 net5249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4736 _00741_ vssd1 vssd1 vccd1 vccd1 net5260 sky130_fd_sc_hd__dlygate4sd3_1
X_22091_ clknet_leaf_47_i_clk net4062 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold4747 net880 vssd1 vssd1 vccd1 vccd1 net5271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4758 rbzero.spi_registers.buf_mapdxw\[1\] vssd1 vssd1 vccd1 vccd1 net5282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4769 net984 vssd1 vssd1 vccd1 vccd1 net5293 sky130_fd_sc_hd__dlygate4sd3_1
X_21042_ net5424 _03519_ _04014_ _04042_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21944_ net169 net1805 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ clknet_leaf_97_i_clk net1126 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20757_ clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__buf_1
XFILLER_0_148_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11490_ _04658_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__06092_ clknet_0__06092_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__06092_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22427_ clknet_leaf_46_i_clk net4765 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
Xhold7362 _08046_ vssd1 vssd1 vccd1 vccd1 net7886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7384 _06689_ vssd1 vssd1 vccd1 vccd1 net7908 sky130_fd_sc_hd__buf_2
XFILLER_0_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6650 rbzero.tex_r1\[31\] vssd1 vssd1 vccd1 vccd1 net7174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6661 net2816 vssd1 vssd1 vccd1 vccd1 net7185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13160_ net3054 vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__inv_2
X_22358_ net490 net1460 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold6672 rbzero.tex_r1\[18\] vssd1 vssd1 vccd1 vccd1 net7196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6683 net2759 vssd1 vssd1 vccd1 vccd1 net7207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6694 rbzero.tex_b0\[11\] vssd1 vssd1 vccd1 vccd1 net7218 sky130_fd_sc_hd__dlygate4sd3_1
X_12111_ rbzero.tex_r1\[21\] rbzero.tex_r1\[20\] _05263_ vssd1 vssd1 vccd1 vccd1 _05280_
+ sky130_fd_sc_hd__mux2_1
Xhold5960 rbzero.tex_g0\[62\] vssd1 vssd1 vccd1 vccd1 net6484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21309_ clknet_leaf_74_i_clk net4040 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_1
X_13091_ _04837_ _06217_ _06244_ net4675 _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__a221o_1
Xhold5971 net1398 vssd1 vssd1 vccd1 vccd1 net6495 sky130_fd_sc_hd__dlygate4sd3_1
X_22289_ net421 net2749 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
Xhold5982 net1461 vssd1 vssd1 vccd1 vccd1 net6506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5993 _04175_ vssd1 vssd1 vccd1 vccd1 net6517 sky130_fd_sc_hd__dlygate4sd3_1
X_12042_ net4254 _05051_ _05209_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__o21ai_1
Xhold290 net5023 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
X_16850_ _09918_ vssd1 vssd1 vccd1 vccd1 _09919_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _08516_ _08517_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16781_ _09722_ _09723_ vssd1 vssd1 vccd1 vccd1 _09851_ sky130_fd_sc_hd__and2_1
X_13993_ _07139_ _07140_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18520_ _02531_ _02536_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__o21a_1
X_15732_ _08768_ _08774_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18451_ net3742 net4586 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__or2_1
X_15663_ _08735_ _08737_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__nor2_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ net32 _06029_ _06032_ _06023_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a22o_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _10376_ _10401_ vssd1 vssd1 vccd1 vccd1 _10402_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _07751_ _07760_ _07762_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__and3_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _04993_ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__or2_1
X_18382_ net3234 net3396 _02413_ _02414_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__o211ai_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _08667_ _08668_ _08666_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17333_ net3474 net4349 vssd1 vssd1 vccd1 vccd1 _10333_ sky130_fd_sc_hd__nand2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _07687_ _07685_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__xor2_2
X_11757_ _04923_ _04924_ net1504 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a21o_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ _08873_ _09216_ vssd1 vssd1 vccd1 vccd1 _10265_ sky130_fd_sc_hd__nor2_1
X_10708_ net6520 net7266 _04214_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ _07622_ _07626_ _07623_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_125_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11688_ _04161_ _04855_ _04856_ net3929 _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a221o_2
X_19003_ _02973_ _02967_ net3914 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__and3b_1
X_16215_ _09281_ net8010 vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ _06572_ _06573_ _06576_ _06577_ _06541_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a41o_1
XFILLER_0_109_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17195_ _10195_ _10196_ vssd1 vssd1 vccd1 vccd1 _10197_ sky130_fd_sc_hd__nor2_4
X_10639_ net2066 net6371 _04181_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _09219_ _09220_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _06441_ _06442_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _05476_ vssd1 vssd1 vccd1 vccd1 _05477_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16077_ _08514_ _08626_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13289_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] _06417_
+ _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3309 rbzero.pov.ready_buffer\[29\] vssd1 vssd1 vccd1 vccd1 net3833 sky130_fd_sc_hd__buf_1
X_19905_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__clkbuf_4
X_15028_ _08006_ _08031_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__nand2_1
Xhold2608 rbzero.side_hot vssd1 vssd1 vccd1 vccd1 net3480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2619 net7788 vssd1 vssd1 vccd1 vccd1 net3143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19836_ _03471_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__clkbuf_4
Xhold1907 _04567_ vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1918 rbzero.tex_g1\[1\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1929 _04325_ vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19767_ _02998_ _03427_ net1687 _03424_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__o211a_1
X_16979_ _09990_ _09169_ _09991_ vssd1 vssd1 vccd1 vccd1 _09992_ sky130_fd_sc_hd__o21a_1
Xinput3 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
X_18718_ _02707_ _02711_ _02721_ _04624_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19698_ net4328 vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__buf_2
XFILLER_0_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18649_ _02649_ _02657_ _04632_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21660_ clknet_leaf_15_i_clk net5377 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_othery\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ _04760_ _04166_ _04852_ _03952_ net4962 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a41o_1
X_21591_ clknet_leaf_23_i_clk net4213 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20542_ net3600 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ net3422 net1510 _03845_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5201 _00753_ vssd1 vssd1 vccd1 vccd1 net5725 sky130_fd_sc_hd__dlygate4sd3_1
X_22212_ net344 net1952 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5212 net1589 vssd1 vssd1 vccd1 vccd1 net5736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5223 _00526_ vssd1 vssd1 vccd1 vccd1 net5747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5234 net1695 vssd1 vssd1 vccd1 vccd1 net5758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5245 net1522 vssd1 vssd1 vccd1 vccd1 net5769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4500 net814 vssd1 vssd1 vccd1 vccd1 net5024 sky130_fd_sc_hd__dlygate4sd3_1
X_22143_ net275 net1140 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
Xhold5256 net1569 vssd1 vssd1 vccd1 vccd1 net5780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4511 _00874_ vssd1 vssd1 vccd1 vccd1 net5035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4522 _00828_ vssd1 vssd1 vccd1 vccd1 net5046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5267 rbzero.spi_registers.buf_texadd2\[6\] vssd1 vssd1 vccd1 vccd1 net5791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5278 net1915 vssd1 vssd1 vccd1 vccd1 net5802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4533 net792 vssd1 vssd1 vccd1 vccd1 net5057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5289 net1993 vssd1 vssd1 vccd1 vccd1 net5813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4544 net788 vssd1 vssd1 vccd1 vccd1 net5068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3810 net3041 vssd1 vssd1 vccd1 vccd1 net4334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4555 net831 vssd1 vssd1 vccd1 vccd1 net5079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22074_ clknet_leaf_13_i_clk net3517 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3821 rbzero.map_overlay.i_mapdx\[3\] vssd1 vssd1 vccd1 vccd1 net4345 sky130_fd_sc_hd__clkbuf_2
Xhold4566 rbzero.spi_registers.texadd3\[23\] vssd1 vssd1 vccd1 vccd1 net5090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3832 _00970_ vssd1 vssd1 vccd1 vccd1 net4356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4577 rbzero.spi_registers.texadd3\[9\] vssd1 vssd1 vccd1 vccd1 net5101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3843 net7915 vssd1 vssd1 vccd1 vccd1 net4367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4588 net822 vssd1 vssd1 vccd1 vccd1 net5112 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03991_ clknet_0__03991_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03991_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3854 net3120 vssd1 vssd1 vccd1 vccd1 net4378 sky130_fd_sc_hd__clkdlybuf4s25_1
X_21025_ _04023_ _04024_ _04025_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o21a_1
Xhold4599 rbzero.spi_registers.buf_othery\[2\] vssd1 vssd1 vccd1 vccd1 net5123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3865 net670 vssd1 vssd1 vccd1 vccd1 net4389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3876 net6074 vssd1 vssd1 vccd1 vccd1 net4400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3887 net3162 vssd1 vssd1 vccd1 vccd1 net4411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3898 net7743 vssd1 vssd1 vccd1 vccd1 net4422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10990_ net6527 net6768 _04366_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__mux2_1
X_20774__201 clknet_1_1__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__inv_2
XFILLER_0_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21927_ clknet_leaf_6_i_clk net1176 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _04760_ _04603_ _04637_ _04165_ net4 net5 vssd1 vssd1 vccd1 vccd1 _05822_
+ sky130_fd_sc_hd__mux4_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ clknet_leaf_97_i_clk net4637 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11611_ rbzero.spi_registers.texadd3\[5\] _04640_ _04642_ rbzero.spi_registers.texadd2\[5\]
+ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_194_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _04989_ vssd1 vssd1 vccd1 vccd1 _05756_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21789_ clknet_leaf_11_i_clk net4340 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _07474_ _07400_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14261_ _06737_ net533 _07366_ _07311_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o22ai_1
X_20298__35 clknet_1_0__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
X_11473_ rbzero.spi_registers.texadd3\[13\] _04640_ _04644_ rbzero.spi_registers.texadd1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ _09012_ _09030_ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _06186_ net3804 _06183_ net4821 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__and4_1
X_14192_ _07288_ _07308_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6480 net1953 vssd1 vssd1 vccd1 vccd1 net7004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6491 rbzero.tex_g0\[11\] vssd1 vssd1 vccd1 vccd1 net7015 sky130_fd_sc_hd__dlygate4sd3_1
X_13143_ net3433 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5790 _00481_ vssd1 vssd1 vccd1 vccd1 net6314 sky130_fd_sc_hd__dlygate4sd3_1
X_17951_ _08634_ _09251_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__or2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _04823_ net3983 _06181_ net3952 vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16902_ net890 _09939_ _09940_ rbzero.wall_tracer.visualWallDist\[-8\] vssd1 vssd1
+ vccd1 vccd1 _00502_ sky130_fd_sc_hd__a22o_1
X_12025_ net4060 net4034 vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nand2_2
X_17882_ _01911_ _01912_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19621_ net5011 net799 _03347_ _03343_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__o211a_1
X_16833_ _09656_ _09765_ _09902_ vssd1 vssd1 vccd1 vccd1 _09903_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16764_ _08317_ _08498_ _08588_ _08556_ vssd1 vssd1 vccd1 vccd1 _09834_ sky130_fd_sc_hd__or4_2
X_19552_ net3038 _03305_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or2_1
X_13976_ _07121_ _07122_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ _08788_ _08789_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__nor2_4
X_18503_ net2977 net1577 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__and2b_1
X_12927_ net4021 _05299_ _04802_ net4002 net34 net36 vssd1 vssd1 vccd1 vccd1 _06084_
+ sky130_fd_sc_hd__mux4_1
X_16695_ _09656_ _09765_ vssd1 vssd1 vccd1 vccd1 _09766_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_158_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19483_ net3151 _03239_ net3075 vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__or3b_1
X_15646_ _08716_ _08719_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__nor2_1
X_18434_ net4513 net4431 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ net44 _06008_ _05997_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a21bo_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11809_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__clkbuf_8
X_18365_ _02398_ _02399_ net3394 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15577_ _08648_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12789_ _05944_ _05947_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _10189_ _10190_ vssd1 vssd1 vccd1 vccd1 _10317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _07671_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__xor2_4
X_18296_ net4467 net4310 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _10246_ _10247_ vssd1 vssd1 vccd1 vccd1 _10248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03985_ _03985_ vssd1 vssd1 vccd1 vccd1 clknet_0__03985_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_142_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14459_ _07605_ _07608_ _07609_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17178_ _10177_ _10178_ _10166_ vssd1 vssd1 vccd1 vccd1 _10180_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16129_ _08570_ _09186_ _09202_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__nand3_1
Xhold3106 rbzero.wall_tracer.visualWallDist\[3\] vssd1 vssd1 vccd1 vccd1 net3630 sky130_fd_sc_hd__buf_1
Xhold3117 net1237 vssd1 vssd1 vccd1 vccd1 net3641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3128 _03846_ vssd1 vssd1 vccd1 vccd1 net3652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3139 _01187_ vssd1 vssd1 vccd1 vccd1 net3663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2405 _03498_ vssd1 vssd1 vccd1 vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2416 net4892 vssd1 vssd1 vccd1 vccd1 net2940 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2427 rbzero.spi_registers.buf_floor\[3\] vssd1 vssd1 vccd1 vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2438 net4400 vssd1 vssd1 vccd1 vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1704 _04489_ vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2449 rbzero.spi_registers.buf_floor\[1\] vssd1 vssd1 vccd1 vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1715 _01366_ vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1726 _04472_ vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
X_19819_ net3974 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
Xhold1737 _01534_ vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1748 _04441_ vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1759 net6052 vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21712_ clknet_leaf_25_i_clk net1831 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21643_ clknet_leaf_34_i_clk net1542 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21574_ clknet_leaf_4_i_clk net5616 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_41 _10329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_52 net4532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_63 _08195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20525_ _03880_ net3343 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_74 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_96 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20456_ net3653 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5020 net1292 vssd1 vssd1 vccd1 vccd1 net5544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5031 _01047_ vssd1 vssd1 vccd1 vccd1 net5555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5042 net1168 vssd1 vssd1 vccd1 vccd1 net5566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20387_ net3638 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_1
Xhold5053 rbzero.spi_registers.texadd3\[13\] vssd1 vssd1 vccd1 vccd1 net5577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5064 net1265 vssd1 vssd1 vccd1 vccd1 net5588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5075 _01036_ vssd1 vssd1 vccd1 vccd1 net5599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4330 _01096_ vssd1 vssd1 vccd1 vccd1 net4854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4341 net1601 vssd1 vssd1 vccd1 vccd1 net4865 sky130_fd_sc_hd__buf_1
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22126_ net258 net2466 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5086 _00710_ vssd1 vssd1 vccd1 vccd1 net5610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4352 _09959_ vssd1 vssd1 vccd1 vccd1 net4876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5097 net1297 vssd1 vssd1 vccd1 vccd1 net5621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4363 net1130 vssd1 vssd1 vccd1 vccd1 net4887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4374 _06261_ vssd1 vssd1 vccd1 vccd1 net4898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3640 net869 vssd1 vssd1 vccd1 vccd1 net4164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4385 net3402 vssd1 vssd1 vccd1 vccd1 net4909 sky130_fd_sc_hd__buf_2
Xhold4396 _02337_ vssd1 vssd1 vccd1 vccd1 net4920 sky130_fd_sc_hd__clkbuf_2
Xhold3651 net657 vssd1 vssd1 vccd1 vccd1 net4175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3662 net7648 vssd1 vssd1 vccd1 vccd1 net4186 sky130_fd_sc_hd__buf_1
X_22057_ clknet_leaf_90_i_clk net3438 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3673 net7651 vssd1 vssd1 vccd1 vccd1 net4197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3684 net7656 vssd1 vssd1 vccd1 vccd1 net4208 sky130_fd_sc_hd__dlygate4sd3_1
X_21008_ _09920_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__clkbuf_4
Xhold2950 net3166 vssd1 vssd1 vccd1 vccd1 net3474 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3695 net4105 vssd1 vssd1 vccd1 vccd1 net4219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2961 _03913_ vssd1 vssd1 vccd1 vccd1 net3485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2972 net1411 vssd1 vssd1 vccd1 vccd1 net3496 sky130_fd_sc_hd__buf_1
Xhold2983 _04619_ vssd1 vssd1 vccd1 vccd1 net3507 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _06951_ _06980_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__xor2_2
Xhold2994 net7751 vssd1 vssd1 vccd1 vccd1 net3518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _06902_ _06910_ _06879_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__o21a_1
X_10973_ net6856 net7109 _04355_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15500_ _08130_ _08137_ _08144_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__o21a_4
XFILLER_0_179_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap87 _02609_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ _04802_ _05844_ _05852_ net4002 vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16480_ _09544_ _09551_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__xnor2_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _06707_ _06703_ _06765_ _06841_ _06842_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ _08502_ _08505_ _08503_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ _05201_ _05786_ _05796_ net73 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18150_ _02181_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__nand2_1
X_15362_ _08436_ net4063 _06178_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__mux2_1
X_12574_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _05541_ vssd1 vssd1 vccd1 vccd1 _05739_
+ sky130_fd_sc_hd__mux2_1
X_17101_ _10100_ _10101_ vssd1 vssd1 vccd1 vccd1 _10103_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14313_ _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__buf_6
X_18081_ _02004_ _02005_ _02002_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11525_ rbzero.spi_registers.texadd3\[19\] rbzero.spi_registers.texadd1\[19\] rbzero.spi_registers.texadd0\[19\]
+ rbzero.spi_registers.texadd2\[19\] _04692_ _04693_ vssd1 vssd1 vccd1 vccd1 _04697_
+ sky130_fd_sc_hd__mux4_2
X_15293_ _06171_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ _10038_ net4556 net4903 vssd1 vssd1 vccd1 vccd1 _10040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14244_ _07294_ _07346_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__nand3_1
X_11456_ _04628_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ _07267_ _07269_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__and2_1
X_11387_ net7185 net6978 _04573_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ net3447 _06281_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _09948_ _09957_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__xor2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17934_ _01887_ _01888_ _01885_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a21oi_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ net3984 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ _05037_ _05027_ _04974_ _05108_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17865_ _01802_ _09231_ _01913_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__o21ai_1
Xnet99_2 clknet_1_1__leaf__04800_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
X_19604_ net5222 _03325_ _03337_ _03330_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16816_ _09881_ _09882_ _09884_ vssd1 vssd1 vccd1 vccd1 _09886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17796_ _01844_ _01845_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19535_ _03000_ _03289_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16747_ _09811_ _09816_ vssd1 vssd1 vccd1 vccd1 _09817_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _07108_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__xor2_2
XFILLER_0_202_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16678_ _09600_ _09616_ _09748_ vssd1 vssd1 vccd1 vccd1 _09749_ sky130_fd_sc_hd__a21oi_1
X_19466_ _02492_ _03238_ net3076 net6302 vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18417_ net4483 net4368 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15629_ _08699_ _08700_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20911__325 clknet_1_1__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__inv_2
X_19397_ _03035_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18348_ _02384_ _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18279_ _02280_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 i_test_wci vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_8
X_21290_ clknet_leaf_89_i_clk net4047 vssd1 vssd1 vccd1 vccd1 reg_rgb\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold801 net5220 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 net5485 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold823 net6444 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
X_20241_ _08275_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__clkbuf_4
Xhold834 net6462 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 net5634 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 net5682 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold867 net5659 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 net5701 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__buf_1
X_20172_ _03440_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__clkbuf_4
Xhold889 net3529 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2202 net5938 vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_196_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2213 net7212 vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 _04315_ vssd1 vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 net7206 vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 rbzero.tex_g0\[63\] vssd1 vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1501 _04421_ vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 _01173_ vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2257 net7176 vssd1 vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 _01430_ vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2268 net5948 vssd1 vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1534 net6989 vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2279 net5919 vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1545 net4390 vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__clkbuf_2
Xhold1556 net6899 vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 _03370_ vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1578 _04249_ vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 net6661 vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21626_ clknet_leaf_5_i_clk net5005 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20886__302 clknet_1_0__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__inv_2
XFILLER_0_30_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21557_ clknet_leaf_2_i_clk net806 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11310_ net6616 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20508_ net3573 net1270 _03867_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__mux2_1
X_12290_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _05457_ vssd1 vssd1 vccd1 vccd1 _05458_
+ sky130_fd_sc_hd__mux2_1
X_21488_ clknet_leaf_15_i_clk net2918 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11241_ net2796 net6539 _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__mux2_1
X_20439_ net3298 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ net6596 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4160 _00665_ vssd1 vssd1 vccd1 vccd1 net4684 sky130_fd_sc_hd__dlygate4sd3_1
X_22109_ net241 net2883 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
X_15980_ _08587_ _08501_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__or2_1
Xhold4182 _01610_ vssd1 vssd1 vccd1 vccd1 net4706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4193 _08257_ vssd1 vssd1 vccd1 vccd1 net4717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3470 net6314 vssd1 vssd1 vccd1 vccd1 net3994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3481 net4042 vssd1 vssd1 vccd1 vccd1 net4005 sky130_fd_sc_hd__clkbuf_2
X_14931_ net7843 _08003_ vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__and2_1
Xhold3492 _03955_ vssd1 vssd1 vccd1 vccd1 net4016 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21002__4 clknet_1_0__leaf__03773_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2780 _01217_ vssd1 vssd1 vccd1 vccd1 net3304 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _10406_ _10416_ _10539_ _09108_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__o22ai_1
Xhold2791 net7820 vssd1 vssd1 vccd1 vccd1 net3315 sky130_fd_sc_hd__dlygate4sd3_1
X_14862_ net7434 _08012_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__nor2_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20991__17 clknet_1_0__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _09549_ _09550_ _09548_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_188_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13813_ _06961_ _06962_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__nor2_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ _10504_ _10472_ vssd1 vssd1 vccd1 vccd1 _10579_ sky130_fd_sc_hd__or2b_1
X_14793_ _07936_ _07942_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16532_ _09096_ _09603_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19320_ _03141_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__clkbuf_4
X_13744_ _06826_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__clkbuf_4
X_10956_ net6433 net6850 _04344_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16463_ _09445_ _09461_ _09534_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_183_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19251_ net4121 _03119_ net604 _03128_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ _06822_ _06823_ _06716_ _06825_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o2bb2a_4
X_10887_ net6918 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__clkbuf_1
X_15414_ net3217 _08304_ _08307_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18202_ _02080_ _02248_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19182_ net5117 _03078_ _03087_ _03074_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12626_ _05784_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand2_1
X_16394_ _08424_ _08574_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _02103_ _02105_ _02179_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15345_ _08418_ _08419_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__nand2_1
X_12557_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _04989_ vssd1 vssd1 vccd1 vccd1 _05722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18064_ _02110_ _02111_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__nand2_1
X_11508_ _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__nand2b_4
X_15276_ net7511 _08350_ _08304_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__a21o_4
X_12488_ _05028_ _05628_ _05636_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a31o_1
XFILLER_0_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 net4346 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
X_17015_ net4597 net4370 vssd1 vssd1 vccd1 vccd1 _10024_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14227_ _06880_ _07082_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__nand2_1
Xhold119 _03021_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11439_ net4010 _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _07276_ _07286_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13109_ net2879 _06244_ _06196_ net2726 _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a221o_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _07236_ _07238_ _07234_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18966_ net3822 _06217_ _01749_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _01965_ _01966_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__nand2_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18897_ _02880_ net4758 _02879_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17848_ _01891_ _01806_ _01896_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__and3_1
XFILLER_0_191_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17779_ _01828_ _01829_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19518_ _02998_ _03275_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19449_ net1571 net3254 _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22460_ clknet_leaf_38_i_clk _01629_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21411_ clknet_leaf_79_i_clk net3239 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22391_ net523 net1994 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21342_ clknet_leaf_42_i_clk net4181 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold620 net4935 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21273_ clknet_leaf_51_i_clk _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold631 _01492_ vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 net4502 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20729__161 clknet_1_1__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__inv_2
Xhold653 net3465 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20224_ net5193 _03731_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold664 net4862 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold675 net3678 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 net4834 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 net4885 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20155_ net5566 _03692_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__or2_1
Xhold2010 _03405_ vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 _04475_ vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2032 net7240 vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2043 _01324_ vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20086_ net3561 _04241_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nor2_1
Xhold2054 net2565 vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2065 _01303_ vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 net6059 vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _01565_ vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2076 net7130 vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1342 _04358_ vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2087 net5968 vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__buf_1
Xhold2098 net7190 vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 net6609 vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1364 net6639 vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 _01383_ vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1386 _03397_ vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1397 _04155_ vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10810_ _04243_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _04928_ _04932_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o21bai_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10741_ net2754 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ net84 _06589_ _06597_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__nand4_4
X_10672_ _04169_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _05279_ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21609_ clknet_leaf_20_i_clk net5265 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13391_ _06527_ _06539_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _08218_ _08237_ net3773 _08239_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__o211a_1
X_12342_ _05508_ _05509_ _04991_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ _06386_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _04614_ _04790_ _04161_ _04601_ _04608_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a2111oi_1
X_14012_ _07157_ _07162_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__nand2b_1
X_11224_ net5872 net7054 _04492_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ net7575 _02801_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20940__351 clknet_1_1__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__inv_2
X_11155_ net2244 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
X_18751_ net3952 _02747_ _09999_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
X_15963_ _09034_ _09033_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__or2b_1
X_11086_ net6318 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17702_ _01751_ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__or2b_1
X_14914_ _06664_ _08006_ _08061_ net7457 vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__a31o_1
X_15894_ _08404_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__inv_2
X_18682_ _02673_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__inv_2
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _10520_ _09484_ _09861_ _01684_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__o22ai_1
X_14845_ _07695_ _07971_ _07693_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__a21o_1
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17564_ _10342_ _10440_ _10439_ vssd1 vssd1 vccd1 vccd1 _10563_ sky130_fd_sc_hd__a21oi_2
X_14776_ _07925_ _07926_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__xnor2_1
X_11988_ _05154_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19303_ net3011 _03147_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__or2_1
X_16515_ _09103_ _09216_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__nor2_1
X_13727_ _06875_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__xnor2_1
X_10939_ net6369 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__clkbuf_1
X_17495_ _10492_ _10491_ vssd1 vssd1 vccd1 vccd1 _10494_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19234_ net5609 _03106_ _03118_ _03115_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__o211a_1
X_16446_ _09301_ _09273_ _09401_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__a21oi_1
X_13658_ _06608_ _06688_ _06753_ _06692_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12609_ _05208_ _05773_ _05619_ _05095_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a211o_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20334__67 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
X_16377_ _09091_ _08707_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__nor2_1
X_19165_ net4197 _03065_ net1142 _03074_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13589_ _06530_ _06631_ _06687_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__mux2_1
Xhold6309 _04566_ vssd1 vssd1 vccd1 vccd1 net6833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15328_ _08341_ _08402_ _08307_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__o21a_1
X_18116_ _02161_ _02163_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__or2_1
X_19096_ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18047_ _01802_ _09602_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__nor2_1
X_15259_ _08333_ net3024 _06177_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4907 net5444 vssd1 vssd1 vccd1 vccd1 net5431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4918 net1054 vssd1 vssd1 vccd1 vccd1 net5442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4929 _00724_ vssd1 vssd1 vccd1 vccd1 net5453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19998_ net4406 _03582_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18949_ net3136 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21960_ net185 net1033 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21891_ clknet_leaf_96_i_clk net1293 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20759__187 clknet_1_0__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__inv_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22443_ clknet_leaf_72_i_clk net3536 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22374_ net506 net2009 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__04010_ clknet_0__04010_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04010_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6821 _03589_ vssd1 vssd1 vccd1 vccd1 net7345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6832 rbzero.spi_registers.spi_counter\[3\] vssd1 vssd1 vccd1 vccd1 net7356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6843 net7725 vssd1 vssd1 vccd1 vccd1 net7367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6854 _09790_ vssd1 vssd1 vccd1 vccd1 net7378 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21325_ clknet_leaf_36_i_clk net4241 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold450 net5280 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
X_21256_ clknet_leaf_52_i_clk net4786 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold461 net5470 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 net6360 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold483 net5429 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
X_20207_ net5626 _03718_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__or2_1
Xhold494 rbzero.pov.ready_buffer\[52\] vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
X_21187_ _02531_ _02537_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20138_ net5410 _03679_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__or2_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _05396_ net3615 _03580_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__mux2_1
X_12960_ _06112_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__or2_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 net6663 vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 _01535_ vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _05077_ vssd1 vssd1 vccd1 vccd1 _05081_
+ sky130_fd_sc_hd__mux2_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 net5759 vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 net6637 vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ net37 vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__inv_2
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 net6649 vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _07769_ _07780_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__xnor2_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _04988_ vssd1 vssd1 vccd1 vccd1 _05012_
+ sky130_fd_sc_hd__mux2_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _07647_ _07648_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__nand2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ net1886 _04941_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a21boi_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16300_ net3103 _08628_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__nand2_1
X_13512_ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__clkbuf_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ net6447 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__clkbuf_1
X_17280_ _10155_ _10156_ _10280_ vssd1 vssd1 vccd1 vccd1 _10281_ sky130_fd_sc_hd__a21bo_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _07615_ _07631_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__xnor2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16231_ _09304_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__clkbuf_4
X_13443_ _06516_ _06495_ _06560_ _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__a2bb2o_2
X_10655_ net6690 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16162_ _09234_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__xnor2_2
X_13374_ net7552 net7582 _04635_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ net4581 _08223_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__or2_1
X_12325_ _04986_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__buf_4
X_16093_ _09118_ _09113_ _09166_ _09167_ _09076_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_121_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15044_ net4386 _08177_ _08138_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__mux2_1
X_19921_ _08398_ _03480_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__nor2_1
X_12256_ _05365_ _05353_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__and2_1
XFILLER_0_181_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11207_ net7107 net7097 _04481_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19852_ net5463 _03475_ _03489_ _03454_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__o211a_1
X_12187_ _05344_ net3910 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__or2b_1
XFILLER_0_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18803_ rbzero.wall_tracer.rayAddendY\[-2\] _02795_ _02714_ vssd1 vssd1 vccd1 vccd1
+ _02796_ sky130_fd_sc_hd__mux2_1
X_11138_ net6792 net2616 _04448_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__mux2_1
X_19783_ _03428_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16995_ net4689 net4570 vssd1 vssd1 vccd1 vccd1 _10006_ sky130_fd_sc_hd__nor2_1
X_18734_ net3883 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__clkbuf_1
X_11069_ net2425 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
X_15946_ _08962_ _08755_ _09020_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18665_ _02579_ net4768 net7609 net3552 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a31o_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _08387_ _08456_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__nor2_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _10526_ _10585_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14828_ _07494_ _07566_ vssd1 vssd1 vccd1 vccd1 _07979_ sky130_fd_sc_hd__nand2_2
X_18596_ net4463 net4446 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__04004_ _04004_ vssd1 vssd1 vccd1 vccd1 clknet_0__04004_ sky130_fd_sc_hd__clkbuf_16
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ _10301_ _10422_ vssd1 vssd1 vccd1 vccd1 _10546_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14759_ _07907_ _07909_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17478_ _10475_ _10476_ vssd1 vssd1 vccd1 vccd1 _10477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19217_ net5780 _03106_ _03109_ _03096_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__o211a_1
X_16429_ _09475_ _09501_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6106 net1829 vssd1 vssd1 vccd1 vccd1 net6630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6117 rbzero.tex_r1\[23\] vssd1 vssd1 vccd1 vccd1 net6641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19148_ net5947 _03065_ _03067_ _03061_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__o211a_1
Xhold6128 net1723 vssd1 vssd1 vccd1 vccd1 net6652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20947__357 clknet_1_1__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__inv_2
Xhold6139 rbzero.tex_g0\[23\] vssd1 vssd1 vccd1 vccd1 net6663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5405 net1684 vssd1 vssd1 vccd1 vccd1 net5929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5416 _00676_ vssd1 vssd1 vccd1 vccd1 net5940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19079_ net2962 net2979 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__or2_1
Xhold5427 _00668_ vssd1 vssd1 vccd1 vccd1 net5951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5438 net2182 vssd1 vssd1 vccd1 vccd1 net5962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4704 net887 vssd1 vssd1 vccd1 vccd1 net5228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5449 net2839 vssd1 vssd1 vccd1 vccd1 net5973 sky130_fd_sc_hd__dlygate4sd3_1
X_21110_ net4143 net4649 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__and2_1
Xhold4715 rbzero.pov.spi_buffer\[45\] vssd1 vssd1 vccd1 vccd1 net5239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4726 rbzero.pov.spi_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net5250 sky130_fd_sc_hd__dlygate4sd3_1
X_22090_ clknet_leaf_48_i_clk _01259_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4737 net901 vssd1 vssd1 vccd1 vccd1 net5261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4748 _01591_ vssd1 vssd1 vccd1 vccd1 net5272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4759 net865 vssd1 vssd1 vccd1 vccd1 net5283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21041_ _04038_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21943_ net168 net2372 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21874_ clknet_leaf_97_i_clk net1223 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20692__127 clknet_1_0__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__inv_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22426_ clknet_leaf_50_i_clk net5457 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20313__48 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XFILLER_0_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7363 rbzero.row_render.size\[9\] vssd1 vssd1 vccd1 vccd1 net7887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6640 _04275_ vssd1 vssd1 vccd1 vccd1 net7164 sky130_fd_sc_hd__dlygate4sd3_1
X_22357_ net489 net2395 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6651 net2635 vssd1 vssd1 vccd1 vccd1 net7175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6662 rbzero.tex_b1\[11\] vssd1 vssd1 vccd1 vccd1 net7186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6673 net2731 vssd1 vssd1 vccd1 vccd1 net7197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _04993_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__clkbuf_8
Xhold6684 rbzero.tex_r1\[25\] vssd1 vssd1 vccd1 vccd1 net7208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5950 _04526_ vssd1 vssd1 vccd1 vccd1 net6474 sky130_fd_sc_hd__dlygate4sd3_1
X_21308_ clknet_leaf_48_i_clk net4012 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold6695 net2692 vssd1 vssd1 vccd1 vccd1 net7219 sky130_fd_sc_hd__dlygate4sd3_1
X_13090_ net3917 net4897 net4913 net3893 vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a22o_1
X_22288_ net420 net2722 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold5961 net1445 vssd1 vssd1 vccd1 vccd1 net6485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5972 rbzero.wall_hot\[0\] vssd1 vssd1 vccd1 vccd1 net6496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5983 rbzero.tex_b0\[26\] vssd1 vssd1 vccd1 vccd1 net6507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5994 net1465 vssd1 vssd1 vccd1 vccd1 net6518 sky130_fd_sc_hd__dlygate4sd3_1
X_12041_ _05105_ _05113_ _05208_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a211o_1
X_21239_ clknet_leaf_62_i_clk _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold280 net5000 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 net5200 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15800_ _08872_ _08873_ _08517_ _08874_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_70_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16780_ _09830_ _09849_ vssd1 vssd1 vccd1 vccd1 _09850_ sky130_fd_sc_hd__xnor2_1
X_13992_ _07119_ _07142_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__and2b_1
XFILLER_0_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _08777_ _08785_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__xnor2_2
X_12943_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xor2_2
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ net3742 net4586 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__nand2_1
X_15662_ _08456_ _08498_ _08736_ _08712_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__o31a_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _06030_ _06031_ net31 vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _10399_ _10400_ vssd1 vssd1 vccd1 vccd1 _10401_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_85_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _04994_ vssd1 vssd1 vccd1 vccd1 _04995_
+ sky130_fd_sc_hd__mux2_1
X_14613_ _07717_ _07734_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__xnor2_2
X_15593_ _08550_ _08625_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__nor2_1
X_18381_ _02413_ _02414_ net3234 net3396 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a211o_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17332_ _10332_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _07693_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__nor2_2
X_11756_ _04922_ _04923_ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nand3_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ net7199 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17263_ _10262_ _10263_ vssd1 vssd1 vccd1 vccd1 _10264_ sky130_fd_sc_hd__and2_1
X_14475_ _07623_ _07625_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__nor2_2
XFILLER_0_154_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11687_ net3936 net3992 net1 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or3b_1
XFILLER_0_153_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ net3913 _02970_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16214_ _09284_ net3025 _09288_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__a21oi_1
X_13426_ net7442 _06431_ _06545_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__o21ai_1
X_17194_ _10192_ _10194_ vssd1 vssd1 vccd1 vccd1 _10196_ sky130_fd_sc_hd__and2_1
X_10638_ net2138 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _08587_ _08574_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__nor2_1
X_13357_ _04635_ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__nand2_2
XFILLER_0_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _05456_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__buf_4
X_16076_ _08309_ _08632_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_23_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13288_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__and2_1
X_19904_ net41 _03473_ _03035_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__o21a_2
X_15027_ _08128_ _08141_ _08069_ vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__mux2_1
X_12239_ rbzero.debug_overlay.vplaneX\[-3\] _05373_ _05405_ _05407_ vssd1 vssd1 vccd1
+ vccd1 _05408_ sky130_fd_sc_hd__a211o_1
Xhold2609 _02806_ vssd1 vssd1 vccd1 vccd1 net3133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19835_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__clkbuf_4
Xhold1908 _01137_ vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1919 net5832 vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_38_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19766_ net6590 _03429_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__or2_1
X_16978_ _09990_ _09169_ net3508 vssd1 vssd1 vccd1 vccd1 _09991_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
X_18717_ net4587 _05401_ _02711_ _02647_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a211oi_1
X_15929_ _09002_ _09003_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19697_ net4327 net3075 net3151 vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__or3b_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18648_ _02655_ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or2_1
X_18579_ net3838 _02569_ _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20610_ _04777_ net2987 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21590_ clknet_leaf_23_i_clk net5676 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20541_ _03902_ net3599 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20472_ _08275_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22211_ net343 net1997 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
Xhold5202 net1558 vssd1 vssd1 vccd1 vccd1 net5726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5213 _00761_ vssd1 vssd1 vccd1 vccd1 net5737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5224 net2788 vssd1 vssd1 vccd1 vccd1 net5748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5235 _00762_ vssd1 vssd1 vccd1 vccd1 net5759 sky130_fd_sc_hd__dlygate4sd3_1
X_22142_ net274 net1374 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
Xhold5246 rbzero.pov.spi_buffer\[59\] vssd1 vssd1 vccd1 vccd1 net5770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4501 rbzero.spi_registers.texadd1\[6\] vssd1 vssd1 vccd1 vccd1 net5025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5257 _00702_ vssd1 vssd1 vccd1 vccd1 net5781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4512 net782 vssd1 vssd1 vccd1 vccd1 net5036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4523 net787 vssd1 vssd1 vccd1 vccd1 net5047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5268 net1217 vssd1 vssd1 vccd1 vccd1 net5792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5279 _00705_ vssd1 vssd1 vccd1 vccd1 net5803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4534 _00857_ vssd1 vssd1 vccd1 vccd1 net5058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4545 _00691_ vssd1 vssd1 vccd1 vccd1 net5069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3800 net1864 vssd1 vssd1 vccd1 vccd1 net4324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3811 net7369 vssd1 vssd1 vccd1 vccd1 net4335 sky130_fd_sc_hd__buf_4
X_22073_ clknet_leaf_9_i_clk net3682 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4556 _00848_ vssd1 vssd1 vccd1 vccd1 net5080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3822 _00669_ vssd1 vssd1 vccd1 vccd1 net4346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4567 net790 vssd1 vssd1 vccd1 vccd1 net5091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3833 net2913 vssd1 vssd1 vccd1 vccd1 net4357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4578 net921 vssd1 vssd1 vccd1 vccd1 net5102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03990_ clknet_0__03990_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03990_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3844 net3103 vssd1 vssd1 vccd1 vccd1 net4368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4589 rbzero.pov.spi_buffer\[31\] vssd1 vssd1 vccd1 vccd1 net5113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21024_ net5271 _03519_ _04014_ _04027_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3855 net7892 vssd1 vssd1 vccd1 vccd1 net4379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3866 rbzero.row_render.size\[8\] vssd1 vssd1 vccd1 vccd1 net4390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3877 net2962 vssd1 vssd1 vccd1 vccd1 net4401 sky130_fd_sc_hd__clkbuf_2
Xhold3899 net3169 vssd1 vssd1 vccd1 vccd1 net4423 sky130_fd_sc_hd__buf_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21926_ clknet_leaf_6_i_clk net1248 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ clknet_leaf_82_i_clk net4750 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ rbzero.spi_registers.texadd1\[5\] _04644_ _04709_ rbzero.spi_registers.texadd0\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _05177_ _05752_ _05754_ _05000_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21788_ clknet_leaf_11_i_clk net5465 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11541_ net4891 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _07311_ _06737_ net532 _07366_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__or4_1
XFILLER_0_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11472_ _04639_ _04638_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_190_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ _06360_ _06361_ _06363_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__o31a_1
X_22409_ net161 net2822 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14191_ _07339_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__xnor2_1
Xhold7193 rbzero.traced_texVinit\[9\] vssd1 vssd1 vccd1 vccd1 net7717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6470 net2550 vssd1 vssd1 vccd1 vccd1 net6994 sky130_fd_sc_hd__dlygate4sd3_1
X_13142_ net3179 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__inv_2
Xhold6481 rbzero.tex_r1\[46\] vssd1 vssd1 vccd1 vccd1 net7005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6492 net1750 vssd1 vssd1 vccd1 vccd1 net7016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17950_ _01997_ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__xnor2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5780 net3197 vssd1 vssd1 vccd1 vccd1 net6304 sky130_fd_sc_hd__clkbuf_2
X_13073_ net4874 vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5791 rbzero.tex_g0\[32\] vssd1 vssd1 vccd1 vccd1 net6315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12024_ net4033 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__buf_4
X_16901_ _09935_ vssd1 vssd1 vccd1 vccd1 _09940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17881_ _01920_ _01930_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19620_ net3100 _03340_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__or2_1
X_16832_ _09762_ _09764_ vssd1 vssd1 vccd1 vccd1 _09902_ sky130_fd_sc_hd__nor2_1
X_19551_ net5190 _03303_ _03307_ _03295_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__o211a_1
X_16763_ _08701_ _08849_ vssd1 vssd1 vccd1 vccd1 _09833_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13975_ _07123_ _07124_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18502_ net3945 _04241_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__nor2_1
X_15714_ _08746_ _08787_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__and2_4
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12926_ _06052_ net36 _06079_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a31o_1
X_19482_ net3118 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__clkbuf_1
X_16694_ _09762_ _09764_ vssd1 vssd1 vccd1 vccd1 _09765_ sky130_fd_sc_hd__xor2_4
XFILLER_0_185_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18433_ net4513 net4431 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__nor2_1
X_15645_ _08716_ _08719_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__nand2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ net30 _06011_ _06014_ _06002_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_115_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11808_ net81 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__buf_6
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18364_ _02390_ _02391_ net3393 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__o21ai_1
X_15576_ _08636_ _08640_ _08647_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _05945_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _10253_ _10315_ vssd1 vssd1 vccd1 vccd1 _10316_ sky130_fd_sc_hd__xnor2_2
X_11739_ net42 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14527_ _07672_ _07674_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__o21a_2
X_18295_ _02339_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03984_ _03984_ vssd1 vssd1 vccd1 vccd1 clknet_0__03984_ sky130_fd_sc_hd__clkbuf_16
X_17246_ _10244_ _10245_ vssd1 vssd1 vccd1 vccd1 _10247_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _07471_ _07354_ _07606_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13409_ _06472_ _06477_ _06433_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a21o_2
X_17177_ _10166_ _10177_ _10178_ vssd1 vssd1 vccd1 vccd1 _10179_ sky130_fd_sc_hd__nand3_1
XFILLER_0_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14389_ _07537_ _07539_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16128_ _08570_ _09186_ _09202_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3107 _08230_ vssd1 vssd1 vccd1 vccd1 net3631 sky130_fd_sc_hd__dlygate4sd3_1
X_16059_ _08724_ _08664_ _09133_ _08665_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__a2bb2o_1
Xhold3118 _03785_ vssd1 vssd1 vccd1 vccd1 net3642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3129 _03847_ vssd1 vssd1 vccd1 vccd1 net3653 sky130_fd_sc_hd__dlygate4sd3_1
X_20997__23 clknet_1_1__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
Xhold2406 net6131 vssd1 vssd1 vccd1 vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2417 net4894 vssd1 vssd1 vccd1 vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2428 net7328 vssd1 vssd1 vccd1 vccd1 net2952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2439 _00649_ vssd1 vssd1 vccd1 vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1705 _01301_ vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
X_20723__156 clknet_1_0__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__inv_2
Xhold1716 net6855 vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
X_19818_ _02967_ net3973 vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and2_1
XFILLER_0_209_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1727 _01317_ vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1738 net7025 vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1749 _01345_ vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
X_19749_ net4401 _03392_ net1575 _03413_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21711_ clknet_leaf_26_i_clk net1669 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21642_ clknet_leaf_29_i_clk net3126 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_20 _05892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21573_ clknet_leaf_4_i_clk net5184 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_31 _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 _10329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ net2956 net3342 _03889_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__mux2_1
XANTENNA_53 net4779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 _08479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_75 net3222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_86 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20455_ _03836_ net3652 vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5010 _01070_ vssd1 vssd1 vccd1 vccd1 net5534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5021 _01060_ vssd1 vssd1 vccd1 vccd1 net5545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5032 rbzero.pov.spi_buffer\[3\] vssd1 vssd1 vccd1 vccd1 net5556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5043 _01050_ vssd1 vssd1 vccd1 vccd1 net5567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20386_ _03791_ net3637 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5054 net1261 vssd1 vssd1 vccd1 vccd1 net5578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4320 net3561 vssd1 vssd1 vccd1 vccd1 net4844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5065 _01094_ vssd1 vssd1 vccd1 vccd1 net5589 sky130_fd_sc_hd__dlygate4sd3_1
X_22125_ net257 net2121 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold5076 rbzero.pov.spi_buffer\[12\] vssd1 vssd1 vccd1 vccd1 net5600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4331 rbzero.pov.spi_buffer\[69\] vssd1 vssd1 vccd1 vccd1 net4855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5087 rbzero.pov.spi_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net5611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4342 _01031_ vssd1 vssd1 vccd1 vccd1 net4866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5098 rbzero.pov.spi_buffer\[53\] vssd1 vssd1 vccd1 vccd1 net5622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4353 _09961_ vssd1 vssd1 vccd1 vccd1 net4877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4364 _00388_ vssd1 vssd1 vccd1 vccd1 net4888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3630 net646 vssd1 vssd1 vccd1 vccd1 net4154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4375 _06267_ vssd1 vssd1 vccd1 vccd1 net4899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3641 net7499 vssd1 vssd1 vccd1 vccd1 net4165 sky130_fd_sc_hd__dlygate4sd3_1
X_22056_ clknet_leaf_90_i_clk net3345 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4386 _04629_ vssd1 vssd1 vccd1 vccd1 net4910 sky130_fd_sc_hd__buf_1
Xhold3652 net7642 vssd1 vssd1 vccd1 vccd1 net4176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4397 rbzero.wall_tracer.mapX\[8\] vssd1 vssd1 vccd1 vccd1 net4921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3663 _00514_ vssd1 vssd1 vccd1 vccd1 net4187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3674 _00683_ vssd1 vssd1 vccd1 vccd1 net4198 sky130_fd_sc_hd__dlygate4sd3_1
X_21007_ _03502_ net1081 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__nor2_1
Xhold2940 net6205 vssd1 vssd1 vccd1 vccd1 net3464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3685 _00769_ vssd1 vssd1 vccd1 vccd1 net4209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2951 net4853 vssd1 vssd1 vccd1 vccd1 net3475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3696 _00963_ vssd1 vssd1 vccd1 vccd1 net4220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2962 _01233_ vssd1 vssd1 vccd1 vccd1 net3486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2973 _03935_ vssd1 vssd1 vccd1 vccd1 net3497 sky130_fd_sc_hd__dlygate4sd3_1
X_20698__133 clknet_1_1__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__inv_2
Xhold2984 _06390_ vssd1 vssd1 vccd1 vccd1 net3508 sky130_fd_sc_hd__buf_4
Xhold2995 rbzero.pov.ready_buffer\[37\] vssd1 vssd1 vccd1 vccd1 net3519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13760_ _06879_ _06902_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__or3_1
X_10972_ net6896 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21909_ clknet_leaf_92_i_clk net5385 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _05825_ _05853_ _05854_ net3965 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a22o_1
Xmax_cap77 _09366_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_6
X_13691_ _06707_ _06708_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15430_ _08503_ _08504_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ _05790_ net6 _05798_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a31o_2
XFILLER_0_183_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _08434_ _08435_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__and2_1
X_12573_ _05736_ _05737_ _05279_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ _10100_ _10101_ vssd1 vssd1 vccd1 vccd1 _10102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14312_ _07405_ _07437_ _07462_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__a21o_1
X_11524_ _04691_ _04694_ _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__and3_1
X_15292_ _08366_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__buf_2
X_18080_ _02126_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17031_ net4902 vssd1 vssd1 vccd1 vccd1 _10039_ sky130_fd_sc_hd__clkbuf_1
X_14243_ _07343_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__xor2_1
X_11455_ net4910 _04626_ _04627_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__or3b_1
XFILLER_0_151_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14174_ _07016_ _07283_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11386_ net6954 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13125_ net3240 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__inv_2
X_18982_ net3923 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _01908_ _01877_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__or2b_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ net3983 vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12007_ _04993_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _01802_ _09231_ _01913_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19603_ net3093 _03327_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__or2_1
X_16815_ _09881_ _09882_ _09884_ vssd1 vssd1 vccd1 vccd1 _09885_ sky130_fd_sc_hd__nand3_1
X_17795_ _01844_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19534_ net5178 _03288_ _03293_ _03295_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__o211a_1
X_16746_ _09676_ _09815_ vssd1 vssd1 vccd1 vccd1 _09816_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13958_ _07062_ _07064_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19465_ _03239_ net3076 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__nand2b_1
X_12909_ net35 net34 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__and2b_1
X_16677_ _09613_ _09615_ vssd1 vssd1 vccd1 vccd1 _09748_ sky130_fd_sc_hd__and2b_1
X_13889_ _06868_ _06872_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__xor2_2
X_18416_ net4483 net4368 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15628_ _08318_ _08702_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19396_ net5398 _03198_ _03210_ _03207_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18347_ net4485 net4353 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15559_ _08633_ _08593_ _08595_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18278_ _02241_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17229_ _10228_ _10229_ vssd1 vssd1 vccd1 vccd1 _10230_ sky130_fd_sc_hd__nor2_1
Xinput40 i_mode[0] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_8
XFILLER_0_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_8
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold802 net5655 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
X_20240_ net3435 _03744_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or2_1
Xhold813 net5622 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 net6446 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold835 _01115_ vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 net3664 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 net3781 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20171_ net3291 _03705_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__or2_1
Xhold868 net5661 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 net5703 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2203 net5940 vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 _04346_ vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2225 _01458_ vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2236 _04271_ vssd1 vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2247 net1982 vssd1 vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1502 _01363_ vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 rbzero.tex_b1\[1\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 _04319_ vssd1 vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2269 net7263 vssd1 vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 net6769 vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _01455_ vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1546 net7661 vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _01529_ vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1568 _00884_ vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 _01518_ vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21625_ clknet_leaf_4_i_clk net5020 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21556_ clknet_leaf_101_i_clk net1380 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20507_ net3367 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21487_ clknet_leaf_15_i_clk net2706 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11240_ _04332_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20438_ _03814_ net3297 vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ net2149 net6594 _04459_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__mux2_1
X_20369_ net719 net3590 _03782_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
Xhold4150 rbzero.debug_overlay.playerY\[1\] vssd1 vssd1 vccd1 vccd1 net4674 sky130_fd_sc_hd__dlygate4sd3_1
X_22108_ net240 net2786 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold4161 net3027 vssd1 vssd1 vccd1 vccd1 net4685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4172 _02660_ vssd1 vssd1 vccd1 vccd1 net4696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4183 net2969 vssd1 vssd1 vccd1 vccd1 net4707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20706__140 clknet_1_0__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__inv_2
XFILLER_0_101_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4194 net7840 vssd1 vssd1 vccd1 vccd1 net4718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3460 _06212_ vssd1 vssd1 vccd1 vccd1 net3984 sky130_fd_sc_hd__clkbuf_4
X_22039_ clknet_leaf_95_i_clk net3698 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3471 rbzero.debug_overlay.playerX\[1\] vssd1 vssd1 vccd1 vccd1 net3995 sky130_fd_sc_hd__buf_2
X_14930_ net7891 _08001_ _08076_ net7566 vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__a211o_1
Xhold3482 _05444_ vssd1 vssd1 vccd1 vccd1 net4006 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3493 _03956_ vssd1 vssd1 vccd1 vccd1 net4017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2770 _01196_ vssd1 vssd1 vccd1 vccd1 net3294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2781 rbzero.pov.ready_buffer\[41\] vssd1 vssd1 vccd1 vccd1 net3305 sky130_fd_sc_hd__dlygate4sd3_1
X_14861_ _07967_ _07794_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__xnor2_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2792 rbzero.pov.ready_buffer\[9\] vssd1 vssd1 vccd1 vccd1 net3316 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ _09669_ _09670_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__and2_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _06961_ _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__and2_1
X_17580_ net7375 _10577_ vssd1 vssd1 vccd1 vccd1 _10578_ sky130_fd_sc_hd__xnor2_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _07534_ _07805_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16531_ net3793 _09304_ _09602_ vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__a21boi_4
X_10955_ net6584 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__clkbuf_1
X_13743_ _06876_ net572 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19250_ _02992_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__clkbuf_4
X_16462_ _09462_ _09443_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__or2b_1
XFILLER_0_196_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ net2057 net6916 _04236_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
X_13674_ _06824_ _06728_ _06724_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18201_ _02246_ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ _08059_ net7764 _08295_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19181_ net1595 _03079_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _05785_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__and2_1
X_16393_ _09358_ _09361_ _09465_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20752__182 clknet_1_0__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__inv_2
X_18132_ _02098_ _02106_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__or2b_1
X_12556_ _05177_ _05718_ _05720_ _05461_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15344_ net2935 _08383_ net4300 vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11507_ _04642_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__inv_2
X_18063_ _02088_ _02109_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__or2_1
X_12487_ _04978_ _05640_ _05644_ _05652_ _05051_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__o311a_1
XFILLER_0_81_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15275_ _08119_ _08124_ _08294_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__a21o_1
Xhold109 net6315 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _10023_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__clkbuf_1
X_14226_ _06837_ _06867_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__or2_1
X_11438_ _04604_ net3908 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__nand2_2
XFILLER_0_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _07260_ _07290_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11369_ net2805 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13108_ net2789 net3804 vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__xor2_1
X_14088_ _07234_ _07236_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__or3_1
X_18965_ net3821 _06219_ _09999_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17916_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__nand2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _06183_ _06179_ _06194_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ _02879_ _02880_ net4758 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__or3_1
X_17847_ _01891_ _01806_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17778_ _09582_ _10416_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19517_ net5124 _03274_ _03284_ _03280_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__o211a_1
X_16729_ _09796_ _09798_ vssd1 vssd1 vccd1 vccd1 _09799_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ net5527 _03198_ _03201_ _03194_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21410_ clknet_leaf_79_i_clk net3205 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22390_ net522 net2154 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21341_ clknet_leaf_42_i_clk net4169 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20360__90 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__inv_2
XFILLER_0_5_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21272_ clknet_leaf_57_i_clk _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold610 net4171 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold621 net4525 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold632 rbzero.pov.ready_buffer\[60\] vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_1
Xhold643 net4504 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_20223_ net5193 _03730_ _03737_ _03735_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold654 _01049_ vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold665 net7881 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold676 net4857 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold687 net7204 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 net5409 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ net5566 _03691_ _03698_ _03696_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__o211a_1
Xhold2000 net6893 vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2011 _00909_ vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2022 _01314_ vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2033 net5915 vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2044 net7140 vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
X_20085_ net6020 _03577_ _03651_ _03636_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__o211a_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2055 _04465_ vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1310 _01327_ vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2066 net6293 vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _03451_ vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 net6735 vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2077 _01400_ vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1343 _01420_ vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2088 net5970 vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1354 net6611 vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2099 _04264_ vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1365 _04443_ vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1376 net6867 vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1387 _00902_ vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _01645_ vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ net7278 net7249 _04236_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ net6628 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12410_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _05476_ vssd1 vssd1 vccd1 vccd1 _05577_
+ sky130_fd_sc_hd__mux2_1
X_21608_ clknet_leaf_20_i_clk net4196 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _06540_ _06481_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__nor2_4
XFILLER_0_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _05493_ vssd1 vssd1 vccd1 vccd1 _05509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21539_ clknet_leaf_28_i_clk net1351 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ _08189_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
X_12272_ _04807_ _05431_ _05440_ _05197_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _07158_ _07160_ _07161_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__a21bo_1
X_11223_ net2509 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ net6547 net2449 _04377_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__mux2_1
X_18750_ _06182_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__xnor2_1
X_15962_ _08992_ _08998_ _09035_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__a21o_1
X_11085_ net6316 net2313 _04415_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__mux2_1
X_17701_ net4433 net4593 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__nand2_1
Xhold3290 _03926_ vssd1 vssd1 vccd1 vccd1 net3814 sky130_fd_sc_hd__dlygate4sd3_1
X_14913_ _07991_ _07989_ _08031_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__a21o_1
X_18681_ _02646_ net3043 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__or2_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _08444_ _08514_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__nor2_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _08872_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__buf_2
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ _06707_ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__buf_2
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17563_ _10471_ _10561_ vssd1 vssd1 vccd1 vccd1 _10562_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ _07774_ _07524_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ net2069 net3040 net2955 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__nand3_1
X_19302_ net4983 _03146_ _03157_ _03155_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__o211a_1
X_16514_ _09064_ _08582_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13726_ _06876_ _06858_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__nor2_1
X_10938_ net2737 net6367 _04344_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
X_17494_ _10491_ _10492_ vssd1 vssd1 vccd1 vccd1 _10493_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20319__54 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_0_168_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19233_ net5057 _03107_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__or2_1
X_16445_ _09516_ _09517_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__nand2_2
XFILLER_0_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10869_ net7247 net7066 _04299_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__mux2_1
X_13657_ _06696_ _06807_ _06692_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ net4239 _05102_ _04984_ _05035_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a2bb2o_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ net1141 _03066_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16376_ _09446_ _09448_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__nand2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _06738_ _06632_ _06695_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__mux2_4
XFILLER_0_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18115_ _01874_ _02063_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15327_ net2935 _08383_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__xnor2_1
X_12539_ _05702_ _05703_ _05261_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__mux2_1
X_19095_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5609 _08193_ vssd1 vssd1 vccd1 vccd1 net6133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18046_ _10259_ _09732_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15258_ net3024 net4355 vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__xor2_1
Xhold4908 net1493 vssd1 vssd1 vccd1 vccd1 net5432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4919 _00680_ vssd1 vssd1 vccd1 vccd1 net5443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14209_ _07356_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__nor2_1
X_15189_ _08273_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
X_19997_ net3301 _03578_ net4562 _03550_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__o211a_1
X_18948_ net3135 _02930_ _02714_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18879_ _02862_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21890_ clknet_leaf_96_i_clk net1264 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22442_ clknet_leaf_72_i_clk net4031 vssd1 vssd1 vccd1 vccd1 rbzero.trace_state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6800 rbzero.pov.spi_counter\[3\] vssd1 vssd1 vccd1 vccd1 net7324 sky130_fd_sc_hd__dlygate4sd3_1
X_22373_ net505 net997 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6811 _03611_ vssd1 vssd1 vccd1 vccd1 net7335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6822 rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1 net7346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6833 _02976_ vssd1 vssd1 vccd1 vccd1 net7357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21324_ clknet_leaf_56_i_clk _00493_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6844 net2985 vssd1 vssd1 vccd1 vccd1 net7368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6855 rbzero.debug_overlay.playerY\[-5\] vssd1 vssd1 vccd1 vccd1 net7379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6877 _08337_ vssd1 vssd1 vccd1 vccd1 net7401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold440 net5313 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
X_21255_ clknet_leaf_52_i_clk net3188 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold451 net5345 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 net5472 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _01542_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
X_20206_ net5626 _03717_ _03727_ _03722_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__o211a_1
Xhold484 net5446 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
X_21186_ _02529_ _02535_ net4658 _02528_ net715 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a32o_1
Xhold495 _03552_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__05891_ clknet_0__05891_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05891_
+ sky130_fd_sc_hd__clkbuf_16
X_20137_ net5410 _03676_ _03688_ _03683_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__o211a_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ net3676 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__clkbuf_1
Xhold1140 net6603 vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 _04432_ vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _05078_ _05079_ _04992_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__mux2_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 net6589 vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 net6849 vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ net4045 net4066 net4083 net4078 _06046_ net37 vssd1 vssd1 vccd1 vccd1 _06047_
+ sky130_fd_sc_hd__mux4_1
Xhold1184 _01409_ vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _03447_ vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _05004_ _05005_ _05007_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__o211a_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818__241 clknet_1_1__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__inv_2
XFILLER_0_200_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ net1010 net1650 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__nand2_1
X_14560_ _07704_ _07710_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__or2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20970__378 clknet_1_1__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__inv_2
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ net1900 net6445 _04225_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
X_13511_ _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__buf_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _07635_ _07634_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__xor2_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16230_ _08328_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__clkbuf_4
X_10654_ net2298 net6688 _04192_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ net4947 _06479_ _06480_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__or3_2
X_16161_ _08590_ _08638_ _09235_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__a21bo_1
X_13373_ _06435_ _06474_ _06522_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15112_ net3166 net3314 _08219_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__mux2_1
X_12324_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _05070_ vssd1 vssd1 vccd1 vccd1 _05492_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16092_ _09107_ _09114_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19920_ net6097 _03530_ net2923 _03496_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__o211a_1
X_12255_ net4063 _05373_ _05368_ net3279 _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a221o_1
X_15043_ _08150_ _08129_ _08175_ _08176_ _08047_ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__a221o_2
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20864__283 clknet_1_1__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__inv_2
X_11206_ net1757 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19851_ _03479_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__or2_1
X_12186_ net3761 _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11137_ net2522 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
X_18802_ _02787_ _02788_ _02794_ _04624_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19782_ _03426_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__buf_4
X_16994_ _09988_ _09997_ _09995_ vssd1 vssd1 vccd1 vccd1 _10005_ sky130_fd_sc_hd__o21a_1
X_18733_ net3882 _06186_ _06394_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
X_11068_ net7113 net6962 _04404_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__mux2_1
X_15945_ _08409_ _08632_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18664_ _02670_ _02671_ rbzero.wall_tracer.rayAddendX\[5\] _09932_ vssd1 vssd1 vccd1
+ vccd1 _02672_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_204_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _08914_ _08923_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__xnor2_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _10596_ _01666_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14827_ _07695_ _07971_ _07976_ _07977_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__a31oi_4
X_18595_ net4463 net4446 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__nor2_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04003_ _04003_ vssd1 vssd1 vccd1 vccd1 clknet_0__04003_ sky130_fd_sc_hd__clkbuf_16
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17546_ _10302_ _10544_ vssd1 vssd1 vccd1 vccd1 _10545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14758_ _07902_ _07908_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__and2_1
XFILLER_0_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13709_ _06660_ _06751_ net582 vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__a21o_4
X_17477_ _09447_ _09794_ _10474_ vssd1 vssd1 vccd1 vccd1 _10476_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14689_ _07795_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19216_ net5547 _03107_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ _09498_ _09500_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6107 rbzero.tex_r0\[23\] vssd1 vssd1 vccd1 vccd1 net6631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19147_ net5014 _03066_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__or2_1
X_16359_ _09424_ _09431_ vssd1 vssd1 vccd1 vccd1 _09432_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6118 net1747 vssd1 vssd1 vccd1 vccd1 net6642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6129 _04257_ vssd1 vssd1 vccd1 vccd1 net6653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5406 rbzero.tex_g1\[47\] vssd1 vssd1 vccd1 vccd1 net5930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5417 rbzero.tex_r0\[62\] vssd1 vssd1 vccd1 vccd1 net5941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19078_ net4401 net2842 _03023_ _03022_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__o211a_1
Xhold5428 rbzero.tex_b0\[59\] vssd1 vssd1 vccd1 vccd1 net5952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5439 _04500_ vssd1 vssd1 vccd1 vccd1 net5963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4705 rbzero.spi_registers.texadd0\[7\] vssd1 vssd1 vccd1 vccd1 net5229 sky130_fd_sc_hd__dlygate4sd3_1
X_18029_ _02075_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4716 net1270 vssd1 vssd1 vccd1 vccd1 net5240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4727 net1232 vssd1 vssd1 vccd1 vccd1 net5251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4738 rbzero.spi_registers.texadd3\[0\] vssd1 vssd1 vccd1 vccd1 net5262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4749 net881 vssd1 vssd1 vccd1 vccd1 net5273 sky130_fd_sc_hd__dlygate4sd3_1
X_21040_ _04039_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__and2b_1
XFILLER_0_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21942_ net167 net2652 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21873_ clknet_leaf_95_i_clk net5253 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ clknet_1_1__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__buf_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7320 rbzero.wall_tracer.stepDistX\[-8\] vssd1 vssd1 vccd1 vccd1 net7844 sky130_fd_sc_hd__dlygate4sd3_1
X_22425_ clknet_leaf_50_i_clk net5426 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7364 net4508 vssd1 vssd1 vccd1 vccd1 net7888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6630 _04183_ vssd1 vssd1 vccd1 vccd1 net7154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7375 rbzero.wall_tracer.stepDistY\[9\] vssd1 vssd1 vccd1 vccd1 net7899 sky130_fd_sc_hd__dlygate4sd3_1
X_22356_ net488 net2725 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold6641 net2645 vssd1 vssd1 vccd1 vccd1 net7165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6652 rbzero.tex_g1\[60\] vssd1 vssd1 vccd1 vccd1 net7176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6663 net2784 vssd1 vssd1 vccd1 vccd1 net7187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6674 _04221_ vssd1 vssd1 vccd1 vccd1 net7198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21307_ clknet_leaf_74_i_clk net3763 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold5940 rbzero.tex_r0\[44\] vssd1 vssd1 vccd1 vccd1 net6464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6685 net2484 vssd1 vssd1 vccd1 vccd1 net7209 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_4_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_206_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5951 net1481 vssd1 vssd1 vccd1 vccd1 net6475 sky130_fd_sc_hd__dlygate4sd3_1
X_22287_ net419 net2112 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
Xhold6696 rbzero.tex_r0\[18\] vssd1 vssd1 vccd1 vccd1 net7220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5962 _04388_ vssd1 vssd1 vccd1 vccd1 net6486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5973 _04639_ vssd1 vssd1 vccd1 vccd1 net6497 sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ net3378 _05095_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5984 net1442 vssd1 vssd1 vccd1 vccd1 net6508 sky130_fd_sc_hd__dlygate4sd3_1
X_21238_ clknet_leaf_62_i_clk _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold270 net7617 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5995 rbzero.tex_r1\[16\] vssd1 vssd1 vccd1 vccd1 net6519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 net5041 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 net5202 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
X_21169_ _09935_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__clkbuf_4
X_13991_ _07113_ _07117_ _07118_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__or3_4
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ _08790_ _08804_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__xnor2_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _06096_ _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nor2_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _08433_ _08516_ _08711_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__o21a_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ net4049 net4891 _04726_ _04777_ net28 net29 vssd1 vssd1 vccd1 vccd1 _06031_
+ sky130_fd_sc_hd__mux4_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17400_ _10377_ _10290_ _10398_ vssd1 vssd1 vccd1 vccd1 _10400_ sky130_fd_sc_hd__nand3_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07751_ _07760_ _07762_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__a21oi_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _04987_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__buf_4
X_18380_ net4429 net4451 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__nand2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08660_ _08662_ _08666_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__a21oi_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17331_ _10331_ net4540 net4903 vssd1 vssd1 vccd1 vccd1 _10332_ sky130_fd_sc_hd__mux2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07641_ _07692_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__nor2_1
X_11755_ net1504 _04923_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nand3_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ net2702 net7197 _04214_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__mux2_1
X_17262_ _10257_ _08708_ _10261_ vssd1 vssd1 vccd1 vccd1 _10263_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14474_ _06923_ _07468_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11686_ net4001 net4972 _04808_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__or3_1
XFILLER_0_181_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19001_ net3913 net3889 _02966_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__and3_1
X_16213_ _09284_ net3025 _09286_ net7371 vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ _06575_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__inv_2
X_17193_ _10192_ _10194_ vssd1 vssd1 vccd1 vccd1 _10195_ sky130_fd_sc_hd__nor2_2
XFILLER_0_154_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ net6371 net6910 _04181_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _09217_ _09218_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__nand2_1
X_13356_ _06443_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _05261_ _05472_ _05474_ _05244_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__o211a_1
X_16075_ _09130_ _09135_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__xor2_1
X_13287_ rbzero.debug_overlay.facingX\[-6\] net3796 vssd1 vssd1 vccd1 vccd1 _06438_
+ sky130_fd_sc_hd__nor2_1
X_19903_ net3159 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
X_15026_ net5684 vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__inv_2
X_12238_ rbzero.debug_overlay.vplaneX\[-4\] _05383_ _05384_ net3838 _04831_ vssd1
+ vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19834_ net40 _03473_ _03034_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__o21a_2
X_12169_ _05336_ _05337_ _04814_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a21oi_1
Xhold1909 net6813 vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_16977_ _09170_ _09121_ vssd1 vssd1 vccd1 vccd1 _09990_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19765_ _02996_ _03427_ net1710 _03424_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15928_ _08968_ _08972_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18716_ _02718_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__xor2_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19696_ net6033 _03359_ net1549 _03384_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18647_ _02627_ _02653_ _02654_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15859_ _08929_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18578_ net3838 net4424 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17529_ _10526_ _10527_ vssd1 vssd1 vccd1 vccd1 _10528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20540_ net668 net3598 _03889_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20471_ net3697 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22210_ net342 net1660 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5203 rbzero.spi_registers.buf_texadd2\[0\] vssd1 vssd1 vccd1 vccd1 net5727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5214 net1590 vssd1 vssd1 vccd1 vccd1 net5738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5225 rbzero.spi_registers.texadd2\[9\] vssd1 vssd1 vccd1 vccd1 net5749 sky130_fd_sc_hd__dlygate4sd3_1
X_22141_ net273 net2190 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5236 net1696 vssd1 vssd1 vccd1 vccd1 net5760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5247 _01095_ vssd1 vssd1 vccd1 vccd1 net5771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4502 net765 vssd1 vssd1 vccd1 vccd1 net5026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4513 rbzero.spi_registers.buf_texadd0\[23\] vssd1 vssd1 vccd1 vccd1 net5037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5258 rbzero.spi_registers.buf_leak\[5\] vssd1 vssd1 vccd1 vccd1 net5782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4524 rbzero.pov.spi_buffer\[32\] vssd1 vssd1 vccd1 vccd1 net5048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5269 _03403_ vssd1 vssd1 vccd1 vccd1 net5793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4535 net793 vssd1 vssd1 vccd1 vccd1 net5059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4546 net789 vssd1 vssd1 vccd1 vccd1 net5070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3801 rbzero.spi_registers.spi_done vssd1 vssd1 vccd1 vccd1 net4325 sky130_fd_sc_hd__dlygate4sd3_1
X_22072_ clknet_leaf_8_i_clk net3673 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3812 _00955_ vssd1 vssd1 vccd1 vccd1 net4336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4557 net832 vssd1 vssd1 vccd1 vccd1 net5081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3823 net632 vssd1 vssd1 vccd1 vccd1 net4347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4568 _00801_ vssd1 vssd1 vccd1 vccd1 net5092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21023_ _04023_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3834 net7445 vssd1 vssd1 vccd1 vccd1 net4358 sky130_fd_sc_hd__clkbuf_4
Xhold4579 _00787_ vssd1 vssd1 vccd1 vccd1 net5103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3845 net7794 vssd1 vssd1 vccd1 vccd1 net4369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3856 net3127 vssd1 vssd1 vccd1 vccd1 net4380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3867 net2069 vssd1 vssd1 vccd1 vccd1 net4391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3878 net7747 vssd1 vssd1 vccd1 vccd1 net4402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3889 _03609_ vssd1 vssd1 vccd1 vccd1 net4413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20700__135 clknet_1_1__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__inv_2
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21925_ clknet_leaf_6_i_clk net1266 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21856_ clknet_leaf_82_i_clk net3703 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21787_ clknet_leaf_11_i_clk net4308 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _04706_ _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11471_ rbzero.spi_registers.texadd3\[14\] _04640_ _04642_ rbzero.spi_registers.texadd2\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20669_ clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__buf_1
XFILLER_0_163_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7150 rbzero.spi_registers.buf_sky\[5\] vssd1 vssd1 vccd1 vccd1 net7674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ _06216_ net4874 _06364_ _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__or4b_1
X_22408_ net160 net2752 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _07277_ _07285_ _07340_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__o21a_1
Xhold7194 net4200 vssd1 vssd1 vccd1 vccd1 net7718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6460 net2408 vssd1 vssd1 vccd1 vccd1 net6984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6471 _04407_ vssd1 vssd1 vccd1 vccd1 net6995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13141_ _06273_ _06275_ _06278_ _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and4b_1
X_20781__207 clknet_1_0__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__inv_2
X_22339_ net471 net2691 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
Xhold6482 net2379 vssd1 vssd1 vccd1 vccd1 net7006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6493 rbzero.tex_r0\[61\] vssd1 vssd1 vccd1 vccd1 net7017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5770 net2590 vssd1 vssd1 vccd1 vccd1 net6294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ net3917 net4897 _06213_ net4090 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__a2bb2o_1
Xhold5781 _02728_ vssd1 vssd1 vccd1 vccd1 net6305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5792 net633 vssd1 vssd1 vccd1 vccd1 net6316 sky130_fd_sc_hd__dlygate4sd3_1
X_12023_ net4059 vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__buf_1
X_16900_ _09933_ vssd1 vssd1 vccd1 vccd1 _09939_ sky130_fd_sc_hd__clkbuf_4
X_17880_ _01928_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16831_ _09792_ _09900_ vssd1 vssd1 vccd1 vccd1 _09901_ sky130_fd_sc_hd__xnor2_2
X_19550_ net3022 _03305_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or2_1
X_16762_ _09725_ _09718_ vssd1 vssd1 vccd1 vccd1 _09832_ sky130_fd_sc_hd__or2b_1
X_13974_ _06826_ _07090_ _06881_ _06923_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__and4b_1
X_20976__384 clknet_1_0__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__inv_2
X_18501_ _02506_ net3212 _02512_ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__or4_1
X_15713_ _08746_ _08787_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__nor2_2
X_12925_ _06080_ _06081_ net36 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__mux2_1
X_19481_ _03261_ net3117 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__or2_1
X_16693_ _09559_ _09630_ _09763_ vssd1 vssd1 vccd1 vccd1 _09764_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_198_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20675__112 clknet_1_1__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__inv_2
XFILLER_0_186_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18432_ _02459_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15644_ _08486_ _08493_ _08717_ _08718_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__o31a_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05201_ _05998_ _06007_ net73 _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__a221o_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _04959_ _04971_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nor3_2
X_18363_ net4489 net4393 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _08562_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__and2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nor2_2
X_17314_ _10314_ _10313_ vssd1 vssd1 vccd1 vccd1 _10315_ sky130_fd_sc_hd__and2b_1
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14526_ _07675_ _07676_ _07623_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__a21o_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _02336_ net4475 _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
X_11738_ _04880_ _04905_ net4093 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ _10244_ _10245_ vssd1 vssd1 vccd1 vccd1 _10246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03983_ _03983_ vssd1 vssd1 vccd1 vccd1 clknet_0__03983_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14457_ _07606_ _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11669_ _04836_ net3893 _04837_ _04776_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13408_ _06545_ _06558_ _06540_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a21o_1
X_17176_ _10171_ _10175_ _10176_ vssd1 vssd1 vccd1 vccd1 _10178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14388_ _07483_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ _09192_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__xnor2_1
X_13339_ net6278 _06430_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16058_ _08490_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__clkbuf_4
Xhold3108 _00427_ vssd1 vssd1 vccd1 vccd1 net3632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3119 _03786_ vssd1 vssd1 vccd1 vccd1 net3643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15009_ _08146_ _08147_ _08069_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__mux2_1
Xhold2407 net4739 vssd1 vssd1 vccd1 vccd1 net2931 sky130_fd_sc_hd__buf_1
Xhold2418 net6096 vssd1 vssd1 vccd1 vccd1 net2942 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2429 _03101_ vssd1 vssd1 vccd1 vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19817_ net3151 net3075 net3972 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__mux2_1
Xhold1706 net6036 vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1717 net6857 vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 rbzero.tex_g1\[48\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _04173_ vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19748_ net6055 _03394_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19679_ net3100 _03374_ net2488 _03371_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21710_ clknet_leaf_19_i_clk net2078 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ clknet_leaf_34_i_clk net1617 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21572_ clknet_leaf_4_i_clk net5261 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_10 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_21 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _08279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20523_ net3582 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_43 i_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 net4779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 _09284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 net3222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_98 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20454_ net888 net3651 _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5000 _00774_ vssd1 vssd1 vccd1 vccd1 net5524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5011 rbzero.spi_registers.texadd3\[6\] vssd1 vssd1 vccd1 vccd1 net5535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5022 rbzero.spi_registers.buf_vshift\[2\] vssd1 vssd1 vccd1 vccd1 net5546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20385_ net3636 net1222 _03782_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__mux2_1
Xhold5033 _01039_ vssd1 vssd1 vccd1 vccd1 net5557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5044 rbzero.pov.spi_buffer\[25\] vssd1 vssd1 vccd1 vccd1 net5568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5055 _00791_ vssd1 vssd1 vccd1 vccd1 net5579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4310 _01099_ vssd1 vssd1 vccd1 vccd1 net4834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22124_ net256 net2199 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold5066 rbzero.pov.spi_buffer\[20\] vssd1 vssd1 vccd1 vccd1 net5590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4321 _03674_ vssd1 vssd1 vccd1 vccd1 net4845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4332 rbzero.pov.spi_buffer\[67\] vssd1 vssd1 vccd1 vccd1 net4856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5077 _01048_ vssd1 vssd1 vccd1 vccd1 net5601 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_84_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold5088 _01038_ vssd1 vssd1 vccd1 vccd1 net5612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4343 rbzero.pov.spi_buffer\[72\] vssd1 vssd1 vccd1 vccd1 net4867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5099 net1337 vssd1 vssd1 vccd1 vccd1 net5623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4354 _00523_ vssd1 vssd1 vccd1 vccd1 net4878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3620 _00515_ vssd1 vssd1 vccd1 vccd1 net4144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4365 net1131 vssd1 vssd1 vccd1 vccd1 net4889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3631 rbzero.traced_texa\[10\] vssd1 vssd1 vccd1 vccd1 net4155 sky130_fd_sc_hd__dlygate4sd3_1
X_22055_ clknet_leaf_90_i_clk net3583 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4376 _06268_ vssd1 vssd1 vccd1 vccd1 net4900 sky130_fd_sc_hd__clkbuf_2
Xhold3642 net923 vssd1 vssd1 vccd1 vccd1 net4166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4387 _06203_ vssd1 vssd1 vccd1 vccd1 net4911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3653 _00517_ vssd1 vssd1 vccd1 vccd1 net4177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4398 net1249 vssd1 vssd1 vccd1 vccd1 net4922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3664 net685 vssd1 vssd1 vccd1 vccd1 net4188 sky130_fd_sc_hd__dlygate4sd3_1
X_21006_ net6347 net4945 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__xnor2_1
Xhold3675 net1143 vssd1 vssd1 vccd1 vccd1 net4199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2930 _03817_ vssd1 vssd1 vccd1 vccd1 net3454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2941 net5663 vssd1 vssd1 vccd1 vccd1 net3465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3686 net1216 vssd1 vssd1 vccd1 vccd1 net4210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2952 net1175 vssd1 vssd1 vccd1 vccd1 net3476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3697 net1015 vssd1 vssd1 vccd1 vccd1 net4221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2963 net5770 vssd1 vssd1 vccd1 vccd1 net3487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2974 _03936_ vssd1 vssd1 vccd1 vccd1 net3498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2985 _08286_ vssd1 vssd1 vccd1 vccd1 net3509 sky130_fd_sc_hd__buf_1
Xhold2996 _03865_ vssd1 vssd1 vccd1 vccd1 net3520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10971_ net2638 net6894 _04355_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ net13 net14 _05867_ _05869_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a32o_1
X_21908_ clknet_leaf_92_i_clk net5389 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap78 _07878_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_2
X_13690_ _06731_ _06840_ _06816_ _06719_ _06724_ _06717_ vssd1 vssd1 vccd1 vccd1 _06841_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xmax_cap89 _04167_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_4
XFILLER_0_210_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ net6349 _05785_ _05799_ _05802_ _05787_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a311o_2
XFILLER_0_210_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21839_ clknet_leaf_80_i_clk net4778 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ net4063 _08412_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ rbzero.tex_b1\[31\] rbzero.tex_b1\[30\] _05476_ vssd1 vssd1 vccd1 vccd1 _05737_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ _07445_ _07436_ _07459_ _07461_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11523_ rbzero.spi_registers.texadd3\[18\] rbzero.spi_registers.texadd1\[18\] rbzero.spi_registers.texadd0\[18\]
+ rbzero.spi_registers.texadd2\[18\] _04692_ _04693_ vssd1 vssd1 vccd1 vccd1 _04695_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _08359_ net7779 _08365_ _08311_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__a22o_2
XFILLER_0_110_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17030_ _06206_ _10036_ _10037_ vssd1 vssd1 vccd1 vccd1 _10038_ sky130_fd_sc_hd__o21ai_1
X_14242_ _07391_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11454_ net2982 net4909 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11385_ net6952 net2816 _04573_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__mux2_1
X_14173_ _07322_ _07323_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6290 net2433 vssd1 vssd1 vccd1 vccd1 net6814 sky130_fd_sc_hd__dlygate4sd3_1
X_13124_ _06271_ net3369 vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor2_1
X_18981_ net3922 net6217 net4902 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17932_ _01760_ _01961_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__nand2_1
X_13055_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__clkbuf_8
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ net694 _05130_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or2b_1
XFILLER_0_206_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17863_ _10259_ _09375_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19602_ net5201 _03325_ _03336_ _03330_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__o211a_1
X_16814_ _09731_ _09746_ _09883_ vssd1 vssd1 vccd1 vccd1 _09884_ sky130_fd_sc_hd__a21bo_1
X_17794_ _01698_ _01723_ _01721_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16745_ _09812_ _09814_ vssd1 vssd1 vccd1 vccd1 _09815_ sky130_fd_sc_hd__nand2_1
X_19533_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13957_ net555 net583 _07107_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19464_ net3075 net3151 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ net35 net34 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nor2_1
X_16676_ _09731_ _09746_ vssd1 vssd1 vccd1 vccd1 _09747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13888_ _07037_ _07038_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__and2_4
XFILLER_0_5_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15627_ _08701_ _08490_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__nand2_1
X_18415_ _02444_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ net1709 _03199_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or2_1
X_12839_ net31 net30 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18346_ net4485 net4353 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__nor2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _08320_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509_ _07474_ _07523_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__nor2_1
X_18277_ _02282_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15489_ _08353_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17228_ _10098_ _10099_ _10096_ vssd1 vssd1 vccd1 vccd1 _10229_ sky130_fd_sc_hd__a21oi_1
Xinput30 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_2
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 i_mode[1] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_6
XFILLER_0_141_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput52 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_8
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold803 net5657 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17159_ _10151_ _10160_ vssd1 vssd1 vccd1 vccd1 _10161_ sky130_fd_sc_hd__xor2_2
Xhold814 net5624 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 _01532_ vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold836 net3513 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold847 net5672 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 net5176 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
X_20170_ net3291 _03704_ _03707_ _03696_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__o211a_1
Xhold869 net7738 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2204 net7168 vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2215 _01431_ vssd1 vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2226 net7271 vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2237 _01498_ vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1503 net6871 vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2248 _04386_ vssd1 vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 net5842 vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 _01454_ vssd1 vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 _04425_ vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1536 net6795 vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1547 _03437_ vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 net6847 vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1569 rbzero.spi_registers.buf_texadd2\[13\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21624_ clknet_leaf_4_i_clk net5145 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20812__236 clknet_1_1__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__inv_2
XFILLER_0_168_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21555_ clknet_leaf_101_i_clk net1087 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20506_ _03880_ net3366 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21486_ clknet_leaf_15_i_clk net2678 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20437_ net3296 net1263 _03823_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11170_ net6443 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20368_ net3643 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4140 _00610_ vssd1 vssd1 vccd1 vccd1 net4664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4151 net3880 vssd1 vssd1 vccd1 vccd1 net4675 sky130_fd_sc_hd__clkbuf_2
X_22107_ net239 net2860 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4162 net7561 vssd1 vssd1 vccd1 vccd1 net4686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4173 _02674_ vssd1 vssd1 vccd1 vccd1 net4697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4184 rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 net4708 sky130_fd_sc_hd__clkbuf_2
Xhold3450 _03463_ vssd1 vssd1 vccd1 vccd1 net3974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4195 net3216 vssd1 vssd1 vccd1 vccd1 net4719 sky130_fd_sc_hd__buf_1
X_22038_ clknet_leaf_95_i_clk net3712 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3461 _02954_ vssd1 vssd1 vccd1 vccd1 net3985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3472 _04828_ vssd1 vssd1 vccd1 vccd1 net3996 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_209_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3483 _05445_ vssd1 vssd1 vccd1 vccd1 net4007 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3494 _03957_ vssd1 vssd1 vccd1 vccd1 net4018 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2760 net7535 vssd1 vssd1 vccd1 vccd1 net3284 sky130_fd_sc_hd__buf_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893__308 clknet_1_0__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__inv_2
Xhold2771 rbzero.pov.ready_buffer\[23\] vssd1 vssd1 vccd1 vccd1 net3295 sky130_fd_sc_hd__dlygate4sd3_1
X_14860_ _07966_ _07842_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__xnor2_2
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2782 _03874_ vssd1 vssd1 vccd1 vccd1 net3306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2793 net731 vssd1 vssd1 vccd1 vccd1 net3317 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13811_ _06928_ _06936_ _06926_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__a21bo_1
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _07774_ _07590_ _07937_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__o31a_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16530_ _09601_ _09368_ _08313_ vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__a21o_2
X_13742_ _06846_ net79 vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__xor2_2
XFILLER_0_202_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ net1697 net6582 _04344_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16461_ _09433_ _09435_ _09532_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__o21ai_1
X_13673_ _06717_ _06731_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__nand2_1
X_10885_ net2721 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__clkbuf_1
X_18200_ _02082_ _02156_ _02154_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a21oi_1
X_15412_ _06166_ _06427_ net4086 vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__mux2_1
X_19180_ net3146 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ net5 net4 vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nor2_2
XFILLER_0_183_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16392_ _09359_ _09360_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18131_ _02176_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15343_ net4300 net2935 _08383_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _04983_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__or2_1
X_20787__213 clknet_1_1__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__inv_2
X_18062_ _02088_ _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11506_ _04650_ _04675_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15274_ _08300_ _06492_ _08319_ net7510 vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__a211o_1
X_12486_ _05646_ _05648_ _05651_ _05034_ _05023_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17013_ _10022_ net4528 _09966_ vssd1 vssd1 vccd1 vccd1 _10023_ sky130_fd_sc_hd__mux2_1
X_14225_ _07328_ _07329_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ net4009 vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14156_ _07301_ _07306_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11368_ net7258 net6806 _04562_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13107_ _06185_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _07159_ _07237_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__nor2_1
X_18964_ net3019 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
X_11299_ net5817 net2289 _04529_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__mux2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__or2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _06183_ _06179_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__o21a_1
X_18895_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _02854_
+ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _01894_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17777_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nand2_1
X_14989_ net4393 net7437 _08027_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19516_ _02996_ _03275_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__or2_1
X_16728_ _09674_ _09797_ vssd1 vssd1 vccd1 vccd1 _09798_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16659_ _09593_ _09595_ vssd1 vssd1 vccd1 vccd1 _09730_ sky130_fd_sc_hd__nor2_1
X_19447_ net3075 net3151 _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19378_ net2020 _03199_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18329_ net4511 net4374 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21340_ clknet_leaf_42_i_clk net4175 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21271_ clknet_leaf_50_i_clk _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 net5563 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 net6356 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 net5546 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20222_ net1228 _03731_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__or2_1
Xhold633 _03487_ vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold644 net5565 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold655 net6418 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold666 net4272 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 net6414 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20153_ net3466 _03692_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__or2_1
Xhold688 _02490_ vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold699 net5411 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2001 net6895 vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2012 net5875 vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2023 net7021 vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
X_20084_ _02864_ _03581_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__or2_1
Xhold2034 _01550_ vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 net6591 vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2045 _04204_ vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2056 _01323_ vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 net6901 vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1322 _00942_ vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2067 net6295 vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1333 net5869 vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2078 net7180 vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2089 net7293 vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1344 net6739 vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 _01367_ vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1366 _01343_ vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1377 net6869 vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1388 net6284 vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 net7224 vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20736__167 clknet_1_1__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__inv_2
XFILLER_0_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ net2568 net6626 _04192_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21607_ clknet_leaf_20_i_clk net5631 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _05070_ vssd1 vssd1 vccd1 vccd1 _05508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21538_ clknet_leaf_28_i_clk net1722 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ net4090 _05369_ _05432_ _05439_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a211oi_1
X_21469_ clknet_leaf_0_i_clk net3098 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14010_ _06876_ _06869_ _06970_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__or3_1
X_11222_ net7054 net7201 _04492_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__mux2_1
X_11153_ net2450 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15961_ _08992_ _08998_ _09035_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__nand3_2
X_11084_ net2025 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
Xhold3280 rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 net3804 sky130_fd_sc_hd__clkbuf_4
X_17700_ net4433 net4593 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__nor2_1
Xhold3291 _01239_ vssd1 vssd1 vccd1 vccd1 net3815 sky130_fd_sc_hd__dlygate4sd3_1
X_14912_ net4456 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__clkbuf_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15892_ _08951_ _08966_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__nor2_1
X_18680_ _02646_ net3043 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__nand2_2
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2590 net7489 vssd1 vssd1 vccd1 vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _08872_ _08873_ _09484_ _09861_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14843_ _07991_ _07993_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__nand2_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17562_ _10558_ _10560_ vssd1 vssd1 vccd1 vccd1 _10561_ sky130_fd_sc_hd__xor2_2
X_14774_ _07232_ _07359_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ net3992 _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nand2_1
X_16513_ _09476_ _09480_ _09584_ vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19301_ net1912 _03147_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or2_1
X_13725_ net553 vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__buf_2
X_10937_ _04332_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__clkbuf_4
X_17493_ _10383_ _08708_ _10378_ _10381_ vssd1 vssd1 vccd1 vccd1 _10492_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_156_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16444_ _09413_ _09515_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__or2_1
X_19232_ net5743 _03106_ _03117_ _03115_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _06638_ _06687_ _06718_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__a21oi_1
X_10868_ net7237 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12607_ net4239 _05097_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a21o_1
X_19163_ net5513 _03065_ _03075_ _03074_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__o211a_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _09328_ _08331_ _08698_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__a2bb2o_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13587_ _06552_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__inv_2
X_10799_ net2760 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__clkbuf_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18114_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15326_ net2935 _08341_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12538_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _05541_ vssd1 vssd1 vccd1 vccd1 _05703_
+ sky130_fd_sc_hd__mux2_1
X_19094_ _04881_ _05816_ _03032_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__and4_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _02091_ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15257_ _08318_ _08326_ _08331_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__or3_2
XFILLER_0_112_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12469_ _05633_ _05634_ _05069_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14208_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__clkbuf_4
Xhold4909 _01086_ vssd1 vssd1 vccd1 vccd1 net5433 sky130_fd_sc_hd__dlygate4sd3_1
X_15188_ net4575 _08188_ net4933 vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ _07288_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19996_ net4561 _03582_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20841__262 clknet_1_0__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__inv_2
X_18947_ _02922_ _02923_ _02928_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18878_ _02864_ rbzero.wall_tracer.rayAddendY\[3\] _02860_ vssd1 vssd1 vccd1 vccd1
+ _02865_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17829_ _10383_ _09420_ _01766_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_179_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22441_ clknet_leaf_39_i_clk net4707 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold6801 rbzero.color_floor\[1\] vssd1 vssd1 vccd1 vccd1 net7325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22372_ net504 net2829 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6823 rbzero.pov.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 net7347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6834 rbzero.spi_registers.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 net7358 sky130_fd_sc_hd__dlygate4sd3_1
X_21323_ clknet_leaf_55_i_clk _00492_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6845 rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 net7369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6856 net4294 vssd1 vssd1 vccd1 vccd1 net7380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6878 _08338_ vssd1 vssd1 vccd1 vccd1 net7402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21254_ clknet_leaf_52_i_clk net3049 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold430 _03680_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold441 net5315 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 net5347 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold463 net5150 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20205_ net3665 _03718_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21185_ _02532_ net4657 net4425 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold474 net5423 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold485 net5448 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold496 net4289 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
X_20136_ net5251 _03679_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__or2_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ _03616_ net3675 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__or2_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _00878_ vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 net6605 vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 _01353_ vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _03433_ vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 _04354_ vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 net6693 vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _00938_ vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _05009_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__buf_4
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ net1010 net1650 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _06626_ _06649_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__nor2_2
X_10722_ net2700 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _07638_ _07640_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__xor2_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ net4947 _06489_ _06491_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__a21o_1
X_10653_ net2225 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16160_ _08621_ _08637_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__nand2_1
X_13372_ _06435_ _06474_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__nand3_1
XFILLER_0_134_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ _08218_ net3055 net4784 _08215_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__o211a_1
X_12323_ _05471_ _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16091_ _09125_ _09147_ _09165_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _08092_ net7836 vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12254_ net3880 _05347_ _05351_ net3893 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11205_ net7097 net2173 _04481_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19850_ net3258 _08364_ _03484_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
X_20899__314 clknet_1_1__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__inv_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12185_ _04604_ _04812_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__nand2_1
X_18801_ _02789_ _02793_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__xnor2_1
X_11136_ net7111 net6792 _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__mux2_1
X_19781_ net3096 _03427_ net1745 _03441_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__o211a_1
X_16993_ _10004_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__clkbuf_1
X_18732_ net3881 _09987_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__o21ai_1
X_11067_ net6680 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
X_15944_ _08958_ _08960_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15875_ _08907_ _08912_ _08926_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__a21o_1
X_18663_ _02654_ _02669_ _02667_ _04623_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a31o_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _01664_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14826_ _07972_ _07693_ _07974_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18594_ net7602 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__inv_2
Xclkbuf_0__04002_ _04002_ vssd1 vssd1 vccd1 vccd1 clknet_0__04002_ sky130_fd_sc_hd__clkbuf_16
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _10540_ _10543_ vssd1 vssd1 vccd1 vccd1 _10544_ sky130_fd_sc_hd__xnor2_1
X_14757_ _07886_ _07901_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11969_ net1600 _05124_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13708_ net573 vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17476_ _09447_ _09794_ _10474_ vssd1 vssd1 vccd1 vccd1 _10475_ sky130_fd_sc_hd__a21oi_1
X_20871__288 clknet_1_1__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__inv_2
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14688_ _07796_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19215_ net5721 _03106_ _03108_ _03096_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__o211a_1
X_16427_ _09495_ _09499_ _09377_ _09378_ _09362_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13639_ _06744_ _06745_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ _09429_ _09430_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19146_ _03039_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__buf_2
Xhold6108 net1777 vssd1 vssd1 vccd1 vccd1 net6632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6119 _04216_ vssd1 vssd1 vccd1 vccd1 net6643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15309_ net4338 _08362_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__nand2_1
Xhold5407 net1941 vssd1 vssd1 vccd1 vccd1 net5931 sky130_fd_sc_hd__dlygate4sd3_1
X_16289_ net3273 _06211_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19077_ net4322 net2979 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__or2_1
Xhold5418 net5804 vssd1 vssd1 vccd1 vccd1 net5942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5429 net1970 vssd1 vssd1 vccd1 vccd1 net5953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4706 net876 vssd1 vssd1 vccd1 vccd1 net5230 sky130_fd_sc_hd__dlygate4sd3_1
X_18028_ _01974_ _01977_ _01975_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4717 _01081_ vssd1 vssd1 vccd1 vccd1 net5241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4728 _01042_ vssd1 vssd1 vccd1 vccd1 net5252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4739 net989 vssd1 vssd1 vccd1 vccd1 net5263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20765__193 clknet_1_1__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__inv_2
XFILLER_0_22_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19979_ rbzero.debug_overlay.facingX\[-6\] _03582_ vssd1 vssd1 vccd1 vccd1 _03586_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21941_ net166 net1523 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
X_21872_ clknet_leaf_100_i_clk net1205 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7310 rbzero.wall_tracer.stepDistX\[-9\] vssd1 vssd1 vccd1 vccd1 net7834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7321 rbzero.row_render.size\[3\] vssd1 vssd1 vccd1 vccd1 net7845 sky130_fd_sc_hd__dlygate4sd3_1
X_22424_ clknet_leaf_54_i_clk net5170 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6620 rbzero.tex_g1\[5\] vssd1 vssd1 vccd1 vccd1 net7144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22355_ net487 net2755 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold6631 net2364 vssd1 vssd1 vccd1 vccd1 net7155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7376 rbzero.texu_hot\[0\] vssd1 vssd1 vccd1 vccd1 net7900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6642 rbzero.tex_g1\[59\] vssd1 vssd1 vccd1 vccd1 net7166 sky130_fd_sc_hd__dlygate4sd3_1
X_20848__268 clknet_1_1__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__inv_2
Xhold6653 net2781 vssd1 vssd1 vccd1 vccd1 net7177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6664 _04516_ vssd1 vssd1 vccd1 vccd1 net7188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5930 _04240_ vssd1 vssd1 vccd1 vccd1 net6454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6675 net2732 vssd1 vssd1 vccd1 vccd1 net7199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21306_ clknet_leaf_74_i_clk net3911 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold5941 net1352 vssd1 vssd1 vccd1 vccd1 net6465 sky130_fd_sc_hd__dlygate4sd3_1
X_22286_ net418 net2059 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
Xhold6686 rbzero.tex_b0\[19\] vssd1 vssd1 vccd1 vccd1 net7210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5952 rbzero.tex_b0\[30\] vssd1 vssd1 vccd1 vccd1 net6476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6697 net2559 vssd1 vssd1 vccd1 vccd1 net7221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5963 net1446 vssd1 vssd1 vccd1 vccd1 net6487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5974 _09944_ vssd1 vssd1 vccd1 vccd1 net6498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5985 _04569_ vssd1 vssd1 vccd1 vccd1 net6509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 net5039 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
X_21237_ clknet_leaf_71_i_clk _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5996 net1448 vssd1 vssd1 vccd1 vccd1 net6520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 net4216 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net5043 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__05942_ clknet_0__05942_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05942_
+ sky130_fd_sc_hd__clkbuf_16
Xhold293 net5098 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
X_21168_ _09933_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20119_ net4838 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__clkbuf_4
X_21099_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__inv_2
X_13990_ _07139_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12941_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__nor2_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15660_ _08733_ _08734_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__xnor2_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _04161_ net3993 net28 vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__mux2_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _07647_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__nand2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _04992_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__clkbuf_8
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _08664_ _08643_ _08540_ _08665_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__and4bb_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _09987_ _10211_ _10212_ _10330_ vssd1 vssd1 vccd1 vccd1 _10331_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _07641_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__and2_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ net757 net2194 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__or2_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _10257_ _08708_ _10261_ vssd1 vssd1 vccd1 vccd1 _10262_ sky130_fd_sc_hd__or3_1
X_10705_ net2828 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__clkbuf_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ _07618_ _07464_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ _04853_ net2987 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19000_ net3891 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16212_ net4355 net7370 _08293_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__mux2_1
X_13424_ _06545_ _06574_ _06540_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a21o_1
X_17192_ _09829_ _09897_ _10193_ vssd1 vssd1 vccd1 vccd1 _10194_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_181_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10636_ net2603 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _09086_ _08582_ _09216_ _08584_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ _06438_ _06444_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ _05248_ _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20907__321 clknet_1_0__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__inv_2
X_16074_ _09137_ _09142_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13286_ _06435_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15025_ _08161_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
X_19902_ _08279_ net3158 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__and2_1
X_12237_ net3837 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__clkbuf_1
X_19833_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__buf_2
X_12168_ _05324_ net4072 vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__and2_1
XFILLER_0_209_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ net6966 net2271 _04437_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux2_1
X_19764_ net6694 _03429_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__or2_1
X_12099_ _05235_ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__or2_1
X_16976_ net4568 net4566 vssd1 vssd1 vccd1 vccd1 _09989_ sky130_fd_sc_hd__or2_1
X_18715_ _02692_ _02704_ _02702_ _02686_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__o211a_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15927_ _08999_ _09000_ _09001_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__a21boi_2
Xinput6 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19695_ net6043 _03361_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18646_ _02653_ _02654_ _02627_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a21oi_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _08929_ _08930_ _08932_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__nand3_1
XFILLER_0_204_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20953__363 clknet_1_0__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__inv_2
X_14809_ _07954_ _07956_ _07958_ _07959_ _07915_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__o2111a_1
X_18577_ net6237 _05403_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15789_ _08448_ _08450_ _08457_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17528_ _10507_ _10508_ _10525_ vssd1 vssd1 vccd1 vccd1 _10527_ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17459_ net4501 net4417 vssd1 vssd1 vccd1 vccd1 _10458_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20470_ _03836_ net3696 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19129_ net5999 _03052_ _03056_ _03048_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5204 net1083 vssd1 vssd1 vccd1 vccd1 net5728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5215 rbzero.spi_registers.texadd0\[0\] vssd1 vssd1 vccd1 vccd1 net5739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22140_ net272 net2178 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
Xhold5226 net1618 vssd1 vssd1 vccd1 vccd1 net5750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5237 rbzero.spi_registers.buf_texadd2\[23\] vssd1 vssd1 vccd1 vccd1 net5761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5248 rbzero.spi_registers.vshift\[0\] vssd1 vssd1 vccd1 vccd1 net5772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4503 _00736_ vssd1 vssd1 vccd1 vccd1 net5027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5259 net1634 vssd1 vssd1 vccd1 vccd1 net5783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4514 net783 vssd1 vssd1 vccd1 vccd1 net5038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4525 net1274 vssd1 vssd1 vccd1 vccd1 net5049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4536 rbzero.spi_registers.buf_texadd0\[16\] vssd1 vssd1 vccd1 vccd1 net5060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22071_ clknet_leaf_13_i_clk net3755 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3802 net796 vssd1 vssd1 vccd1 vccd1 net4326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4547 rbzero.spi_registers.buf_texadd0\[1\] vssd1 vssd1 vccd1 vccd1 net5071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4558 rbzero.spi_registers.texadd1\[14\] vssd1 vssd1 vccd1 vccd1 net5082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3813 net735 vssd1 vssd1 vccd1 vccd1 net4337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3824 net7479 vssd1 vssd1 vccd1 vccd1 net4348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4569 net791 vssd1 vssd1 vccd1 vccd1 net5093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21022_ _04024_ _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__or2b_1
Xhold3835 _00977_ vssd1 vssd1 vccd1 vccd1 net4359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3846 net3102 vssd1 vssd1 vccd1 vccd1 net4370 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3857 net7780 vssd1 vssd1 vccd1 vccd1 net4381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3868 net7450 vssd1 vssd1 vccd1 vccd1 net4392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3879 net3155 vssd1 vssd1 vccd1 vccd1 net4403 sky130_fd_sc_hd__buf_1
XFILLER_0_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21924_ clknet_leaf_6_i_clk net1317 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ clknet_leaf_97_i_clk net4462 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21786_ clknet_leaf_10_i_clk net4337 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7140 rbzero.spi_registers.buf_texadd1\[17\] vssd1 vssd1 vccd1 vccd1 net7664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22407_ net159 net2573 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
Xhold7151 rbzero.spi_registers.texadd2\[14\] vssd1 vssd1 vccd1 vccd1 net7675 sky130_fd_sc_hd__dlygate4sd3_1
X_20599_ net2938 _03782_ net3562 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_104_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6450 net2286 vssd1 vssd1 vccd1 vccd1 net6974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ net3851 _06279_ _06270_ _06280_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6461 rbzero.tex_g1\[14\] vssd1 vssd1 vccd1 vccd1 net6985 sky130_fd_sc_hd__dlygate4sd3_1
X_22338_ net470 net1426 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
Xhold6472 net2551 vssd1 vssd1 vccd1 vccd1 net6996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6483 _04189_ vssd1 vssd1 vccd1 vccd1 net7007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6494 net1932 vssd1 vssd1 vccd1 vccd1 net7018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5760 rbzero.spi_registers.buf_texadd1\[9\] vssd1 vssd1 vccd1 vccd1 net6284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13071_ net4896 vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__inv_2
X_22269_ net401 net2463 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5771 _03271_ vssd1 vssd1 vccd1 vccd1 net6295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5782 rbzero.spi_registers.mosi vssd1 vssd1 vccd1 vccd1 net6306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5793 _04422_ vssd1 vssd1 vccd1 vccd1 net6317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12022_ net4033 _04831_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16830_ _09898_ _09899_ vssd1 vssd1 vccd1 vccd1 _09900_ sky130_fd_sc_hd__xor2_2
XFILLER_0_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16761_ _09719_ _09724_ vssd1 vssd1 vccd1 vccd1 _09831_ sky130_fd_sc_hd__or2_1
X_13973_ _06861_ _06837_ _06918_ _06895_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o22ai_1
X_18500_ _02513_ _02517_ _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__or3_1
X_15712_ _08777_ _08785_ _08786_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__a21oi_2
X_12924_ _04162_ _06065_ _06066_ net3993 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a22o_1
X_16692_ _09627_ _09629_ vssd1 vssd1 vccd1 vccd1 _09763_ sky130_fd_sc_hd__nor2_1
X_19480_ net1726 net3116 net3077 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18431_ _02458_ net4573 _02411_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
X_15643_ _08472_ _08485_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ net52 _06012_ _06008_ net51 vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a22o_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _04933_ _04958_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__and2_1
X_15574_ _08551_ _08561_ _08558_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__a21bo_1
X_18362_ net4489 net4393 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12786_ net25 net24 vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nor2_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17313_ _10310_ _10312_ vssd1 vssd1 vccd1 vccd1 _10314_ sky130_fd_sc_hd__nand2_1
X_14525_ _07083_ _06922_ _07463_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__or3_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11737_ net4092 _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18293_ net4920 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03982_ _03982_ vssd1 vssd1 vccd1 vccd1 clknet_0__03982_ sky130_fd_sc_hd__clkbuf_16
X_17244_ _10108_ _10112_ _10113_ _10115_ _10107_ vssd1 vssd1 vccd1 vccd1 _10245_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_127_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ _07366_ _07353_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__nor2_1
X_11668_ net4033 net3880 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ net6150 _06431_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17175_ _10171_ _10175_ _10176_ vssd1 vssd1 vccd1 vccd1 _10177_ sky130_fd_sc_hd__nand3_2
X_10619_ net6518 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__clkbuf_1
X_14387_ _07481_ _07482_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11599_ rbzero.spi_registers.texadd0\[0\] _04680_ _04769_ _04770_ _04159_ vssd1 vssd1
+ vccd1 vccd1 _04771_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _09199_ _09200_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__nor2_1
X_13338_ _06486_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16057_ _09094_ _09131_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__mux2_4
Xhold3109 net682 vssd1 vssd1 vccd1 vccd1 net3633 sky130_fd_sc_hd__clkbuf_2
X_15008_ _06690_ _07989_ _08002_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__a21o_1
Xhold2408 net4741 vssd1 vssd1 vccd1 vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2419 net7733 vssd1 vssd1 vccd1 vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
X_19816_ net3153 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1707 net6038 vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1718 _01414_ vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1729 net932 vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19747_ net4322 _03392_ net1538 _03413_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__o211a_1
X_16959_ _09946_ _09947_ _09974_ _09967_ vssd1 vssd1 vccd1 vccd1 _09975_ sky130_fd_sc_hd__and4_1
XFILLER_0_212_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20877__294 clknet_1_0__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__inv_2
X_19678_ net7195 _03375_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18629_ _02637_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02639_
+ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_3_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21640_ clknet_leaf_29_i_clk net3080 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21571_ clknet_leaf_17_i_clk net4126 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_11 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _08873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20522_ _03880_ net3581 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__and2_1
XANTENNA_44 rbzero.wall_tracer.visualWallDist\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_55 net6146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_66 _10454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_77 net4090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20453_ net3250 vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_99 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5001 net1119 vssd1 vssd1 vccd1 vccd1 net5525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5012 net1194 vssd1 vssd1 vccd1 vccd1 net5536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5023 net1146 vssd1 vssd1 vccd1 vccd1 net5547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20384_ net3430 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
Xhold5034 rbzero.map_overlay.i_mapdx\[5\] vssd1 vssd1 vccd1 vccd1 net5558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4300 _06201_ vssd1 vssd1 vccd1 vccd1 net4824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5045 _01061_ vssd1 vssd1 vccd1 vccd1 net5569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22123_ net255 net1385 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold4311 net1210 vssd1 vssd1 vccd1 vccd1 net4835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5056 net1262 vssd1 vssd1 vccd1 vccd1 net5580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5067 net1280 vssd1 vssd1 vccd1 vccd1 net5591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4322 _01102_ vssd1 vssd1 vccd1 vccd1 net4846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5078 rbzero.pov.spi_buffer\[21\] vssd1 vssd1 vccd1 vccd1 net5602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4333 _01103_ vssd1 vssd1 vccd1 vccd1 net4857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5089 rbzero.spi_registers.texadd1\[13\] vssd1 vssd1 vccd1 vccd1 net5613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4344 net1508 vssd1 vssd1 vccd1 vccd1 net4868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3610 _00518_ vssd1 vssd1 vccd1 vccd1 net4134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4355 net2808 vssd1 vssd1 vccd1 vccd1 net4879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3621 net653 vssd1 vssd1 vccd1 vccd1 net4145 sky130_fd_sc_hd__dlygate4sd3_1
X_22054_ clknet_leaf_90_i_clk net3278 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4366 gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 net4890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3632 net7555 vssd1 vssd1 vccd1 vccd1 net4156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4377 _09963_ vssd1 vssd1 vccd1 vccd1 net4901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3643 net7644 vssd1 vssd1 vccd1 vccd1 net4167 sky130_fd_sc_hd__buf_1
Xhold4388 net6269 vssd1 vssd1 vccd1 vccd1 net4912 sky130_fd_sc_hd__buf_1
Xhold3654 net679 vssd1 vssd1 vccd1 vccd1 net4178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4399 _00525_ vssd1 vssd1 vccd1 vccd1 net4923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3665 net7711 vssd1 vssd1 vccd1 vccd1 net4189 sky130_fd_sc_hd__dlygate4sd3_1
X_21005_ net4945 net65 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nor2_1
Xhold2931 _03818_ vssd1 vssd1 vccd1 vccd1 net3455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3676 net7717 vssd1 vssd1 vccd1 vccd1 net4200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2942 net1177 vssd1 vssd1 vccd1 vccd1 net3466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3687 net7657 vssd1 vssd1 vccd1 vccd1 net4211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2953 _03916_ vssd1 vssd1 vccd1 vccd1 net3477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3698 rbzero.spi_registers.buf_texadd1\[16\] vssd1 vssd1 vccd1 vccd1 net4222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2964 net1247 vssd1 vssd1 vccd1 vccd1 net3488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2975 _01244_ vssd1 vssd1 vccd1 vccd1 net3499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2986 _08291_ vssd1 vssd1 vccd1 vccd1 net3510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2997 _03866_ vssd1 vssd1 vccd1 vccd1 net3521 sky130_fd_sc_hd__dlygate4sd3_1
X_10970_ net2766 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21907_ clknet_leaf_92_i_clk net1492 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ _04241_ _05785_ _05796_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a31o_2
XFILLER_0_183_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21838_ clknet_leaf_81_i_clk net3546 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _05476_ vssd1 vssd1 vccd1 vccd1 _05736_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21769_ clknet_leaf_4_i_clk net1720 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _07391_ _07434_ _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ rbzero.spi_registers.texadd3\[17\] rbzero.spi_registers.texadd1\[17\] rbzero.spi_registers.texadd0\[17\]
+ rbzero.spi_registers.texadd2\[17\] _04692_ _04693_ vssd1 vssd1 vccd1 vccd1 _04694_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15290_ _08364_ _08361_ _08341_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14241_ _07337_ _07363_ _07390_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ net4909 net2982 _04626_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_34_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14172_ _07310_ _07321_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11384_ net2512 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6280 net2277 vssd1 vssd1 vccd1 vccd1 net6804 sky130_fd_sc_hd__dlygate4sd3_1
X_13123_ net3852 vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__inv_2
Xhold6291 _04471_ vssd1 vssd1 vccd1 vccd1 net6815 sky130_fd_sc_hd__dlygate4sd3_1
X_18980_ net3921 _02956_ _09999_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _01958_ _01960_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__or2_1
X_13054_ _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__clkbuf_8
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5590 net1566 vssd1 vssd1 vccd1 vccd1 net6114 sky130_fd_sc_hd__dlygate4sd3_1
X_12005_ net3992 _05153_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__o21a_2
XFILLER_0_178_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17862_ _01831_ _01824_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19601_ net3050 _03327_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__or2_1
X_16813_ _09743_ _09745_ vssd1 vssd1 vccd1 vccd1 _09883_ sky130_fd_sc_hd__nand2_1
X_17793_ _01823_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__xnor2_1
X_19532_ _08274_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__clkbuf_4
X_16744_ _08707_ _09813_ _08962_ vssd1 vssd1 vccd1 vccd1 _09814_ sky130_fd_sc_hd__or3b_1
X_13956_ _07102_ net535 vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__and2b_1
X_19463_ net1727 _03241_ net1791 _03233_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__o211a_1
X_12907_ _06059_ _06060_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__a21o_2
X_16675_ _09743_ _09745_ vssd1 vssd1 vccd1 vccd1 _09746_ sky130_fd_sc_hd__xor2_1
X_13887_ _07030_ _07025_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18414_ _02443_ net4458 _02411_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ _08328_ _08329_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__nor2_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ net32 net33 vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nor2_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ net5147 _03198_ _03209_ _03207_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18345_ _02375_ _02376_ _02377_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__o21a_1
X_15557_ _06208_ _08631_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__nand2_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _05927_ _05928_ net19 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ _07657_ _07658_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__nand2_2
X_15488_ _08353_ _08405_ _08424_ _08557_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__or4_1
X_18276_ _02287_ _02321_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17227_ _10226_ _10227_ vssd1 vssd1 vccd1 vccd1 _10228_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput20 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput31 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_4
X_14439_ _07589_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__clkbuf_4
Xinput42 i_mode[2] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_4
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_8
XFILLER_0_141_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17158_ _10154_ _10159_ vssd1 vssd1 vccd1 vccd1 _10160_ sky130_fd_sc_hd__xor2_2
Xhold804 net3816 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 net3842 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold826 net5668 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 _01104_ vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 net6424 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _08836_ _08946_ _09181_ _09183_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17089_ _09826_ _10088_ _10089_ vssd1 vssd1 vccd1 vccd1 _10091_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold859 net6503 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2205 net7170 vssd1 vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2216 net7273 vssd1 vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2227 _04180_ vssd1 vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2238 rbzero.tex_g1\[50\] vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1504 net6873 vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _01394_ vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 _01268_ vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1526 _01359_ vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1537 _04282_ vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1548 net6165 vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _04196_ vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21623_ clknet_leaf_5_i_clk net5864 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21554_ clknet_leaf_101_i_clk net918 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20505_ net3365 net1290 _03867_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21485_ clknet_leaf_93_i_clk net2124 vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20436_ net3758 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20367_ _08279_ net3642 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4130 _01606_ vssd1 vssd1 vccd1 vccd1 net4654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22106_ net238 net2321 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold4141 net3482 vssd1 vssd1 vccd1 vccd1 net4665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4152 _00980_ vssd1 vssd1 vccd1 vccd1 net4676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4163 net3852 vssd1 vssd1 vccd1 vccd1 net4687 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4174 _00588_ vssd1 vssd1 vccd1 vccd1 net4698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3440 net6286 vssd1 vssd1 vccd1 vccd1 net3964 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4185 _02818_ vssd1 vssd1 vccd1 vccd1 net4709 sky130_fd_sc_hd__dlygate4sd3_1
X_22037_ clknet_leaf_95_i_clk net3767 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3451 net6313 vssd1 vssd1 vccd1 vccd1 net3975 sky130_fd_sc_hd__clkbuf_1
Xhold3462 _00617_ vssd1 vssd1 vccd1 vccd1 net3986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3473 _02948_ vssd1 vssd1 vccd1 vccd1 net3997 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3484 _00458_ vssd1 vssd1 vccd1 vccd1 net4008 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2750 net5449 vssd1 vssd1 vccd1 vccd1 net3274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3495 _01254_ vssd1 vssd1 vccd1 vccd1 net4019 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2761 rbzero.pov.ready_buffer\[54\] vssd1 vssd1 vccd1 vccd1 net3285 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2772 net713 vssd1 vssd1 vccd1 vccd1 net3296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2783 _03875_ vssd1 vssd1 vccd1 vccd1 net3307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2794 _03804_ vssd1 vssd1 vccd1 vccd1 net3318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _06952_ _06960_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__xnor2_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _07938_ _07940_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13741_ _06887_ _06891_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__and2_1
X_10953_ net2235 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16460_ _09421_ _09436_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ _06657_ _06705_ _06733_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ net6916 net2747 _04236_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15411_ _08472_ _08485_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__xnor2_1
X_12623_ net7 net6 vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__nor2_2
X_16391_ _09352_ _09354_ _09351_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20346__78 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18130_ _01833_ _02084_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15342_ net4300 net7404 vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__nand2_1
X_12554_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _04994_ vssd1 vssd1 vccd1 vccd1 _05719_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ _04648_ _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18061_ _02090_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__xnor2_1
X_15273_ net4086 _06152_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nor2_1
X_12485_ _05649_ _05650_ _05002_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17012_ _10018_ _10020_ _10021_ vssd1 vssd1 vccd1 vccd1 _10022_ sky130_fd_sc_hd__o21ai_1
X_14224_ _07264_ _07265_ _07318_ _07319_ net568 vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__a32o_1
XFILLER_0_184_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11436_ net4009 _04607_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ _07302_ _07305_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__nor2_1
X_11367_ net6510 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13106_ _06186_ net3804 _06183_ net4821 vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__or4_1
X_14086_ _07204_ _07206_ _07208_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__o21a_1
X_18963_ net3018 _02943_ _02714_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11298_ net5955 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _10581_ _01855_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a21oi_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ net3804 _06178_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a21o_1
X_18894_ _02860_ _02862_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17845_ _10379_ _09310_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17776_ _09108_ _10406_ _01711_ _10539_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14988_ _08127_ _08108_ _08129_ net7436 net6162 vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__a221o_4
XFILLER_0_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19515_ net5406 _03274_ _03283_ _03280_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__o211a_1
X_16727_ _09051_ _09662_ vssd1 vssd1 vccd1 vccd1 _09797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13939_ _06861_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19446_ net4326 _03238_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__nand2_1
X_16658_ _09727_ _09728_ vssd1 vssd1 vccd1 vccd1 _09729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_83_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15609_ _08444_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_173_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19377_ net5504 _03198_ _03200_ _03194_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16589_ _09561_ _09579_ _09659_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18328_ _02363_ _02361_ _02362_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18259_ _02303_ _02304_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21270_ clknet_leaf_56_i_clk _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold601 net3584 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 _04157_ vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 net5548 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
X_20221_ net5212 _03730_ _03736_ _03735_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__o211a_1
Xhold634 net4307 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold645 net5567 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03779_ clknet_0__03779_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03779_
+ sky130_fd_sc_hd__clkbuf_16
Xhold656 _04208_ vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold667 net6448 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_21_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold678 net6416 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
X_20152_ net3466 _03691_ _03697_ _03696_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold689 _00573_ vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2002 _01416_ vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2013 net5877 vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2024 net7023 vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ net3317 _03577_ net4635 _03636_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__o211a_1
Xhold2035 net7220 vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _04553_ vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 _01556_ vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 net6887 vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 _04174_ vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2068 net6296 vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 net6721 vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _01308_ vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2079 _04184_ vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1345 _03399_ vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1356 net6757 vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1367 net6625 vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1378 _01531_ vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1389 _03373_ vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21606_ clknet_leaf_20_i_clk net5489 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21537_ clknet_leaf_27_i_clk net1828 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ _05433_ _05434_ _05436_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__or4_1
X_21468_ clknet_leaf_24_i_clk net3053 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11221_ net6495 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
X_20419_ _03814_ net3324 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__and2_1
X_21399_ clknet_leaf_64_i_clk _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11152_ net2449 net53 _04377_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20654__93 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__inv_2
X_20901__316 clknet_1_1__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__inv_2
X_15960_ _09009_ _09033_ _09034_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__a21o_1
X_11083_ net2024 net6316 _04415_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3270 net4973 vssd1 vssd1 vccd1 vccd1 net3794 sky130_fd_sc_hd__dlygate4sd3_1
X_14911_ net4455 _08059_ _08027_ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__mux2_1
Xhold3281 net6189 vssd1 vssd1 vccd1 vccd1 net3805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3292 net5556 vssd1 vssd1 vccd1 vccd1 net3816 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _08955_ _08956_ _08965_ _08964_ _08957_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__o32a_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2580 net3939 vssd1 vssd1 vccd1 vccd1 net3104 sky130_fd_sc_hd__dlygate4sd3_1
X_17630_ _01680_ _01681_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__and2_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _07984_ _07992_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__xnor2_4
Xhold2591 net7817 vssd1 vssd1 vccd1 vccd1 net3115 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1890 _01289_ vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ _10375_ _10436_ _10559_ vssd1 vssd1 vccd1 vccd1 _10560_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14773_ _07618_ _07590_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__nor2_1
X_11985_ net2869 _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19300_ net4995 _03146_ _03156_ _03155_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__o211a_1
X_16512_ _09478_ _09479_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__nand2_1
X_10936_ net2675 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13724_ _06869_ _06867_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__or2_1
X_17492_ _10489_ _10490_ vssd1 vssd1 vccd1 vccd1 _10491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19231_ net5236 _03107_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16443_ _09413_ _09515_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__nand2_1
X_10867_ net7235 net2682 _04299_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__mux2_1
X_13655_ _06589_ _06799_ _06805_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_186_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ net4239 _05097_ _05209_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__o21ai_1
X_19162_ net2541 _03066_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__or2_1
X_16374_ _08962_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__buf_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _06736_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10798_ net7207 net6578 _04266_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__mux2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18113_ _01984_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__xnor2_1
X_12537_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _04989_ vssd1 vssd1 vccd1 vccd1 _05702_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15325_ net3262 _08399_ _08303_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19093_ net3937 net3930 net4002 _04802_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and4b_1
XFILLER_0_186_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18044_ _02023_ _02020_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12468_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _05072_ vssd1 vssd1 vccd1 vccd1 _05634_
+ sky130_fd_sc_hd__mux2_1
X_15256_ _08330_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11419_ net5769 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
X_14207_ _07307_ _07357_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__nand2_2
X_15187_ _08272_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
X_12399_ _05000_ _05561_ _05565_ _05023_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14138_ _07008_ _07261_ _07287_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__or3_1
X_19995_ net3788 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ _07217_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__or2_1
X_18946_ _02913_ _02917_ _02927_ _04623_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18877_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17828_ _01822_ _01799_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__or2b_1
XFILLER_0_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _01684_ _10407_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19429_ net5018 _03224_ _03229_ _03220_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22440_ clknet_leaf_39_i_clk net4681 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20325__59 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22371_ net503 net2733 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6802 _03097_ vssd1 vssd1 vccd1 vccd1 net7326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6813 _03603_ vssd1 vssd1 vccd1 vccd1 net7337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21322_ clknet_leaf_72_i_clk _00491_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6835 rbzero.spi_registers.spi_counter\[0\] vssd1 vssd1 vccd1 vccd1 net7359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6846 net4335 vssd1 vssd1 vccd1 vccd1 net7370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6857 _09404_ vssd1 vssd1 vccd1 vccd1 net7381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6879 _08339_ vssd1 vssd1 vccd1 vccd1 net7403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold420 net5276 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21253_ clknet_leaf_52_i_clk net3068 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold431 net5599 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold442 net5341 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold453 net5419 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
X_20204_ net3665 _03717_ _03726_ _03722_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__o211a_1
Xhold464 net5152 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
X_21184_ _02529_ net4425 _04143_ _02528_ net701 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a32o_1
Xhold475 net5425 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold486 net7498 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold497 net5401 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20135_ net5251 _03676_ _03687_ _03683_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__o211a_1
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ net4799 net3674 _03580_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__mux2_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 net6065 vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 net5794 vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _01486_ vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 net6703 vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 _00928_ vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 _01423_ vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _03432_ vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1197 net5787 vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _04936_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20968_ clknet_1_0__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__buf_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ net6445 net2699 _04225_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13440_ _06495_ _06590_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_181_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10652_ net6688 net6782 _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13371_ _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ _04978_ _05475_ _05480_ _05489_ _05027_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__o311a_1
X_15110_ net4783 _08223_ vssd1 vssd1 vccd1 vccd1 _08226_ sky130_fd_sc_hd__or2_1
X_16090_ _09125_ _09147_ _09148_ _09164_ _09146_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_181_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15041_ _08031_ _08141_ net7478 vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__mux2_1
X_12253_ net2942 _05378_ _05379_ net2940 vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11204_ net2174 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20825__247 clknet_1_1__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__inv_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ _05329_ net4073 vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__xnor2_2
X_18800_ _02791_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__or2_1
X_11135_ _04403_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__buf_4
X_19780_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__buf_4
X_16992_ _10003_ net4507 _09966_ vssd1 vssd1 vccd1 vccd1 _10004_ sky130_fd_sc_hd__mux2_1
X_18731_ _06205_ _06189_ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__or3_1
X_11066_ net6678 net2424 _04404_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_1
X_15943_ _09000_ _09001_ _08999_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__a21o_1
X_18662_ _02654_ _02667_ _02669_ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _08907_ _08912_ _08926_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__nand3_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _01662_ _01663_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__and2_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _07975_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__inv_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18593_ net4667 net7601 _02603_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__and3_1
Xclkbuf_0__04001_ _04001_ vssd1 vssd1 vccd1 vccd1 clknet_0__04001_ sky130_fd_sc_hd__clkbuf_16
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _10541_ _10542_ vssd1 vssd1 vccd1 vccd1 _10543_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _07905_ _07906_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__and2_1
X_20719__152 clknet_1_1__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__inv_2
X_11968_ net2993 _05125_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__xnor2_1
X_13707_ _06737_ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__xnor2_4
X_10919_ net5844 net5931 _04333_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17475_ _09562_ _09420_ vssd1 vssd1 vccd1 vccd1 _10474_ sky130_fd_sc_hd__nor2_1
X_11899_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14687_ _07811_ _07836_ _07837_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__a21oi_2
X_19214_ net5428 _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__or2_1
X_16426_ _09493_ _09494_ _09365_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13638_ _06662_ _06784_ _06787_ _06788_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19145_ _03036_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__clkbuf_4
X_16357_ _08310_ _09311_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ _06717_ _06719_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6109 _04290_ vssd1 vssd1 vccd1 vccd1 net6633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15308_ net4338 _08362_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ net4318 net2842 net643 _03022_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__o211a_1
Xhold5408 _04335_ vssd1 vssd1 vccd1 vccd1 net5932 sky130_fd_sc_hd__dlygate4sd3_1
X_16288_ _09358_ _09361_ vssd1 vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__xor2_2
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5419 rbzero.map_overlay.i_otherx\[1\] vssd1 vssd1 vccd1 vccd1 net5943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18027_ _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nand2_1
X_15239_ _08299_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4707 _00713_ vssd1 vssd1 vccd1 vccd1 net5231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4718 rbzero.spi_registers.buf_mapdyw\[0\] vssd1 vssd1 vccd1 vccd1 net5242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4729 net1233 vssd1 vssd1 vccd1 vccd1 net5253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19978_ net951 _03578_ net4443 _03550_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18929_ _02864_ net3700 _05391_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__or3b_2
XFILLER_0_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21940_ clknet_leaf_9_i_clk net4863 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21871_ clknet_leaf_100_i_clk net1244 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20930__342 clknet_1_1__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__inv_2
XFILLER_0_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7300 _10086_ vssd1 vssd1 vccd1 vccd1 net7824 sky130_fd_sc_hd__dlygate4sd3_1
X_22423_ clknet_leaf_55_i_clk net5336 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
Xhold7322 rbzero.row_render.size\[0\] vssd1 vssd1 vccd1 vccd1 net7846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6610 rbzero.tex_b0\[49\] vssd1 vssd1 vccd1 vccd1 net7134 sky130_fd_sc_hd__dlygate4sd3_1
X_22354_ net486 net1455 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold6621 net2325 vssd1 vssd1 vccd1 vccd1 net7145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6632 rbzero.tex_g1\[55\] vssd1 vssd1 vccd1 vccd1 net7156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7377 net4375 vssd1 vssd1 vccd1 vccd1 net7901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6643 net2625 vssd1 vssd1 vccd1 vccd1 net7167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7388 _06722_ vssd1 vssd1 vccd1 vccd1 net7912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6654 rbzero.tex_b0\[44\] vssd1 vssd1 vccd1 vccd1 net7178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7399 _08301_ vssd1 vssd1 vccd1 vccd1 net7923 sky130_fd_sc_hd__dlygate4sd3_1
X_21305_ clknet_leaf_74_i_clk net3990 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold6665 net2785 vssd1 vssd1 vccd1 vccd1 net7189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5920 rbzero.tex_r1\[10\] vssd1 vssd1 vccd1 vccd1 net6444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6676 rbzero.tex_b1\[31\] vssd1 vssd1 vccd1 vccd1 net7200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5931 net1454 vssd1 vssd1 vccd1 vccd1 net6455 sky130_fd_sc_hd__dlygate4sd3_1
X_22285_ net417 net2783 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold5942 _04267_ vssd1 vssd1 vccd1 vccd1 net6466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6687 net2656 vssd1 vssd1 vccd1 vccd1 net7211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6698 rbzero.tex_b0\[32\] vssd1 vssd1 vccd1 vccd1 net7222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5953 net1417 vssd1 vssd1 vccd1 vccd1 net6477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5964 rbzero.tex_r0\[49\] vssd1 vssd1 vccd1 vccd1 net6488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 net7517 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
X_21236_ clknet_leaf_59_i_clk _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5975 rbzero.tex_r0\[19\] vssd1 vssd1 vccd1 vccd1 net6499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 net7472 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5986 net1443 vssd1 vssd1 vccd1 vccd1 net6510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5997 _04223_ vssd1 vssd1 vccd1 vccd1 net6521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 net4325 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 net5064 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 net5100 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
X_21167_ net4111 _09941_ _09942_ _09284_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__a22o_1
X_20118_ net3561 net4837 net2122 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__or3b_1
X_21098_ _04087_ net4937 _04089_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20049_ net3323 _03613_ net4464 _03602_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__o211a_1
X_12940_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__and2_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _06026_ _06028_ net31 vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__mux2_1
XANTENNA_101 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _07644_ _07646_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__or2_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__buf_4
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _08311_ net4954 vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__nor2_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ net757 net2194 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14541_ _07690_ _07691_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__and2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ net7197 net7280 _04214_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _10258_ _10260_ vssd1 vssd1 vccd1 vccd1 _10261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14472_ _06922_ _07466_ _06923_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__and3b_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _04726_ net4891 net3868 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16211_ _09174_ _09177_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__xor2_4
XFILLER_0_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ net6910 net7181 _04181_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__mux2_1
X_13423_ net6146 _06431_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ _09895_ _09896_ vssd1 vssd1 vccd1 vccd1 _10193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _08559_ _08560_ _08581_ _09216_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13354_ net7582 _06156_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_91_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12305_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _05230_ vssd1 vssd1 vccd1 vccd1 _05473_
+ sky130_fd_sc_hd__mux2_1
X_16073_ _09140_ _09145_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13285_ net4561 net7146 vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__nand2_1
X_15024_ net4378 _08160_ _08138_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__mux2_1
X_12236_ _05403_ _05377_ _05379_ rbzero.debug_overlay.vplaneX\[-7\] _05404_ vssd1
+ vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a221o_1
X_19901_ net6140 _03521_ net3157 _03474_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19832_ net5467 _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and2_1
X_12167_ _05329_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__inv_2
X_11118_ net6672 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
X_19763_ net1608 _03427_ net1904 _03424_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__o211a_1
X_12098_ rbzero.tex_r1\[1\] rbzero.tex_r1\[0\] _05072_ vssd1 vssd1 vccd1 vccd1 _05267_
+ sky130_fd_sc_hd__mux2_1
X_16975_ net4568 net4566 vssd1 vssd1 vccd1 vccd1 _09988_ sky130_fd_sc_hd__nand2_1
X_18714_ _02716_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__nand2_1
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net6620 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
X_15926_ _08347_ _08367_ _08432_ _08455_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19694_ net6047 _03359_ net1671 _03384_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__o211a_1
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
XFILLER_0_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18645_ _02630_ _02634_ _02652_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08909_ _08931_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__nor2_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _07913_ _07914_ _07905_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_204_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18576_ _02579_ _02584_ net4692 net3406 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__a31o_1
X_15788_ _08840_ _08843_ _08862_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__a21bo_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _10507_ _10508_ _10525_ vssd1 vssd1 vccd1 vccd1 _10526_ sky130_fd_sc_hd__a21o_1
X_14739_ _07444_ _07805_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ _10457_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16409_ net3537 _08313_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17389_ _08717_ _09216_ vssd1 vssd1 vccd1 vccd1 _10389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19128_ net5190 _03053_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5205 _03396_ vssd1 vssd1 vccd1 vccd1 net5729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5216 net1827 vssd1 vssd1 vccd1 vccd1 net5740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19059_ net3038 net2843 _03013_ _03011_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__o211a_1
Xhold5227 _00763_ vssd1 vssd1 vccd1 vccd1 net5751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5238 net1115 vssd1 vssd1 vccd1 vccd1 net5762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4504 net766 vssd1 vssd1 vccd1 vccd1 net5028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5249 net1650 vssd1 vssd1 vccd1 vccd1 net5773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4515 _00876_ vssd1 vssd1 vccd1 vccd1 net5039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4526 _01068_ vssd1 vssd1 vccd1 vccd1 net5050 sky130_fd_sc_hd__dlygate4sd3_1
X_22070_ clknet_leaf_13_i_clk net3815 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4537 net758 vssd1 vssd1 vccd1 vccd1 net5061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4548 net769 vssd1 vssd1 vccd1 vccd1 net5072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3803 _03357_ vssd1 vssd1 vccd1 vccd1 net4327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3814 net7731 vssd1 vssd1 vccd1 vccd1 net4338 sky130_fd_sc_hd__clkbuf_2
X_21021_ net1011 net5271 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4559 net878 vssd1 vssd1 vccd1 vccd1 net5083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3825 net3046 vssd1 vssd1 vccd1 vccd1 net4349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3836 net2916 vssd1 vssd1 vccd1 vccd1 net4360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3847 net7488 vssd1 vssd1 vccd1 vccd1 net4371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3858 net3138 vssd1 vssd1 vccd1 vccd1 net4382 sky130_fd_sc_hd__buf_1
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3869 net3148 vssd1 vssd1 vccd1 vccd1 net4393 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21923_ clknet_leaf_6_i_clk net1323 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ clknet_leaf_82_i_clk net3810 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21785_ clknet_leaf_93_i_clk net626 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7130 rbzero.spi_registers.texadd2\[16\] vssd1 vssd1 vccd1 vccd1 net7654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22406_ net158 net2365 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
Xhold7141 rbzero.spi_registers.buf_texadd3\[8\] vssd1 vssd1 vccd1 vccd1 net7665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7152 rbzero.traced_texa\[-11\] vssd1 vssd1 vccd1 vccd1 net7676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20598_ net3252 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_1
Xhold6440 net1813 vssd1 vssd1 vccd1 vccd1 net6964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6451 rbzero.tex_b0\[47\] vssd1 vssd1 vccd1 vccd1 net6975 sky130_fd_sc_hd__dlygate4sd3_1
X_22337_ net469 net2501 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6462 net2004 vssd1 vssd1 vccd1 vccd1 net6986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6473 rbzero.tex_g0\[59\] vssd1 vssd1 vccd1 vccd1 net6997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6484 net2406 vssd1 vssd1 vccd1 vccd1 net7008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6495 rbzero.tex_b1\[5\] vssd1 vssd1 vccd1 vccd1 net7019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5750 rbzero.spi_registers.buf_leak\[2\] vssd1 vssd1 vccd1 vccd1 net6274 sky130_fd_sc_hd__dlygate4sd3_1
X_13070_ net3853 vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__inv_2
X_22268_ net400 net2211 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
Xhold5761 net1912 vssd1 vssd1 vccd1 vccd1 net6285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5772 _00818_ vssd1 vssd1 vccd1 vccd1 net6296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5783 net1467 vssd1 vssd1 vccd1 vccd1 net6307 sky130_fd_sc_hd__dlygate4sd3_1
X_12021_ _04627_ _04817_ _04820_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__o22a_1
Xhold5794 net634 vssd1 vssd1 vccd1 vccd1 net6318 sky130_fd_sc_hd__dlygate4sd3_1
X_21219_ clknet_leaf_43_i_clk net4889 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22199_ net331 net2872 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16760_ _09700_ _09709_ _09707_ vssd1 vssd1 vccd1 vccd1 _09830_ sky130_fd_sc_hd__a21o_1
X_13972_ _06885_ _06922_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nor2_1
X_15711_ _08749_ _08776_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__nor2_1
X_12923_ _04760_ _04603_ _04637_ _04165_ net34 net35 vssd1 vssd1 vccd1 vccd1 _06080_
+ sky130_fd_sc_hd__mux4_1
X_16691_ _09691_ _09761_ vssd1 vssd1 vccd1 vccd1 _09762_ sky130_fd_sc_hd__xnor2_4
X_20937__348 clknet_1_1__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__inv_2
XFILLER_0_88_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18430_ _02456_ _02457_ _01971_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__o21ai_1
X_15642_ _08498_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__buf_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ net29 net28 vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__and2_2
XFILLER_0_186_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11805_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__clkbuf_8
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _02397_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__clkbuf_1
X_15573_ _08636_ _08640_ _08647_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__nand3_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ net26 net27 vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__nor2_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17312_ _10310_ _10312_ vssd1 vssd1 vccd1 vccd1 _10313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _07232_ _06918_ _07463_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__or3_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _04803_ net2987 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and2_1
X_18292_ _06204_ _08314_ _06388_ net4919 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _10235_ _10243_ vssd1 vssd1 vccd1 vccd1 _10244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03981_ _03981_ vssd1 vssd1 vccd1 vccd1 clknet_0__03981_ sky130_fd_sc_hd__clkbuf_16
X_14455_ _07367_ _07399_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__or2_1
X_11667_ net3821 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13406_ _06544_ _06552_ _06554_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__or4_4
X_17174_ _09871_ _09874_ _09872_ vssd1 vssd1 vccd1 vccd1 _10176_ sky130_fd_sc_hd__a21bo_1
X_10618_ net2427 net6516 _04170_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14386_ net587 net3333 _07467_ _07536_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__a31o_1
X_11598_ rbzero.spi_registers.texadd1\[0\] _04644_ _04709_ vssd1 vssd1 vccd1 vccd1
+ _04770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16125_ _09197_ _09198_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _06447_ _06487_ _06446_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20682__118 clknet_1_0__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__inv_2
X_16056_ _08490_ _08755_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13268_ rbzero.wall_tracer.rcp_sel\[0\] _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15007_ _08132_ _07993_ _07991_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__mux2_1
X_12219_ net3857 _05372_ _05375_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a211o_1
X_13199_ net2839 _06229_ _06244_ net2905 vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__a22o_1
Xhold2409 net5462 vssd1 vssd1 vccd1 vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
X_19815_ _02967_ net3152 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__and2_1
Xhold1708 net6039 vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 net2448 vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_19746_ net1537 _03394_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__or2_1
X_16958_ _09948_ _09957_ vssd1 vssd1 vccd1 vccd1 _09974_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15909_ _08872_ _08517_ _08874_ _08873_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__o22ai_1
X_19677_ net3070 _03374_ net2594 _03371_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__o211a_1
X_16889_ _09935_ vssd1 vssd1 vccd1 vccd1 _09938_ sky130_fd_sc_hd__buf_4
XFILLER_0_177_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18628_ _02637_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02638_
+ sky130_fd_sc_hd__nand2_1
X_18559_ net3241 rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1 vccd1 _02574_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21570_ clknet_leaf_17_i_clk net4985 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ net3580 net1493 _03889_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__mux2_1
XANTENNA_23 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _09286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 rbzero.wall_tracer.visualWallDist\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 net6146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_67 _10454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20452_ net3559 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_89 _05995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5002 rbzero.spi_registers.texadd2\[18\] vssd1 vssd1 vccd1 vccd1 net5526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20383_ _03791_ net3429 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__and2_1
Xhold5013 _00784_ vssd1 vssd1 vccd1 vccd1 net5537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5024 _00832_ vssd1 vssd1 vccd1 vccd1 net5548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5035 net1185 vssd1 vssd1 vccd1 vccd1 net5559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22122_ net254 net2184 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold4301 _00386_ vssd1 vssd1 vccd1 vccd1 net4825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5046 rbzero.pov.spi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net5570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5057 rbzero.pov.spi_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net5581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4312 rbzero.pov.sclk_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net4836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4323 rbzero.pov.spi_buffer\[64\] vssd1 vssd1 vccd1 vccd1 net4847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5068 _01056_ vssd1 vssd1 vccd1 vccd1 net5592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5079 _01057_ vssd1 vssd1 vccd1 vccd1 net5603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4334 rbzero.pov.spi_buffer\[68\] vssd1 vssd1 vccd1 vccd1 net4858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4345 _01108_ vssd1 vssd1 vccd1 vccd1 net4869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3600 net7628 vssd1 vssd1 vccd1 vccd1 net4124 sky130_fd_sc_hd__dlygate4sd3_1
X_20988__15 clknet_1_1__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
Xhold3611 net683 vssd1 vssd1 vccd1 vccd1 net4135 sky130_fd_sc_hd__dlygate4sd3_1
X_22053_ clknet_leaf_90_i_clk net3614 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4356 rbzero.pov.spi_buffer\[71\] vssd1 vssd1 vccd1 vccd1 net4880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4367 net2986 vssd1 vssd1 vccd1 vccd1 net4891 sky130_fd_sc_hd__clkbuf_4
Xhold3622 net7635 vssd1 vssd1 vccd1 vccd1 net4146 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3633 net689 vssd1 vssd1 vccd1 vccd1 net4157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4378 _09964_ vssd1 vssd1 vccd1 vccd1 net4902 sky130_fd_sc_hd__clkbuf_4
Xhold3644 _00510_ vssd1 vssd1 vccd1 vccd1 net4168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4389 _06245_ vssd1 vssd1 vccd1 vccd1 net4913 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3655 rbzero.traced_texa\[1\] vssd1 vssd1 vccd1 vccd1 net4179 sky130_fd_sc_hd__buf_1
Xhold2910 net5693 vssd1 vssd1 vccd1 vccd1 net3434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3666 net1072 vssd1 vssd1 vccd1 vccd1 net4190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2921 _02889_ vssd1 vssd1 vccd1 vccd1 net3445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3677 net1257 vssd1 vssd1 vccd1 vccd1 net4201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2932 _01190_ vssd1 vssd1 vccd1 vccd1 net3456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2943 _03812_ vssd1 vssd1 vccd1 vccd1 net3467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3688 _00760_ vssd1 vssd1 vccd1 vccd1 net4212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2954 _03917_ vssd1 vssd1 vccd1 vccd1 net3478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3699 net4214 vssd1 vssd1 vccd1 vccd1 net4223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2965 _03914_ vssd1 vssd1 vccd1 vccd1 net3489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2976 net4559 vssd1 vssd1 vccd1 vccd1 net3500 sky130_fd_sc_hd__buf_1
XFILLER_0_173_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2987 _08292_ vssd1 vssd1 vccd1 vccd1 net3511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2998 _01212_ vssd1 vssd1 vccd1 vccd1 net3522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21906_ clknet_leaf_93_i_clk net1414 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21837_ clknet_leaf_83_i_clk net3879 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12570_ _05051_ _05709_ _05717_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21768_ clknet_leaf_8_i_clk net1991 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ net6497 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21699_ clknet_leaf_5_i_clk net743 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14240_ _07337_ _07363_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a21oi_4
X_11452_ net4026 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_151_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14171_ _07310_ _07321_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11383_ net6970 net6952 _04573_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6270 net1795 vssd1 vssd1 vccd1 vccd1 net6794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6281 rbzero.tex_b0\[24\] vssd1 vssd1 vccd1 vccd1 net6805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ net3462 _06276_ net3500 _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__o22a_1
Xhold6292 net2434 vssd1 vssd1 vccd1 vccd1 net6816 sky130_fd_sc_hd__dlygate4sd3_1
X_20294__31 clknet_1_1__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5580 net642 vssd1 vssd1 vccd1 vccd1 net6104 sky130_fd_sc_hd__dlymetal6s2s_1
X_13053_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__buf_6
X_17930_ _01976_ _01977_ _01870_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12004_ net2869 _05154_ _05156_ _05172_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a221o_1
X_17861_ _01825_ _01830_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__nand2_1
Xhold4890 _00796_ vssd1 vssd1 vccd1 vccd1 net5414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16812_ _09879_ _09880_ _09868_ vssd1 vssd1 vccd1 vccd1 _09882_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19600_ net5197 _03325_ _03335_ _03330_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__o211a_1
X_17792_ _01841_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19531_ _02998_ _03289_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or2_1
X_16743_ _08372_ _08795_ vssd1 vssd1 vccd1 vccd1 _09813_ sky130_fd_sc_hd__or2_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13955_ _07081_ _07105_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_199_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19462_ _02492_ _02498_ _03238_ net1790 vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a31o_1
X_12906_ net36 net39 _06049_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__and4b_1
XFILLER_0_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16674_ _08613_ _09744_ _09611_ _09612_ _09604_ vssd1 vssd1 vccd1 vccd1 _09745_ sky130_fd_sc_hd__a32o_1
X_13886_ _07032_ net570 _07036_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__a21bo_4
X_18413_ _10010_ _02442_ _01747_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o21ai_1
X_15625_ _08310_ _08331_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _05995_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
X_19393_ net1903 _03199_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18344_ _02382_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ net3539 _08304_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__nor2_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _04159_ net4891 _04726_ _04777_ net16 net17 vssd1 vssd1 vccd1 vccd1 _05928_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _07652_ _07655_ _07656_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__nand3_1
X_18275_ _02315_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__xnor2_1
X_11719_ net4013 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__clkinv_4
X_15487_ _08558_ _08561_ _08551_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_86_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12699_ net13 _05857_ _05859_ net12 vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a31o_1
X_17226_ _08724_ _09666_ vssd1 vssd1 vccd1 vccd1 _10227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_4
X_14438_ _07305_ _07588_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
Xinput32 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_2
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput43 i_reg_csb vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_4
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_8
X_17157_ _10157_ _10158_ vssd1 vssd1 vccd1 vccd1 _10159_ sky130_fd_sc_hd__xnor2_2
Xhold805 net5557 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _07488_ _07519_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__xor2_1
Xhold816 net5569 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16108_ _08836_ _09182_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__xnor2_4
Xhold827 net5670 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 net3597 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _09826_ _10088_ _10089_ vssd1 vssd1 vccd1 vccd1 _10090_ sky130_fd_sc_hd__a21oi_2
Xhold849 net6426 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16039_ _09082_ _09112_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2206 _01537_ vssd1 vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2217 _04434_ vssd1 vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2228 _01577_ vssd1 vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2239 net7230 vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1505 _01142_ vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 net7068 vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 net6955 vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 _01488_ vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 net6745 vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19729_ net5795 _03408_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__or2_1
XFILLER_0_212_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21622_ clknet_leaf_4_i_clk net5580 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ clknet_leaf_5_i_clk net1051 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20504_ _08274_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__buf_2
XFILLER_0_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21484_ clknet_leaf_93_i_clk net623 vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20435_ _03814_ net3757 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20366_ net1623 net3641 _03782_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22105_ net237 net2607 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold4131 net1505 vssd1 vssd1 vccd1 vccd1 net4655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4142 rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 net4666 sky130_fd_sc_hd__buf_2
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4153 net641 vssd1 vssd1 vccd1 vccd1 net4677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4164 net7562 vssd1 vssd1 vccd1 vccd1 net4688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4175 net3690 vssd1 vssd1 vccd1 vccd1 net4699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3430 _03576_ vssd1 vssd1 vccd1 vccd1 net3954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4186 _02821_ vssd1 vssd1 vccd1 vccd1 net4710 sky130_fd_sc_hd__dlygate4sd3_1
X_22036_ clknet_leaf_95_i_clk net3785 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3441 _05824_ vssd1 vssd1 vccd1 vccd1 net3965 sky130_fd_sc_hd__clkbuf_4
Xhold4197 _02855_ vssd1 vssd1 vccd1 vccd1 net4721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3452 _09914_ vssd1 vssd1 vccd1 vccd1 net3976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3463 net6048 vssd1 vssd1 vccd1 vccd1 net3987 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3474 _02949_ vssd1 vssd1 vccd1 vccd1 net3998 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3485 net7364 vssd1 vssd1 vccd1 vccd1 net4009 sky130_fd_sc_hd__clkbuf_4
Xhold2740 _00419_ vssd1 vssd1 vccd1 vccd1 net3264 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2751 net1239 vssd1 vssd1 vccd1 vccd1 net3275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3496 net7307 vssd1 vssd1 vccd1 vccd1 net4020 sky130_fd_sc_hd__clkbuf_2
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2762 net639 vssd1 vssd1 vccd1 vccd1 net3286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2773 _03834_ vssd1 vssd1 vccd1 vccd1 net3297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2784 _01216_ vssd1 vssd1 vccd1 vccd1 net3308 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2795 _03805_ vssd1 vssd1 vccd1 vccd1 net3319 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13740_ _06889_ _06887_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__nand3_2
X_10952_ net6582 net2234 _04344_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _06820_ _06821_ _06788_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__o21ai_1
X_10883_ net2748 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__clkbuf_1
X_15410_ _08456_ _08484_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12622_ net9 net8 vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nor2_1
X_16390_ _09443_ _09462_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15341_ net645 _08415_ _08303_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _05541_ vssd1 vssd1 vccd1 vccd1 _05718_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18060_ _02093_ _02107_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__xnor2_1
X_11504_ _04646_ _04647_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__nor2_1
X_15272_ _08346_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__buf_2
X_12484_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _05218_ vssd1 vssd1 vccd1 vccd1 _05650_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17011_ _10010_ _09284_ vssd1 vssd1 vccd1 vccd1 _10021_ sky130_fd_sc_hd__nand2_1
X_14223_ _07281_ _07330_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _04601_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ net6508 net2804 _04562_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__mux2_1
X_14154_ _07303_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13105_ net2802 net4897 _06244_ net2879 _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11297_ net5953 net5817 _04529_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
X_14085_ _07207_ _07235_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__or2_1
X_18962_ _04624_ _02941_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a21o_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nor2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ net6186 _06189_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o21a_1
X_18893_ net4662 net7598 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__and2_1
XFILLER_0_206_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _01892_ _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20794__219 clknet_1_1__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__inv_2
X_17775_ _09108_ _01711_ _10539_ _10406_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__o22ai_1
X_14987_ _08070_ _08093_ _08111_ _08128_ _08069_ net7759 vssd1 vssd1 vccd1 vccd1 _08129_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_117_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16726_ _09091_ _09312_ _09419_ _08724_ vssd1 vssd1 vccd1 vccd1 _09796_ sky130_fd_sc_hd__o22a_1
X_19514_ net1608 _03275_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13938_ _06826_ _06922_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19445_ _02507_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16657_ _09139_ _09484_ _09603_ _09138_ vssd1 vssd1 vccd1 vccd1 _09728_ sky130_fd_sc_hd__o22ai_1
X_13869_ _07013_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__xnor2_1
X_15608_ _08681_ _08682_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19376_ net1644 _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__or2_1
X_16588_ _09580_ _09560_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__or2b_1
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18327_ _02367_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15539_ _08604_ _08591_ _08605_ _08534_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18258_ _01778_ _09418_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nor2_1
X_20688__124 clknet_1_1__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__inv_2
XFILLER_0_142_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ net4540 net4411 vssd1 vssd1 vccd1 vccd1 _10210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18189_ _02204_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold602 net5475 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20220_ net1284 _03731_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__or2_1
Xhold613 _01649_ vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 net6394 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold635 net6402 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03778_ clknet_0__03778_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03778_
+ sky130_fd_sc_hd__clkbuf_16
Xhold646 net3589 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _01552_ vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold668 net6450 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20151_ net3660 _03692_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__or2_1
Xhold679 _01412_ vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2003 net7031 vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
X_20082_ net4634 _03581_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__or2_1
Xhold2014 net7142 vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _01404_ vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2036 _04295_ vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _01150_ vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2047 net7160 vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1313 _01583_ vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2058 _04556_ vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 net6927 vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 _03452_ vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1335 net7664 vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1346 _00904_ vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 _04508_ vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1368 net6627 vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1379 net6623 vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21605_ clknet_leaf_1_i_clk net5525 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21536_ clknet_leaf_36_i_clk net1916 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21467_ clknet_leaf_24_i_clk net3094 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11220_ net2508 net6493 _04492_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20418_ net3323 net1276 _03801_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__mux2_1
X_21398_ clknet_leaf_64_i_clk _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11151_ net5937 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11082_ net5836 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
Xhold3260 _03851_ vssd1 vssd1 vccd1 vccd1 net3784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3271 net3200 vssd1 vssd1 vccd1 vccd1 net3795 sky130_fd_sc_hd__dlymetal6s2s_1
X_22019_ clknet_leaf_99_i_clk net3469 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14910_ net7433 _08052_ _08058_ _08047_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__a31o_1
XFILLER_0_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3282 _00595_ vssd1 vssd1 vccd1 vccd1 net3806 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15890_ _08957_ _08964_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__xnor2_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3293 net1328 vssd1 vssd1 vccd1 vccd1 net3817 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2570 _00636_ vssd1 vssd1 vccd1 vccd1 net3094 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2581 _03248_ vssd1 vssd1 vccd1 vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
X_14841_ _07584_ _07978_ _07581_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__o21ai_2
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2592 rbzero.spi_registers.buf_floor\[5\] vssd1 vssd1 vccd1 vccd1 net3116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _10433_ _10435_ vssd1 vssd1 vccd1 vccd1 _10559_ sky130_fd_sc_hd__nor2_1
Xhold1880 _01360_ vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1891 net7086 vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_14772_ _07894_ _07896_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__xnor2_1
X_11984_ net3040 net2955 net2069 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16511_ _09582_ _08588_ _09469_ _09468_ _09467_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__o32a_1
XFILLER_0_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13723_ _06870_ _06871_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__nand2_1
X_10935_ net6367 net7227 _04333_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__mux2_1
X_17491_ _10130_ _09312_ _10488_ vssd1 vssd1 vccd1 vccd1 _10490_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19230_ net5669 _03106_ _03116_ _03115_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__o211a_1
X_16442_ _09513_ _09514_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _06803_ _06804_ _06765_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__o21a_1
X_10866_ net7117 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12605_ _05735_ _05769_ _04975_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__mux2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ net5678 _03065_ _03073_ _03074_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16373_ _09187_ _09328_ _08962_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__or3b_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _06711_ _06735_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__nor2_4
X_10797_ net6706 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _02157_ _02159_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15324_ _08398_ net4294 _06177_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__mux2_1
X_19092_ _09929_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nor2_2
X_12536_ net947 net3128 _05120_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18043_ _01825_ _02022_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ _08328_ net7477 vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__or2_1
X_12467_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _05072_ vssd1 vssd1 vccd1 vccd1 _05633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ _07301_ _07306_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11418_ net5767 net1521 _04243_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15186_ net4605 _08186_ _08260_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__mux2_1
X_12398_ _04993_ _05562_ _05564_ _05009_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _07008_ _07261_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__o21ai_2
X_11349_ net6838 net2027 _04551_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__mux2_1
X_19994_ _03261_ net3787 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ _07216_ _07209_ _07214_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nor3_1
X_18945_ _02913_ _02917_ _02927_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_197_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ _06152_ _06169_ _06171_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18876_ _02854_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17827_ _01776_ _01793_ _01791_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17758_ _10520_ _09861_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16709_ _09768_ vssd1 vssd1 vccd1 vccd1 _09779_ sky130_fd_sc_hd__inv_2
X_17689_ _01739_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19428_ net1566 _03225_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19359_ net4257 _03186_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22370_ net502 net2704 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6803 net7365 vssd1 vssd1 vccd1 vccd1 net7327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6814 rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 net7338 sky130_fd_sc_hd__dlygate4sd3_1
X_21321_ clknet_leaf_72_i_clk _00490_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6825 _03587_ vssd1 vssd1 vccd1 vccd1 net7349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6836 rbzero.spi_registers.spi_cmd\[3\] vssd1 vssd1 vccd1 vccd1 net7360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6847 _09287_ vssd1 vssd1 vccd1 vccd1 net7371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 _01442_ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21252_ clknet_leaf_52_i_clk net3202 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold421 net5378 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 net5297 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
X_20203_ net3412 _03718_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or2_1
Xhold443 net5343 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 net5421 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21183_ net4424 net701 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__or2_1
Xhold465 net5262 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 net5405 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 rbzero.traced_texa\[-9\] vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkdlybuf4s25_1
X_20134_ net1204 _03679_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__or2_1
Xhold498 net5403 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20065_ net719 _03577_ net4641 _03636_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__o211a_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20742__173 clknet_1_0__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__inv_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 net5782 vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _03417_ vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _03192_ vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 net6607 vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 net6705 vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 net7665 vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 net4671 vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _00927_ vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 net5789 vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10720_ net2260 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10651_ _04169_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ _06520_ _06475_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _05482_ _05485_ _05488_ _05061_ _05023_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21519_ clknet_leaf_35_i_clk net3147 vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15040_ _08174_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12252_ net3024 _05377_ _05382_ rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1
+ vccd1 _05421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11203_ net2173 net7225 _04481_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12183_ net4038 net4072 _05337_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11134_ net6658 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
X_16991_ _06206_ _09998_ _10002_ vssd1 vssd1 vccd1 vccd1 _10003_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_82_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11065_ net6451 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
X_15942_ _08999_ _09000_ _09001_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__nand3_1
X_18730_ _06185_ _06188_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__nor2_1
Xhold3090 _01222_ vssd1 vssd1 vccd1 vccd1 net3614 sky130_fd_sc_hd__dlygate4sd3_1
X_18661_ _02650_ _02668_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _08929_ _08930_ _08932_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__a21o_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _01662_ _01663_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nor2_1
X_14824_ _07972_ _07974_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ net4667 _02602_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_97_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04000_ _04000_ vssd1 vssd1 vccd1 vccd1 clknet_0__04000_ sky130_fd_sc_hd__clkbuf_16
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17543_ _09138_ _09139_ _10168_ vssd1 vssd1 vccd1 vccd1 _10542_ sky130_fd_sc_hd__a21oi_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _07367_ _07805_ _07904_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__o21ai_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _05126_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13706_ _06846_ net79 vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__nor2_8
X_10918_ net933 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__clkbuf_1
X_17474_ _10401_ _10376_ vssd1 vssd1 vccd1 vccd1 _10473_ sky130_fd_sc_hd__or2b_1
X_14686_ _07812_ _07835_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_20_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11898_ _04982_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__buf_4
X_16425_ _09481_ _09497_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__xnor2_2
X_19213_ _03039_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13637_ _06762_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__clkbuf_2
X_10849_ net2011 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19144_ net5978 _03052_ _03064_ _03061_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__o211a_1
X_16356_ _09427_ _09428_ vssd1 vssd1 vccd1 vccd1 _09429_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13568_ _06608_ _06688_ _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15307_ net4338 _08381_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__nand2_1
X_12519_ _05683_ _05684_ _05068_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__mux2_1
X_19075_ _02992_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__buf_4
X_16287_ _09359_ _09360_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_35_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ _06565_ _06587_ _06632_ _06629_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__and4_1
Xhold5409 net1942 vssd1 vssd1 vccd1 vccd1 net5933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18026_ net4497 net4619 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__nand2_1
X_15238_ _08312_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4708 rbzero.pov.spi_buffer\[33\] vssd1 vssd1 vccd1 vccd1 net5232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4719 net843 vssd1 vssd1 vccd1 vccd1 net5243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15169_ net4411 _08152_ _08260_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19977_ rbzero.debug_overlay.facingX\[-7\] _03582_ vssd1 vssd1 vccd1 vccd1 _03585_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18928_ _02910_ _02911_ _02895_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18859_ net3700 net4799 _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21870_ clknet_leaf_100_i_clk net1329 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20772__199 clknet_1_1__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__inv_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7301 rbzero.wall_tracer.stepDistY\[-8\] vssd1 vssd1 vccd1 vccd1 net7825 sky130_fd_sc_hd__dlygate4sd3_1
X_22422_ clknet_leaf_55_i_clk net5273 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7312 _06716_ vssd1 vssd1 vccd1 vccd1 net7836 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6600 rbzero.tex_b0\[22\] vssd1 vssd1 vccd1 vccd1 net7124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6611 net2346 vssd1 vssd1 vccd1 vccd1 net7135 sky130_fd_sc_hd__dlygate4sd3_1
X_22353_ net485 net2369 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
Xhold7356 rbzero.texu_hot\[1\] vssd1 vssd1 vccd1 vccd1 net7880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6622 net3194 vssd1 vssd1 vccd1 vccd1 net7146 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold7367 _06838_ vssd1 vssd1 vccd1 vccd1 net7891 sky130_fd_sc_hd__clkbuf_2
Xhold6633 net2452 vssd1 vssd1 vccd1 vccd1 net7157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7378 rbzero.wall_tracer.stepDistX\[9\] vssd1 vssd1 vccd1 vccd1 net7902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6644 rbzero.tex_r1\[15\] vssd1 vssd1 vccd1 vccd1 net7168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6655 net2316 vssd1 vssd1 vccd1 vccd1 net7179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5910 _04356_ vssd1 vssd1 vccd1 vccd1 net6434 sky130_fd_sc_hd__dlygate4sd3_1
X_21304_ clknet_leaf_12_i_clk net3871 vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_1
X_22284_ net416 net2627 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
Xhold5921 net1347 vssd1 vssd1 vccd1 vccd1 net6445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6666 rbzero.tex_r0\[46\] vssd1 vssd1 vccd1 vccd1 net7190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5932 rbzero.tex_g0\[28\] vssd1 vssd1 vccd1 vccd1 net6456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6677 net2508 vssd1 vssd1 vccd1 vccd1 net7201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6688 rbzero.tex_g1\[37\] vssd1 vssd1 vccd1 vccd1 net7212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5943 net1353 vssd1 vssd1 vccd1 vccd1 net6467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6699 net2619 vssd1 vssd1 vccd1 vccd1 net7223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5954 _04565_ vssd1 vssd1 vccd1 vccd1 net6478 sky130_fd_sc_hd__dlygate4sd3_1
X_21235_ clknet_leaf_59_i_clk _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5965 net1424 vssd1 vssd1 vccd1 vccd1 net6489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 net5008 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5976 net1477 vssd1 vssd1 vccd1 vccd1 net6500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 net4978 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5987 rbzero.tex_g1\[24\] vssd1 vssd1 vccd1 vccd1 net6511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 net5044 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _03323_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5998 net1449 vssd1 vssd1 vccd1 vccd1 net6522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 net5066 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21166_ net4962 net65 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nor2_1
Xhold295 net5075 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20117_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__buf_2
X_21097_ _04082_ _04086_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nand2_1
X_20048_ net4463 _03614_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ net3937 _06012_ _06008_ net3930 _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a221o_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _04953_ _04971_ _04980_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__nor3_4
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ net224 net1972 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _07585_ _07637_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__xor2_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _04920_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ net6361 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14471_ _07598_ _07621_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__xnor2_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _04164_ _04790_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or3b_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16210_ net3024 net4306 net4087 vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13422_ _06559_ _06562_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and2b_1
X_17190_ _10125_ _10191_ vssd1 vssd1 vccd1 vccd1 _10192_ sky130_fd_sc_hd__xnor2_1
X_10634_ net7155 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ _08596_ _08597_ _08598_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_107_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13353_ net3356 _06430_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12304_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _05263_ vssd1 vssd1 vccd1 vccd1 _05472_
+ sky130_fd_sc_hd__mux2_1
X_16072_ _09127_ _09144_ _09146_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ net4561 net7146 vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__or2_2
X_20749__179 clknet_1_0__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__inv_2
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19900_ net3156 _03471_ _03520_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__a22o_1
X_15023_ _08150_ _08104_ _08159_ net6162 vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__a211o_2
X_12235_ rbzero.debug_overlay.vplaneX\[-9\] _05382_ _05378_ rbzero.debug_overlay.vplaneX\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19831_ _03034_ _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__nand2_2
X_12166_ _05326_ _05329_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or3_1
X_11117_ net6670 net1935 _04437_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__mux2_1
X_19762_ net6624 _03429_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__or2_1
X_12097_ _05010_ _05258_ _05260_ _05265_ _05030_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a221o_1
X_16974_ net3508 vssd1 vssd1 vccd1 vccd1 _09987_ sky130_fd_sc_hd__buf_4
X_18713_ _02647_ net4787 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__nand2_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ net6618 net2662 _04392_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
X_15925_ _08559_ _08433_ _08456_ _08560_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__o22ai_2
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ net6071 _03361_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__or2_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15856_ _08898_ _08907_ _08908_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__and3_1
X_18644_ _02630_ _02634_ _02652_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__nand3_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ _07910_ _07957_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__and2_1
XFILLER_0_203_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15787_ _08560_ _08394_ _08841_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__or3_1
X_18575_ _04633_ _02587_ _02588_ _09933_ rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a32o_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _06098_ _06101_ _06096_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__a21o_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914__327 clknet_1_1__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__inv_2
XFILLER_0_15_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17526_ _10523_ _10524_ vssd1 vssd1 vccd1 vccd1 _10525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _07887_ _07888_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__xnor2_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17457_ _10456_ net3474 net4903 vssd1 vssd1 vccd1 vccd1 _10457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14669_ _07801_ _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16408_ _09476_ _09480_ vssd1 vssd1 vccd1 vccd1 _09481_ sky130_fd_sc_hd__xor2_2
X_17388_ _10386_ _10387_ vssd1 vssd1 vccd1 vccd1 _10388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ net4351 _08296_ _09411_ _09412_ _08239_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19127_ net5966 _03052_ _03055_ _03048_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5206 _00901_ vssd1 vssd1 vccd1 vccd1 net5730 sky130_fd_sc_hd__dlygate4sd3_1
X_19058_ net3022 _03009_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__or2_1
Xhold5217 _00706_ vssd1 vssd1 vccd1 vccd1 net5741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5228 net1619 vssd1 vssd1 vccd1 vccd1 net5752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5239 _03423_ vssd1 vssd1 vccd1 vccd1 net5763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4505 rbzero.spi_registers.buf_texadd0\[10\] vssd1 vssd1 vccd1 vccd1 net5029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18009_ _02019_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__xnor2_2
Xhold4516 net784 vssd1 vssd1 vccd1 vccd1 net5040 sky130_fd_sc_hd__dlygate4sd3_1
X_20808__232 clknet_1_0__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__inv_2
Xhold4527 net1275 vssd1 vssd1 vccd1 vccd1 net5051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4538 _00869_ vssd1 vssd1 vccd1 vccd1 net5062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21020_ net1011 net5271 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nor2_1
Xhold4549 _00854_ vssd1 vssd1 vccd1 vccd1 net5073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3804 _03391_ vssd1 vssd1 vccd1 vccd1 net4328 sky130_fd_sc_hd__dlygate4sd3_1
X_20960__369 clknet_1_1__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__inv_2
Xhold3815 _00958_ vssd1 vssd1 vccd1 vccd1 net4339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3826 net7880 vssd1 vssd1 vccd1 vccd1 net4350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3837 net7827 vssd1 vssd1 vccd1 vccd1 net4361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3848 net3114 vssd1 vssd1 vccd1 vccd1 net4372 sky130_fd_sc_hd__buf_1
XFILLER_0_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3859 net7737 vssd1 vssd1 vccd1 vccd1 net4383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21922_ clknet_leaf_6_i_clk net1363 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21853_ clknet_leaf_81_i_clk net3618 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20854__274 clknet_1_0__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__inv_2
XFILLER_0_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21784_ clknet_leaf_76_i_clk _00953_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20735_ clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__buf_1
XFILLER_0_212_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7120 rbzero.traced_texa\[0\] vssd1 vssd1 vccd1 vccd1 net7644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22405_ net157 net2604 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
Xhold7131 rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 net7655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7142 rbzero.spi_registers.buf_texadd3\[23\] vssd1 vssd1 vccd1 vccd1 net7666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7153 rbzero.row_render.texu\[2\] vssd1 vssd1 vccd1 vccd1 net7677 sky130_fd_sc_hd__dlygate4sd3_1
X_20597_ _03924_ net3251 vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__and2_1
Xhold6430 net2269 vssd1 vssd1 vccd1 vccd1 net6954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6441 rbzero.tex_g0\[16\] vssd1 vssd1 vccd1 vccd1 net6965 sky130_fd_sc_hd__dlygate4sd3_1
X_22336_ net468 net2171 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
Xhold6452 net1961 vssd1 vssd1 vccd1 vccd1 net6976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7197 rbzero.traced_texVinit\[10\] vssd1 vssd1 vccd1 vccd1 net7721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6463 rbzero.tex_g1\[61\] vssd1 vssd1 vccd1 vccd1 net6987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6474 net2301 vssd1 vssd1 vccd1 vccd1 net6998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6485 rbzero.tex_b0\[8\] vssd1 vssd1 vccd1 vccd1 net7009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5740 gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 net6264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5751 net2553 vssd1 vssd1 vccd1 vccd1 net6275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22267_ net399 net2019 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
Xhold6496 net2436 vssd1 vssd1 vccd1 vccd1 net7020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5762 gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 net6286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5773 rbzero.spi_registers.buf_texadd3\[0\] vssd1 vssd1 vccd1 vccd1 net6297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5784 rbzero.wall_tracer.mapY\[5\] vssd1 vssd1 vccd1 vccd1 net6308 sky130_fd_sc_hd__dlygate4sd3_1
X_12020_ net4065 net4094 _05188_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o22a_1
X_21218_ clknet_leaf_43_i_clk net5708 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_22198_ net330 net1879 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21149_ net3535 net3981 net2982 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__o21ai_1
X_13971_ _07092_ _07091_ _07089_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__a21o_1
X_15710_ _08778_ _08784_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12922_ net3965 _05825_ _06046_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__mux2_1
X_16690_ _09759_ _09760_ vssd1 vssd1 vccd1 vccd1 _09761_ sky130_fd_sc_hd__nor2_2
XFILLER_0_198_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15641_ _08714_ _08715_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__xnor2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12853_ net53 _05998_ _06010_ _06002_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__a211oi_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _04971_ _04973_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _02396_ net4453 _02338_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15572_ _08642_ _08602_ _08645_ _08646_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__a31o_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _05943_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _10149_ _10188_ _10311_ vssd1 vssd1 vccd1 vccd1 _10312_ sky130_fd_sc_hd__a21oi_2
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ _07655_ _07673_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__nand2_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _09987_ _02334_ _02335_ _09992_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a31o_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _04892_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _10241_ _10242_ vssd1 vssd1 vccd1 vccd1 _10243_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__03980_ _03980_ vssd1 vssd1 vccd1 vccd1 clknet_0__03980_ sky130_fd_sc_hd__clkbuf_16
X_14454_ _07474_ _07358_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__nor2_1
X_11666_ net4971 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ _06485_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__xnor2_2
X_10617_ net1836 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__clkbuf_1
X_17173_ _09096_ _10174_ _10170_ vssd1 vssd1 vccd1 vccd1 _10175_ sky130_fd_sc_hd__o21bai_1
X_14385_ _07533_ _07535_ _07465_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ rbzero.spi_registers.texadd3\[0\] _04640_ _04642_ rbzero.spi_registers.texadd2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _09197_ _09198_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13336_ _06455_ _06445_ _06458_ _06462_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _08517_ _09096_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__or2_1
X_13267_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15006_ _08145_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
X_12218_ rbzero.debug_overlay.facingY\[-8\] _05377_ _05380_ _05386_ vssd1 vssd1 vccd1
+ vccd1 _05387_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _06222_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19814_ net1467 net3151 _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
X_12149_ _05314_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1709 rbzero.tex_g1\[31\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_19745_ net6104 _03407_ net1639 _03413_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__o211a_1
X_16957_ _09971_ _09972_ vssd1 vssd1 vccd1 vccd1 _09973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15908_ _08975_ _08976_ _08982_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__a21bo_1
X_19676_ net6928 _03375_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16888_ _09933_ vssd1 vssd1 vccd1 vccd1 _09937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18627_ net4666 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__clkbuf_4
X_15839_ _08891_ _08894_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__xor2_2
XFILLER_0_149_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ _02572_ rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1 vccd1 _02573_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ _10413_ _10403_ vssd1 vssd1 vccd1 vccd1 _10508_ sky130_fd_sc_hd__or2b_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ net3747 _02504_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or2_1
XANTENNA_13 _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20520_ net3277 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _09286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_46 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_57 _03273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20451_ _03836_ net3558 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__and2_1
XANTENNA_68 rbzero.tex_b0\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20382_ net3428 net1232 _03782_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5003 net1151 vssd1 vssd1 vccd1 vccd1 net5527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5014 net1195 vssd1 vssd1 vccd1 vccd1 net5538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5025 net1147 vssd1 vssd1 vccd1 vccd1 net5549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22121_ net253 net2181 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5036 _00671_ vssd1 vssd1 vccd1 vccd1 net5560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4302 net2389 vssd1 vssd1 vccd1 vccd1 net4826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5047 net3268 vssd1 vssd1 vccd1 vccd1 net5571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5058 net1276 vssd1 vssd1 vccd1 vccd1 net5582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4313 net4794 vssd1 vssd1 vccd1 vccd1 net4837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4324 _01100_ vssd1 vssd1 vccd1 vccd1 net4848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5069 rbzero.spi_registers.texadd2\[1\] vssd1 vssd1 vccd1 vccd1 net5593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4335 rbzero.pov.spi_buffer\[61\] vssd1 vssd1 vccd1 vccd1 net4859 sky130_fd_sc_hd__dlygate4sd3_1
X_22052_ clknet_leaf_90_i_clk net3716 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4346 net1509 vssd1 vssd1 vccd1 vccd1 net4870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3601 _00740_ vssd1 vssd1 vccd1 vccd1 net4125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3612 net7537 vssd1 vssd1 vccd1 vccd1 net4136 sky130_fd_sc_hd__buf_1
Xhold4357 net1302 vssd1 vssd1 vccd1 vccd1 net4881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4368 rbzero.debug_overlay.playerY\[-7\] vssd1 vssd1 vccd1 vccd1 net4892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3623 _00507_ vssd1 vssd1 vccd1 vccd1 net4147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3634 net7486 vssd1 vssd1 vccd1 vccd1 net4158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4379 _10039_ vssd1 vssd1 vccd1 vccd1 net4903 sky130_fd_sc_hd__buf_4
Xhold3645 net674 vssd1 vssd1 vccd1 vccd1 net4169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2900 _03860_ vssd1 vssd1 vccd1 vccd1 net3424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3656 net7553 vssd1 vssd1 vccd1 vccd1 net4180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2911 net1395 vssd1 vssd1 vccd1 vccd1 net3435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2922 net4760 vssd1 vssd1 vccd1 vccd1 net3446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3667 net7646 vssd1 vssd1 vccd1 vccd1 net4191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2944 _03813_ vssd1 vssd1 vccd1 vccd1 net3468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3689 net1219 vssd1 vssd1 vccd1 vccd1 net4213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2955 _01235_ vssd1 vssd1 vccd1 vccd1 net3479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2966 _03915_ vssd1 vssd1 vccd1 vccd1 net3490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2977 net4572 vssd1 vssd1 vccd1 vccd1 net3501 sky130_fd_sc_hd__buf_1
XFILLER_0_138_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2988 _00464_ vssd1 vssd1 vccd1 vccd1 net3512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2999 rbzero.pov.ready_buffer\[71\] vssd1 vssd1 vccd1 vccd1 net3523 sky130_fd_sc_hd__dlygate4sd3_1
X_21905_ clknet_leaf_93_i_clk net1476 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21836_ clknet_leaf_83_i_clk net3860 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20358__88 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__inv_2
X_21767_ clknet_leaf_8_i_clk net2016 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11520_ net7318 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21698_ clknet_leaf_2_i_clk net912 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ net4930 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__clkbuf_4
X_20649_ net1173 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14170_ _07312_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__xnor2_1
X_11382_ net2657 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6260 net2020 vssd1 vssd1 vccd1 vccd1 net6784 sky130_fd_sc_hd__dlygate4sd3_1
X_13121_ net3373 vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__inv_2
Xhold6271 rbzero.tex_r0\[30\] vssd1 vssd1 vccd1 vccd1 net6795 sky130_fd_sc_hd__dlygate4sd3_1
X_22319_ net451 net2062 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6282 net2481 vssd1 vssd1 vccd1 vccd1 net6806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6293 rbzero.tex_r1\[49\] vssd1 vssd1 vccd1 vccd1 net6817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5570 _02659_ vssd1 vssd1 vccd1 vccd1 net6094 sky130_fd_sc_hd__dlygate4sd3_1
X_13052_ _04627_ _06207_ _04626_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__nand3b_4
Xhold5581 _00896_ vssd1 vssd1 vccd1 vccd1 net6105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5592 _02600_ vssd1 vssd1 vccd1 vccd1 net6116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12003_ net3992 _05155_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4880 net1022 vssd1 vssd1 vccd1 vccd1 net5404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17860_ _01808_ _01818_ _01816_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a21o_1
Xhold4891 net1030 vssd1 vssd1 vccd1 vccd1 net5415 sky130_fd_sc_hd__dlygate4sd3_1
X_16811_ _09868_ _09879_ _09880_ vssd1 vssd1 vccd1 vccd1 _09881_ sky130_fd_sc_hd__nand3_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17791_ _01839_ _01840_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__and2_1
X_19530_ net5547 _03288_ _03292_ _03280_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16742_ _09562_ _08707_ _09306_ _08962_ vssd1 vssd1 vccd1 vccd1 _09812_ sky130_fd_sc_hd__a2bb2o_1
X_13954_ net3405 _07084_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _05207_ _06052_ _06046_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a31o_1
X_16673_ _09740_ _09608_ _09305_ vssd1 vssd1 vccd1 vccd1 _09744_ sky130_fd_sc_hd__a21oi_1
X_19461_ net3106 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__clkbuf_1
X_13885_ _06869_ _06973_ _07033_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__or3_4
XFILLER_0_199_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18412_ _02440_ _02441_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__xnor2_1
X_15624_ _08698_ _08490_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ reg_gpout\[3\] clknet_1_1__leaf__05994_ net45 vssd1 vssd1 vccd1 vccd1 _05995_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ net5263 _03198_ _03208_ _03207_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ _08629_ _08611_ _08312_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _02381_ net4491 _02338_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12767_ _04162_ net3993 net16 vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _07652_ _07655_ _07656_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18274_ _02316_ _02319_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__xnor2_1
X_11718_ net1506 _04887_ _04821_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o21a_1
X_15486_ _08559_ _08542_ _08550_ _08560_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ _05207_ _05853_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17225_ _09797_ _10224_ _10225_ vssd1 vssd1 vccd1 vccd1 _10226_ sky130_fd_sc_hd__o21a_1
X_14437_ _07303_ _07304_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__and2_1
Xinput11 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_4
X_11649_ net4930 net4026 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__nand2_1
Xinput22 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_4
Xinput33 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17156_ _08684_ _09477_ vssd1 vssd1 vccd1 vccd1 _10158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_4
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput55 i_vec_csb vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_4
X_14368_ _07504_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__xnor2_1
Xhold806 net5651 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ _08938_ _08944_ _08943_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__a21o_1
Xhold817 net5625 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 net6464 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13319_ _06437_ _06469_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__xnor2_2
X_17087_ _09804_ _09806_ _09802_ vssd1 vssd1 vccd1 vccd1 _10089_ sky130_fd_sc_hd__a21oi_1
Xhold839 _01091_ vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14299_ _07414_ _07449_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16038_ _09082_ _09112_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2207 net7196 vssd1 vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2218 _01351_ vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 net7277 vssd1 vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1506 net6947 vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 _04296_ vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1528 _04558_ vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_17989_ _09231_ _08705_ _02037_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__or3_1
Xhold1539 net6697 vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19728_ net3022 _03407_ net4236 _03400_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19659_ net6170 _03362_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21621_ clknet_leaf_3_i_clk net4114 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21552_ clknet_leaf_5_i_clk net1067 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20503_ net3442 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21483_ clknet_leaf_76_i_clk _00652_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20966__375 clknet_1_0__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__inv_2
X_20434_ net3756 net1288 _03823_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20665__103 clknet_1_1__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__inv_2
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20365_ net3270 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4110 rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 net4634 sky130_fd_sc_hd__buf_2
X_22104_ net236 net2655 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold4121 _03593_ vssd1 vssd1 vccd1 vccd1 net4645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4132 rbzero.debug_overlay.vplaneX\[-8\] vssd1 vssd1 vccd1 vccd1 net4656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4143 _02601_ vssd1 vssd1 vccd1 vccd1 net4667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4154 rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 net4678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4165 net3851 vssd1 vssd1 vccd1 vccd1 net4689 sky130_fd_sc_hd__buf_1
Xhold3420 rbzero.spi_registers.ss_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net3944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3431 _00984_ vssd1 vssd1 vccd1 vccd1 net3955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4176 rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 net4700 sky130_fd_sc_hd__dlygate4sd3_1
X_22035_ clknet_leaf_95_i_clk net3836 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4187 _00605_ vssd1 vssd1 vccd1 vccd1 net4711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3442 _03958_ vssd1 vssd1 vccd1 vccd1 net3966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4198 _02859_ vssd1 vssd1 vccd1 vccd1 net4722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3453 _09915_ vssd1 vssd1 vccd1 vccd1 net3977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3464 _04810_ vssd1 vssd1 vccd1 vccd1 net3988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2730 rbzero.spi_registers.buf_sky\[0\] vssd1 vssd1 vccd1 vccd1 net3254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3475 net6250 vssd1 vssd1 vccd1 vccd1 net3999 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2741 rbzero.wall_tracer.mapX\[5\] vssd1 vssd1 vccd1 vccd1 net3265 sky130_fd_sc_hd__clkbuf_2
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3486 _04613_ vssd1 vssd1 vccd1 vccd1 net4010 sky130_fd_sc_hd__clkbuf_2
Xhold2752 _03890_ vssd1 vssd1 vccd1 vccd1 net3276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3497 _05817_ vssd1 vssd1 vccd1 vccd1 net4021 sky130_fd_sc_hd__buf_4
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2763 _03903_ vssd1 vssd1 vccd1 vccd1 net3287 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2774 _03835_ vssd1 vssd1 vccd1 vccd1 net3298 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2785 rbzero.pov.ready_buffer\[72\] vssd1 vssd1 vccd1 vccd1 net3309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2796 _01184_ vssd1 vssd1 vccd1 vccd1 net3320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ net5856 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13670_ _06662_ _06754_ _06755_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10882_ net2747 net52 _04236_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12621_ _05783_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21819_ clknet_leaf_91_i_clk net4523 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15340_ _08414_ net3003 _06177_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__mux2_1
X_12552_ _05035_ _05712_ _05716_ _05030_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _04652_ _04672_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15271_ _08311_ net7761 _08344_ _08345_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__a2bb2o_2
X_12483_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _05218_ vssd1 vssd1 vccd1 vccd1 _05649_
+ sky130_fd_sc_hd__mux2_1
X_17010_ _10014_ _10017_ _10019_ vssd1 vssd1 vccd1 vccd1 _10020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14222_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _04161_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14153_ net559 net560 vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11365_ net2278 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6090 net1738 vssd1 vssd1 vccd1 vccd1 net6614 sky130_fd_sc_hd__dlygate4sd3_1
X_13104_ _04886_ _06185_ _06196_ net2726 _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14084_ _06865_ _06957_ _06955_ _07232_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__o22a_1
X_18961_ net4634 _05391_ _02917_ _08246_ _02893_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__o311a_1
X_11296_ net1462 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17912_ _01760_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__xnor2_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _06190_ _06178_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__xnor2_1
X_18892_ _02854_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02878_
+ sky130_fd_sc_hd__or2_1
X_17843_ _10380_ _09249_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__nor2_1
X_17774_ _09593_ _10543_ _10541_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__o21ai_4
X_14986_ _06690_ _08120_ _08029_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19513_ net5459 _03274_ _03282_ _03280_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__o211a_1
X_16725_ _09133_ _09794_ vssd1 vssd1 vccd1 vccd1 _09795_ sky130_fd_sc_hd__nand2_1
X_13937_ _07049_ _07048_ _07047_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19444_ net5091 _03036_ _03237_ _03233_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16656_ _08584_ _09086_ _09483_ _09603_ vssd1 vssd1 vccd1 vccd1 _09727_ sky130_fd_sc_hd__or4_1
X_13868_ _07014_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ _08529_ _08449_ _08424_ _08394_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__o22ai_1
X_12819_ net3937 _05957_ _05958_ net3930 _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a221o_1
X_19375_ _03084_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__buf_2
X_16587_ _09553_ _09555_ _09657_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__o21ai_4
X_13799_ _06947_ _06937_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__or2b_1
X_18326_ _02366_ net4591 _02338_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15538_ net3722 _08304_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__nor2_2
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18257_ _08634_ _09538_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__nor2_1
X_15469_ _08300_ net8016 vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17208_ net4540 net4411 vssd1 vssd1 vccd1 vccd1 _10209_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18188_ _02233_ _02234_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nor2_1
Xhold603 net6348 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 net6386 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
X_17139_ _10139_ _10140_ vssd1 vssd1 vccd1 vccd1 _10141_ sky130_fd_sc_hd__xor2_2
XFILLER_0_170_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold625 net6396 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03777_ clknet_0__03777_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03777_
+ sky130_fd_sc_hd__clkbuf_16
Xhold636 net6404 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold647 net5612 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ net3660 _03691_ _03695_ _03696_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__o211a_1
Xhold658 net6354 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 _01372_ vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20081_ net4748 _03577_ _03649_ _03636_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2004 _04428_ vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 _04408_ vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2026 net6993 vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 _01476_ vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2048 _04182_ vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1303 net5739 vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 net6707 vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 _01147_ vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 _00943_ vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1336 _03383_ vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1347 net6719 vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 _01284_ vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 _01557_ vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21604_ clknet_leaf_2_i_clk net4172 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21535_ clknet_leaf_36_i_clk net2468 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21466_ clknet_leaf_24_i_clk net3051 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20351__83 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__inv_2
XFILLER_0_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20417_ net3349 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__clkbuf_1
X_21397_ clknet_leaf_62_i_clk _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11150_ net5920 net5935 _04448_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ net5834 net2024 _04415_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
X_20279_ net3496 _03756_ _03768_ _03761_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__o211a_1
Xhold3250 _00431_ vssd1 vssd1 vccd1 vccd1 net3774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3261 _01205_ vssd1 vssd1 vccd1 vccd1 net3785 sky130_fd_sc_hd__dlygate4sd3_1
X_22018_ clknet_leaf_99_i_clk net3663 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3272 rbzero.wall_tracer.rayAddendX\[2\] vssd1 vssd1 vccd1 vccd1 net3796 sky130_fd_sc_hd__clkbuf_2
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3283 rbzero.debug_overlay.vplaneY\[-4\] vssd1 vssd1 vccd1 vccd1 net3807 sky130_fd_sc_hd__buf_2
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3294 _03789_ vssd1 vssd1 vccd1 vccd1 net3818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2560 _00983_ vssd1 vssd1 vccd1 vccd1 net3084 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ net7434 vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__buf_2
Xhold2571 net6196 vssd1 vssd1 vccd1 vccd1 net3095 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2582 _03249_ vssd1 vssd1 vccd1 vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2593 _03262_ vssd1 vssd1 vccd1 vccd1 net3117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1870 net5887 vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1881 rbzero.tex_r1\[47\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ _07920_ _07921_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__nand2_1
X_11983_ _04161_ _05129_ _05130_ _05131_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o221a_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1892 _04530_ vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
X_16510_ _08684_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13722_ _06868_ _06872_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10934_ net7103 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17490_ _10130_ _09312_ _10488_ vssd1 vssd1 vccd1 vccd1 _10489_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16441_ _09262_ _09396_ _09395_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _06743_ _06707_ _06767_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ net7115 net2695 _04299_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _05051_ _05743_ _05751_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _09350_ _09355_ _09444_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__a21bo_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19160_ _02992_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13584_ _06716_ _06729_ _06732_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a2bb2o_1
X_10796_ net6704 net2759 _04266_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _01986_ _02060_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a21oi_2
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ net4294 _08375_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__xor2_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ net4093 _05693_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091_ _05299_ net3898 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15254_ net7476 _08314_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__nand2_2
X_18042_ _02040_ _02047_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ _05279_ _05631_ _05034_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ _06867_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__clkbuf_4
X_11417_ net5926 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
X_15185_ _08271_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
X_12397_ _04982_ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14136_ _07276_ _07286_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__xor2_1
X_11348_ net6537 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19993_ net3786 net3305 _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__mux2_1
X_14067_ _07192_ _07197_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__xnor2_1
X_18944_ _02910_ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__xnor2_1
X_11279_ net2105 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ _06172_ _06173_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18875_ _02854_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _02862_
+ sky130_fd_sc_hd__xor2_1
X_17826_ _01874_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20660__98 clknet_1_0__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__inv_2
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17757_ _01806_ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14969_ _06721_ _08093_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16708_ _09771_ _09774_ _09772_ vssd1 vssd1 vccd1 vccd1 _09778_ sky130_fd_sc_hd__o21ba_1
X_17688_ _01736_ _01738_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19427_ net5143 _03224_ _03228_ _03220_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__o211a_1
X_16639_ _09700_ _09709_ vssd1 vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19358_ net5750 _03185_ _03189_ _03181_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18309_ _02351_ net4687 _02338_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19289_ net5477 _03146_ _03150_ _03142_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__o211a_1
Xhold6804 _03100_ vssd1 vssd1 vccd1 vccd1 net7328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6815 _00865_ vssd1 vssd1 vccd1 vccd1 net7339 sky130_fd_sc_hd__dlygate4sd3_1
X_21320_ clknet_leaf_72_i_clk _00489_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6837 gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 net7361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6848 rbzero.wall_tracer.stepDistX\[4\] vssd1 vssd1 vccd1 vccd1 net7372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold400 net7487 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
X_21251_ clknet_leaf_51_i_clk net3464 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold411 net3300 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold422 net5380 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20202_ net3412 _03717_ _03725_ _03722_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__o211a_1
Xhold433 net5299 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 rbzero.spi_registers.buf_texadd0\[12\] vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
X_21182_ _03502_ net1128 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nor2_1
Xhold455 net4762 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 net5264 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold477 net5407 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold488 net7520 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
X_20133_ net5551 _03676_ _03686_ _03683_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__o211a_1
Xhold499 net4247 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
X_20064_ net4640 _03581_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__or2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 net4730 vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _03082_ vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20777__204 clknet_1_0__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__inv_2
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _00918_ vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 net4228 vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _03366_ vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 _01499_ vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 _03438_ vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 net4673 vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 net6061 vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 net6651 vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ net6566 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12320_ _05486_ _05487_ _05068_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21518_ clknet_leaf_33_i_clk net1636 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12251_ rbzero.debug_overlay.playerY\[-2\] _05374_ _05372_ net3917 vssd1 vssd1 vccd1
+ vccd1 _05420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21449_ clknet_leaf_45_i_clk net3924 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ net6738 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12182_ _05341_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11133_ net6656 net2521 _04437_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ _09999_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10002_ sky130_fd_sc_hd__or3_2
X_11064_ net6449 net1765 _04404_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__mux2_1
X_15941_ _08955_ _08956_ _08965_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__o21ai_1
Xhold3080 net4669 vssd1 vssd1 vccd1 vccd1 net3604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3091 rbzero.pov.ready_buffer\[4\] vssd1 vssd1 vccd1 vccd1 net3615 sky130_fd_sc_hd__dlygate4sd3_1
X_18660_ _02637_ net4463 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__xor2_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _08909_ _08935_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__xnor2_2
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2390 rbzero.pov.ready_buffer\[51\] vssd1 vssd1 vccd1 vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
X_17611_ _10486_ _10495_ _10493_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _07572_ _07973_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__nor2_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18591_ _02594_ _02595_ _02596_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17542_ _09138_ _09139_ _10168_ vssd1 vssd1 vccd1 vccd1 _10541_ sky130_fd_sc_hd__or3_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14754_ _07367_ _07805_ _07904_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__or3_1
X_11966_ net2993 _05125_ net1793 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__o21ai_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ net5931 net2253 _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _06847_ _06850_ _06855_ _06733_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__o22ai_2
X_17473_ _10355_ _10370_ _10368_ vssd1 vssd1 vccd1 vccd1 _10472_ sky130_fd_sc_hd__a21o_1
X_14685_ _07812_ _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__xor2_2
XFILLER_0_184_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _05037_ vssd1 vssd1 vccd1 vccd1 _05067_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19212_ _03036_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__clkbuf_4
X_16424_ _09492_ _09496_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__xnor2_2
X_13636_ _06743_ _06785_ _06786_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__or3b_1
X_10848_ net7058 net6702 _04288_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19143_ net5216 _03053_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__or2_1
X_16355_ _09425_ _09426_ vssd1 vssd1 vccd1 vccd1 _09428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ _06697_ _06698_ _06600_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ net6489 net2499 _04255_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20315__50 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12518_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _05218_ vssd1 vssd1 vccd1 vccd1 _05684_
+ sky130_fd_sc_hd__mux2_1
X_15306_ net7404 vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ _08559_ _09222_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19074_ net642 net2979 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13498_ _06628_ _06630_ _06643_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__or4b_2
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18025_ net4497 net4619 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ _08311_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__buf_6
X_12449_ reg_rgb\[15\] _05615_ _05204_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__mux2_2
XFILLER_0_125_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20330__64 clknet_1_1__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4709 net1433 vssd1 vssd1 vccd1 vccd1 net5233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15168_ _08262_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _07267_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__xor2_1
X_20726__158 clknet_1_1__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__inv_2
X_19976_ net3422 _03578_ net4364 _03550_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__o211a_1
X_15099_ _08190_ net3067 net6279 _08215_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18927_ _02864_ _05391_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18858_ _02844_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17809_ _01739_ _01746_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__nor2_1
X_18789_ _02779_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22421_ clknet_leaf_57_i_clk net4977 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7302 net4434 vssd1 vssd1 vccd1 vccd1 net7826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6601 net2711 vssd1 vssd1 vccd1 vccd1 net7125 sky130_fd_sc_hd__dlygate4sd3_1
X_22352_ net484 net2339 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold6612 rbzero.tex_b0\[13\] vssd1 vssd1 vccd1 vccd1 net7136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7357 net4350 vssd1 vssd1 vccd1 vccd1 net7881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6623 _02715_ vssd1 vssd1 vccd1 vccd1 net7147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7368 rbzero.wall_tracer.stepDistY\[8\] vssd1 vssd1 vccd1 vccd1 net7892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6634 _04324_ vssd1 vssd1 vccd1 vccd1 net7158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5900 rbzero.tex_b1\[45\] vssd1 vssd1 vccd1 vccd1 net6424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21303_ clknet_leaf_47_i_clk _00472_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold6645 net2728 vssd1 vssd1 vccd1 vccd1 net7169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5911 net1207 vssd1 vssd1 vccd1 vccd1 net6435 sky130_fd_sc_hd__dlygate4sd3_1
X_22283_ net415 net1122 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold6656 rbzero.tex_r1\[52\] vssd1 vssd1 vccd1 vccd1 net7180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5922 _04230_ vssd1 vssd1 vccd1 vccd1 net6446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6667 net2622 vssd1 vssd1 vccd1 vccd1 net7191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6678 rbzero.tex_r0\[47\] vssd1 vssd1 vccd1 vccd1 net7202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5933 net1332 vssd1 vssd1 vccd1 vccd1 net6457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5944 rbzero.tex_b0\[46\] vssd1 vssd1 vccd1 vccd1 net6468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6689 net2737 vssd1 vssd1 vccd1 vccd1 net7213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5955 net1418 vssd1 vssd1 vccd1 vccd1 net6479 sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ clknet_leaf_59_i_clk _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold230 net4996 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold241 net5025 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5966 _04261_ vssd1 vssd1 vccd1 vccd1 net6490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 net4980 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5977 _04294_ vssd1 vssd1 vccd1 vccd1 net6501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5988 net1427 vssd1 vssd1 vccd1 vccd1 net6512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 net5046 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5999 rbzero.spi_registers.buf_floor\[4\] vssd1 vssd1 vccd1 vccd1 net6523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _03324_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_2
X_21165_ _04139_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__buf_1
Xhold285 net5196 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 net5077 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
X_20116_ net4845 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__buf_4
X_21096_ net4936 net1886 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__nand2_1
X_20047_ net3177 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _04989_ vssd1 vssd1 vccd1 vccd1 _04990_
+ sky130_fd_sc_hd__mux2_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ net223 net1969 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _04918_ _04919_ net2909 vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ net2827 net6359 _04214_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__mux2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _07444_ _07439_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__nor2_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _04599_ _04602_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nor2_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20831__253 clknet_1_0__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__inv_2
XFILLER_0_181_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13421_ _06547_ _06549_ _06539_ _06550_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__and4_1
XFILLER_0_187_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10633_ net2602 net7153 _04181_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16140_ _09207_ _09214_ vssd1 vssd1 vccd1 vccd1 _09215_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _04635_ _06500_ _06502_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12303_ _05030_ _05455_ _05462_ _05470_ _05051_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__o311a_1
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16071_ _09140_ _09145_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__nor2_1
X_13283_ net6259 _06430_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ net7458 _08157_ _08158_ _08068_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ net4656 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19830_ net41 net40 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__or2_2
X_12165_ net4071 _05330_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a21o_1
X_11116_ net2666 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
X_19761_ net1572 _03427_ net1560 _03424_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__o211a_1
X_12096_ _05261_ _05264_ _05034_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16973_ _09965_ _09985_ _09986_ _09966_ net5420 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18712_ _02647_ net4787 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__or2_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net1996 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
X_15924_ _08387_ _08493_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__nor2_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_102_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19692_ net4401 _03359_ net1713 _03384_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__o211a_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ _02650_ _02651_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__or2_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _08869_ _08911_ _08928_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__a21o_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _07907_ _07909_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__or2_1
X_18574_ net3838 _02586_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15786_ _08857_ _08860_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__nand2_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _06153_ _06102_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nand2_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _10514_ _10522_ vssd1 vssd1 vccd1 vccd1 _10524_ sky130_fd_sc_hd__or2_1
X_14737_ _07532_ _07590_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__nor2_1
X_11949_ _04909_ _05053_ _05094_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17456_ _09987_ _10336_ _10337_ _10455_ vssd1 vssd1 vccd1 vccd1 _10456_ sky130_fd_sc_hd__a31o_1
X_14668_ _07444_ _07524_ _07800_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16407_ _09478_ _09479_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__xor2_2
XFILLER_0_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _06697_ _06698_ _06621_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__a21oi_1
X_17387_ _08872_ _09595_ vssd1 vssd1 vccd1 vccd1 _10387_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ _07705_ _07708_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19126_ net5132 _03053_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__or2_1
X_16338_ net7407 _09410_ _08633_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19057_ net3022 net2843 _03012_ _03011_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__o211a_1
Xhold5207 net1573 vssd1 vssd1 vccd1 vccd1 net5731 sky130_fd_sc_hd__dlygate4sd3_1
X_16269_ _09341_ _09342_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__nor2_1
Xhold5218 rbzero.spi_registers.texadd0\[3\] vssd1 vssd1 vccd1 vccd1 net5742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5229 rbzero.spi_registers.buf_leak\[1\] vssd1 vssd1 vccd1 vccd1 net5753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18008_ _02055_ _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__nor2_1
Xhold4506 net703 vssd1 vssd1 vccd1 vccd1 net5030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4517 rbzero.spi_registers.texadd0\[20\] vssd1 vssd1 vccd1 vccd1 net5041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4528 rbzero.spi_registers.texadd1\[15\] vssd1 vssd1 vccd1 vccd1 net5052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4539 net759 vssd1 vssd1 vccd1 vccd1 net5063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3805 _00921_ vssd1 vssd1 vccd1 vccd1 net4329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3816 net3033 vssd1 vssd1 vccd1 vccd1 net4340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3827 net1189 vssd1 vssd1 vccd1 vccd1 net4351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3838 net3065 vssd1 vssd1 vccd1 vccd1 net4362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3849 net7816 vssd1 vssd1 vccd1 vccd1 net4373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19959_ _03470_ _03564_ _03531_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21921_ clknet_leaf_93_i_clk net1401 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21852_ clknet_leaf_81_i_clk net3677 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21783_ clknet_leaf_31_i_clk net3928 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20889__305 clknet_1_0__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__inv_2
XFILLER_0_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7110 rbzero.spi_registers.texadd0\[12\] vssd1 vssd1 vccd1 vccd1 net7634 sky130_fd_sc_hd__dlygate4sd3_1
X_22404_ net156 net2139 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
Xhold7121 rbzero.pov.ready_buffer\[27\] vssd1 vssd1 vccd1 vccd1 net7645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7132 rbzero.spi_registers.texadd2\[15\] vssd1 vssd1 vccd1 vccd1 net7656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7143 rbzero.spi_registers.buf_texadd1\[19\] vssd1 vssd1 vccd1 vccd1 net7667 sky130_fd_sc_hd__dlygate4sd3_1
X_20596_ net3156 net1187 net3250 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__mux2_1
Xhold7154 rbzero.pov.ready_buffer\[30\] vssd1 vssd1 vccd1 vccd1 net7678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6420 net2445 vssd1 vssd1 vccd1 vccd1 net6944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6431 rbzero.tex_b0\[36\] vssd1 vssd1 vccd1 vccd1 net6955 sky130_fd_sc_hd__dlygate4sd3_1
X_22335_ net467 net2624 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6442 net1935 vssd1 vssd1 vccd1 vccd1 net6966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7187 rbzero.traced_texVinit\[1\] vssd1 vssd1 vccd1 vccd1 net7711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6453 rbzero.tex_b0\[15\] vssd1 vssd1 vccd1 vccd1 net6977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7198 net4230 vssd1 vssd1 vccd1 vccd1 net7722 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold6464 net2057 vssd1 vssd1 vccd1 vccd1 net6988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6475 _04391_ vssd1 vssd1 vccd1 vccd1 net6999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5730 _08214_ vssd1 vssd1 vccd1 vccd1 net6254 sky130_fd_sc_hd__dlygate4sd3_1
X_22266_ net398 net2832 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
Xhold6486 net2215 vssd1 vssd1 vccd1 vccd1 net7010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5741 net3897 vssd1 vssd1 vccd1 vccd1 net6265 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold6497 rbzero.tex_g1\[10\] vssd1 vssd1 vccd1 vccd1 net7021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5752 _03269_ vssd1 vssd1 vccd1 vccd1 net6276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5763 net3964 vssd1 vssd1 vccd1 vccd1 net6287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5774 net1559 vssd1 vssd1 vccd1 vccd1 net6298 sky130_fd_sc_hd__dlygate4sd3_1
X_21217_ clknet_leaf_43_i_clk net4826 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5785 net3034 vssd1 vssd1 vccd1 vccd1 net6309 sky130_fd_sc_hd__dlygate4sd3_1
X_22197_ net329 net2239 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold5796 _02944_ vssd1 vssd1 vccd1 vccd1 net6320 sky130_fd_sc_hd__dlygate4sd3_1
X_21148_ net3535 net3981 _08195_ net3507 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__o211a_1
X_21079_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__inv_2
X_13970_ _07092_ _07089_ _07091_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__nand3_1
X_12921_ net37 net36 _06077_ net38 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__a31o_1
XFILLER_0_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15640_ _08456_ _08498_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__nor2_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ net40 _06007_ _06008_ net41 _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a221o_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _04962_ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__xnor2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _08596_ _08597_ _08613_ _08644_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ reg_gpout\[2\] clknet_1_1__leaf__05942_ net45 vssd1 vssd1 vccd1 vccd1 _05943_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_150_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _10186_ _10187_ vssd1 vssd1 vccd1 vccd1 _10311_ sky130_fd_sc_hd__nor2_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _07652_ _07653_ _07654_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__a21o_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11734_ net3620 _04164_ _04759_ _04894_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a221o_1
X_18290_ net4475 net4315 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__or2_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17241_ _10132_ _10134_ _10240_ vssd1 vssd1 vccd1 vccd1 _10242_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14453_ _07602_ _07603_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__nand2_2
X_11665_ net3921 _04600_ _04606_ net3821 _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10616_ net6516 net6902 _04170_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13404_ _06540_ net82 _06517_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__o21ai_2
X_17172_ _10172_ _10173_ vssd1 vssd1 vccd1 vccd1 _10174_ sky130_fd_sc_hd__and2_2
XFILLER_0_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14384_ _07534_ _07532_ _07464_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11596_ _04718_ _04764_ _04767_ _04727_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__o31a_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16123_ _08433_ _08498_ _08733_ _08731_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ _06449_ _06450_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__nand2_1
X_16054_ _09098_ _09128_ vssd1 vssd1 vccd1 vccd1 _09129_ sky130_fd_sc_hd__nand2_1
X_13266_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__xor2_4
XFILLER_0_84_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12217_ rbzero.debug_overlay.facingY\[-1\] _05381_ _05382_ rbzero.debug_overlay.facingY\[-9\]
+ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a221o_1
X_15005_ net4451 _08144_ _08138_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__mux2_1
X_13197_ _04868_ net3984 _06185_ _06350_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__a221o_1
XFILLER_0_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19813_ net3971 net2978 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__nand2_2
X_12148_ _04836_ _04603_ _05315_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19744_ net1638 _03408_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ _04992_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__buf_4
X_16956_ net4922 _09968_ vssd1 vssd1 vccd1 vccd1 _09972_ sky130_fd_sc_hd__nor2_1
X_15907_ _08977_ _08974_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19675_ net3088 _03374_ net1693 _03371_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16887_ net4391 _09934_ _09936_ _08144_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a22o_1
X_18626_ _02621_ _02632_ _02633_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a31o_1
X_20838__259 clknet_1_1__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__inv_2
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _08844_ _08852_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18557_ net3241 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__buf_1
X_15769_ _08840_ _08843_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17508_ _10405_ _10412_ vssd1 vssd1 vccd1 vccd1 _10507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18488_ _02504_ _02508_ net3211 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a21oi_1
X_17439_ _10437_ _10438_ vssd1 vssd1 vccd1 vccd1 _10439_ sky130_fd_sc_hd__nor2_1
XANTENNA_14 _05069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_36 _10205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20450_ net1098 net3557 _03823_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__mux2_1
XANTENNA_58 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 rbzero.wall_tracer.visualWallDist\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19109_ net5402 _03040_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20381_ net3191 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5004 _00772_ vssd1 vssd1 vccd1 vccd1 net5528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5015 rbzero.pov.spi_buffer\[18\] vssd1 vssd1 vccd1 vccd1 net5539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22120_ net252 net2414 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold5026 rbzero.pov.spi_buffer\[5\] vssd1 vssd1 vccd1 vccd1 net5550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5037 rbzero.spi_registers.buf_otherx\[2\] vssd1 vssd1 vccd1 vccd1 net5561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4303 net688 vssd1 vssd1 vccd1 vccd1 net4827 sky130_fd_sc_hd__buf_1
Xhold5048 _03681_ vssd1 vssd1 vccd1 vccd1 net5572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4314 _03677_ vssd1 vssd1 vccd1 vccd1 net4838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5059 _01053_ vssd1 vssd1 vccd1 vccd1 net5583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4325 net4859 vssd1 vssd1 vccd1 vccd1 net4849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22051_ clknet_leaf_90_i_clk net3576 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4336 rbzero.pov.spi_buffer\[73\] vssd1 vssd1 vccd1 vccd1 net4860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3602 net620 vssd1 vssd1 vccd1 vccd1 net4126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3613 _00519_ vssd1 vssd1 vccd1 vccd1 net4137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4358 _01107_ vssd1 vssd1 vccd1 vccd1 net4882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4369 net2940 vssd1 vssd1 vccd1 vccd1 net4893 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3624 net693 vssd1 vssd1 vccd1 vccd1 net4148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3635 net924 vssd1 vssd1 vccd1 vccd1 net4159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2901 _01209_ vssd1 vssd1 vccd1 vccd1 net3425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3646 net7636 vssd1 vssd1 vccd1 vccd1 net4170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3657 net687 vssd1 vssd1 vccd1 vccd1 net4181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2912 _03896_ vssd1 vssd1 vccd1 vccd1 net3436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2923 net4506 vssd1 vssd1 vccd1 vccd1 net3447 sky130_fd_sc_hd__buf_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3668 _00754_ vssd1 vssd1 vccd1 vccd1 net4192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3679 net7506 vssd1 vssd1 vccd1 vccd1 net4203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2934 net6108 vssd1 vssd1 vccd1 vccd1 net3458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2945 _01188_ vssd1 vssd1 vccd1 vccd1 net3469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2967 _01234_ vssd1 vssd1 vccd1 vccd1 net3491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2978 net4574 vssd1 vssd1 vccd1 vccd1 net3502 sky130_fd_sc_hd__buf_1
Xhold2989 net4858 vssd1 vssd1 vccd1 vccd1 net3513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21904_ clknet_leaf_93_i_clk net1342 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21835_ clknet_leaf_83_i_clk net4603 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21766_ clknet_leaf_18_i_clk net5840 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21697_ clknet_leaf_3_i_clk net4117 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ net3402 net2982 net3507 _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__o31ai_1
X_20648_ net6363 _03026_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11381_ net7211 net6970 _04573_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20579_ _03924_ net3680 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6250 net2305 vssd1 vssd1 vccd1 vccd1 net6774 sky130_fd_sc_hd__dlygate4sd3_1
X_13120_ net3284 vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__inv_2
X_22318_ net450 net1761 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold6261 rbzero.tex_r1\[22\] vssd1 vssd1 vccd1 vccd1 net6785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6272 net2060 vssd1 vssd1 vccd1 vccd1 net6796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6283 _04571_ vssd1 vssd1 vccd1 vccd1 net6807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6294 net2066 vssd1 vssd1 vccd1 vccd1 net6818 sky130_fd_sc_hd__dlygate4sd3_1
X_20943__354 clknet_1_0__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__inv_2
X_13051_ net4909 net6168 vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__nor2b_2
X_22249_ net381 net1429 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5571 net3371 vssd1 vssd1 vccd1 vccd1 net6095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5582 net1770 vssd1 vssd1 vccd1 vccd1 net6106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5593 net3595 vssd1 vssd1 vccd1 vccd1 net6117 sky130_fd_sc_hd__dlygate4sd3_1
X_12002_ _04161_ _05158_ _05171_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__o21ai_1
Xhold4870 rbzero.spi_registers.texadd0\[15\] vssd1 vssd1 vccd1 vccd1 net5394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4881 rbzero.spi_registers.buf_othery\[1\] vssd1 vssd1 vccd1 vccd1 net5405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4892 rbzero.spi_registers.texadd0\[16\] vssd1 vssd1 vccd1 vccd1 net5416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16810_ _09875_ _09876_ _09878_ vssd1 vssd1 vccd1 vccd1 _09880_ sky130_fd_sc_hd__a21o_1
X_17790_ _01839_ _01840_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16741_ _09810_ _09699_ _09697_ vssd1 vssd1 vccd1 vccd1 _09811_ sky130_fd_sc_hd__a21o_1
X_13953_ _07102_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_202_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19460_ _03088_ net3105 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__or2_1
X_12904_ _06046_ _06052_ net41 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__and3b_1
X_16672_ _09734_ _09742_ vssd1 vssd1 vccd1 vccd1 _09743_ sky130_fd_sc_hd__xor2_1
XFILLER_0_159_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _07033_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__xnor2_2
X_18411_ _02432_ _02434_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
X_15623_ _08313_ _08315_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ net1559 _03199_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__or2_1
X_12835_ _05446_ _05948_ _05954_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__o22a_2
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ net7818 _02380_ _10047_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__o21ai_1
X_15554_ net3120 _08628_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__nand2_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _05923_ _05925_ net19 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__mux2_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _07605_ _07608_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18273_ _02317_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11717_ net2791 net2789 net2879 net2802 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__or4_1
X_15485_ _08367_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__clkbuf_4
X_12697_ net40 _05852_ _05854_ net41 vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17224_ _09328_ _09419_ _09794_ _09051_ vssd1 vssd1 vccd1 vccd1 _10225_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14436_ _06859_ _07524_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__nor2_1
X_11648_ net4909 net6168 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nand2_4
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
Xinput23 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_2
Xinput34 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_4
X_17155_ _10155_ _10156_ vssd1 vssd1 vccd1 vccd1 _10157_ sky130_fd_sc_hd__xnor2_2
Xinput45 i_reg_outs_enb vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_4
XFILLER_0_13_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14367_ _07508_ _07513_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__o21a_1
X_11579_ _04674_ _04652_ _04672_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput56 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_4
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold807 net5653 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ _08945_ _08996_ _09178_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__a22o_4
Xhold818 net5627 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ _06465_ _06468_ _06466_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a21o_1
X_17086_ _09828_ _09793_ vssd1 vssd1 vccd1 vccd1 _10088_ sky130_fd_sc_hd__or2b_1
Xhold829 net6466 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ _07082_ _07419_ _06931_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16037_ _09083_ _09101_ _09111_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ net2768 net2388 _06179_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2208 net7198 vssd1 vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2219 net7238 vssd1 vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1507 net6949 vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1518 _01475_ vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
X_17988_ _02035_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1529 _01145_ vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19727_ net4235 _03408_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__or2_1
X_16939_ _09949_ _09955_ _09956_ vssd1 vssd1 vccd1 vccd1 _09957_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19658_ net3112 _03360_ net2275 _03354_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18609_ net87 _02613_ _02619_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19589_ _03294_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21620_ clknet_leaf_3_i_clk net4120 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21551_ clknet_leaf_3_i_clk net4129 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20502_ _03858_ net3441 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21482_ clknet_leaf_21_i_clk net2950 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20433_ net3293 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20364_ _08279_ net3269 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__and2_1
Xhold4100 net739 vssd1 vssd1 vccd1 vccd1 net4624 sky130_fd_sc_hd__dlygate4sd3_1
X_22103_ net235 net762 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4111 _03650_ vssd1 vssd1 vccd1 vccd1 net4635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4122 _00992_ vssd1 vssd1 vccd1 vccd1 net4646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4133 _02534_ vssd1 vssd1 vccd1 vccd1 net4657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4144 _02604_ vssd1 vssd1 vccd1 vccd1 net4668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4155 net2158 vssd1 vssd1 vccd1 vccd1 net4679 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3410 _02998_ vssd1 vssd1 vccd1 vccd1 net3934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4166 net4771 vssd1 vssd1 vccd1 vccd1 net4690 sky130_fd_sc_hd__dlygate4sd3_1
X_22034_ clknet_leaf_96_i_clk net3654 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3421 net2841 vssd1 vssd1 vccd1 vccd1 net3945 sky130_fd_sc_hd__buf_1
XFILLER_0_140_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4177 net1364 vssd1 vssd1 vccd1 vccd1 net4701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3432 rbzero.spi_registers.spi_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net3956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4188 net3863 vssd1 vssd1 vccd1 vccd1 net4712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3443 _01255_ vssd1 vssd1 vccd1 vccd1 net3967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3454 _09916_ vssd1 vssd1 vccd1 vccd1 net3978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4199 _02861_ vssd1 vssd1 vccd1 vccd1 net4723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2720 _03632_ vssd1 vssd1 vccd1 vccd1 net3244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3465 _04811_ vssd1 vssd1 vccd1 vccd1 net3989 sky130_fd_sc_hd__clkbuf_2
Xhold2731 _03242_ vssd1 vssd1 vccd1 vccd1 net3255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3476 _00616_ vssd1 vssd1 vccd1 vccd1 net4000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3487 _05348_ vssd1 vssd1 vccd1 vccd1 net4011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2742 net6142 vssd1 vssd1 vccd1 vccd1 net3266 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2753 _03891_ vssd1 vssd1 vccd1 vccd1 net3277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3498 _03963_ vssd1 vssd1 vccd1 vccd1 net4022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2764 _03904_ vssd1 vssd1 vccd1 vccd1 net3288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2775 _01198_ vssd1 vssd1 vccd1 vccd1 net3299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2786 net1034 vssd1 vssd1 vccd1 vccd1 net3310 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2797 net4482 vssd1 vssd1 vccd1 vccd1 net3321 sky130_fd_sc_hd__dlygate4sd3_1
X_10950_ net2234 net5854 _04344_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10881_ net5777 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire80 _05008_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_2
XFILLER_0_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ reg_hsync _05782_ _05204_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__mux2_2
XFILLER_0_211_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21818_ clknet_leaf_91_i_clk net4445 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _05004_ _05713_ _05715_ _05010_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21749_ clknet_leaf_102_i_clk net1646 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _04650_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nand2_1
X_12482_ _05019_ _05647_ _05009_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__o21a_1
X_15270_ net4306 _08341_ _06209_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14221_ _07365_ _07370_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11433_ _04164_ _04603_ _04607_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__o31a_1
XFILLER_0_184_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _07251_ _07253_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__xnor2_1
X_11364_ net6804 net6508 _04562_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6080 net1664 vssd1 vssd1 vccd1 vccd1 net6604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6091 _04539_ vssd1 vssd1 vccd1 vccd1 net6615 sky130_fd_sc_hd__dlygate4sd3_1
X_13103_ net2791 _06183_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__xnor2_1
X_14083_ _07214_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__or2_1
X_18960_ _02939_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__xnor2_1
X_11295_ net6506 net5953 _04529_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17911_ _01958_ _01960_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__xor2_1
Xhold5390 rbzero.tex_r1\[28\] vssd1 vssd1 vccd1 vccd1 net5914 sky130_fd_sc_hd__dlygate4sd3_1
X_13034_ net3804 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__inv_2
X_18891_ _02854_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02877_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17842_ _01675_ _08793_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__or2_1
XFILLER_0_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17773_ _01702_ _01704_ _01701_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a21bo_1
X_14985_ _06663_ _08030_ _08032_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19512_ net1572 _03275_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__or2_1
X_16724_ _09305_ _09536_ vssd1 vssd1 vccd1 vccd1 _09794_ sky130_fd_sc_hd__nor2_1
X_13936_ _07049_ _07047_ _07048_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19443_ net2873 _03039_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__or2_1
X_16655_ _09718_ _09725_ vssd1 vssd1 vccd1 vccd1 _09726_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ _07016_ _07017_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15606_ _08529_ _08393_ _08405_ _08422_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__or4_1
X_19374_ _03035_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__clkbuf_4
X_12818_ net4972 _05946_ _05956_ net4002 vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__a22o_1
X_16586_ _09542_ _09556_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _06908_ _06909_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__xor2_2
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18325_ net7782 _02365_ _10029_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15537_ net3539 _08327_ _08379_ _08611_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__or4_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ net40 _05903_ _05905_ net41 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18256_ _02180_ _02301_ _02197_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15468_ _08130_ _08137_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ _10208_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__clkbuf_1
X_14419_ _07504_ _07518_ _07569_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__o21a_1
X_18187_ _02205_ _02232_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__nor2_1
X_15399_ net4358 _08434_ net4288 vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17138_ _08873_ _08582_ vssd1 vssd1 vccd1 vccd1 _10140_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold604 _04142_ vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 net6388 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__03776_ clknet_0__03776_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03776_
+ sky130_fd_sc_hd__clkbuf_16
Xhold626 _01512_ vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold637 _01482_ vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 net6362 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
X_17069_ _10070_ _10071_ _10072_ vssd1 vssd1 vccd1 vccd1 _10073_ sky130_fd_sc_hd__o21ai_1
Xhold659 _04156_ vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20080_ _05391_ _03581_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__or2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _01357_ vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 _01375_ vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 net6995 vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2038 net5910 vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1304 net5741 vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2049 _01576_ vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 net6709 vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1326 net6669 vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1337 net6030 vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1348 _03434_ vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 net6235 vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20972__380 clknet_1_1__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__inv_2
XFILLER_0_71_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21603_ clknet_leaf_102_i_clk net5529 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21534_ clknet_leaf_36_i_clk net2195 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21465_ clknet_leaf_24_i_clk net3113 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20416_ _03814_ net3348 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21396_ clknet_leaf_61_i_clk _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ net5987 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20278_ net3514 net4839 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3240 rbzero.pov.ready_buffer\[31\] vssd1 vssd1 vccd1 vccd1 net3764 sky130_fd_sc_hd__buf_1
X_22017_ clknet_leaf_98_i_clk net3609 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3251 rbzero.pov.ready_buffer\[38\] vssd1 vssd1 vccd1 vccd1 net3775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3262 rbzero.debug_overlay.facingX\[-1\] vssd1 vssd1 vccd1 vccd1 net3786 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3273 net6326 vssd1 vssd1 vccd1 vccd1 net3797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3284 _03644_ vssd1 vssd1 vccd1 vccd1 net3808 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2550 net7311 vssd1 vssd1 vccd1 vccd1 net3074 sky130_fd_sc_hd__clkbuf_2
Xhold3295 _03790_ vssd1 vssd1 vccd1 vccd1 net3819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2561 rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 net3085 sky130_fd_sc_hd__clkbuf_2
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 net3052 vssd1 vssd1 vccd1 vccd1 net3096 sky130_fd_sc_hd__buf_4
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2583 _00806_ vssd1 vssd1 vccd1 vccd1 net3107 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2594 _03263_ vssd1 vssd1 vccd1 vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1860 _01528_ vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1871 _01526_ vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
X_14770_ _07532_ _07805_ _07919_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1882 net7007 vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
X_11982_ net4041 _05133_ _05129_ _04161_ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a221o_1
Xhold1893 _01171_ vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
X_13721_ _06870_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__xnor2_2
X_10933_ net2674 net7101 _04333_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16440_ _09414_ _09512_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10864_ net6826 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__clkbuf_1
X_13652_ _06800_ _06802_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12603_ _04979_ _05755_ _05759_ _05028_ _05767_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__o311a_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _09356_ _09349_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ net2422 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__clkbuf_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ net7433 _06715_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__nor2_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18110_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__nor2_1
X_15322_ _08374_ _08395_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__a21bo_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _05699_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
X_19090_ net4020 net3897 net3964 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18041_ _02045_ _02046_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ _08327_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12465_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _05457_ vssd1 vssd1 vccd1 vccd1 _05631_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_90 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_90/HI o_rgb[0] sky130_fd_sc_hd__conb_1
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14204_ _06859_ _07354_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__or2_1
X_11416_ net5924 net5767 _04243_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__mux2_1
X_12396_ rbzero.tex_g1\[47\] rbzero.tex_g1\[46\] _04987_ vssd1 vssd1 vccd1 vccd1 _05563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15184_ net4619 _08184_ _08260_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__mux2_1
X_11347_ net6535 net2331 _04551_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_1
X_14135_ _07277_ _07285_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19992_ _03580_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11278_ net5890 net6780 _04514_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
X_14066_ _07209_ _07214_ _07216_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__o21a_1
X_18943_ _02924_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13017_ _06122_ _06140_ _06141_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__and3_1
X_18874_ net1581 _02557_ _02853_ net4723 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__o211ai_1
X_17825_ _01795_ _01872_ _01873_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _01804_ _01805_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__or2_1
X_14968_ _08069_ _08111_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__nand2_1
X_16707_ net4519 _08296_ _09776_ _09777_ _08239_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13919_ _07042_ _07068_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__a21oi_1
X_17687_ _01736_ _01738_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14899_ net4310 _08048_ _08027_ vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19426_ net1543 _03225_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__or2_1
X_16638_ _09707_ _09708_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19357_ net1806 _03186_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__or2_1
X_16569_ _09529_ _09640_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18308_ _06206_ net7805 _10011_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19288_ net1667 _03147_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18239_ _02188_ _02283_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6805 rbzero.pov.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 net7329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6827 _03591_ vssd1 vssd1 vccd1 vccd1 net7351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6838 _04815_ vssd1 vssd1 vccd1 vccd1 net7362 sky130_fd_sc_hd__dlygate4sd3_1
X_21250_ clknet_leaf_50_i_clk net3264 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6849 net3272 vssd1 vssd1 vccd1 vccd1 net7373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold401 net5135 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold412 net4563 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 net5355 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
X_20201_ net5533 _03718_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold434 net5181 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold445 net609 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
X_21181_ net6349 net4951 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold456 net4764 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 net5301 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
X_20132_ net3737 _03679_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__or2_1
Xhold478 net5286 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 rbzero.pov.ready_buffer\[67\] vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20063_ net4729 _03613_ _03638_ _03636_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__o211a_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 net6561 vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
X_20703__137 clknet_1_1__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__inv_2
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 net5997 vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1123 net6585 vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 net6617 vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 _00880_ vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 net6581 vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 net6173 vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 _00897_ vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 net6063 vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21517_ clknet_leaf_37_i_clk net5704 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _05194_ _05418_ net4014 _05193_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21448_ clknet_leaf_45_i_clk net3986 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ net1923 net6736 _04481_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12181_ _05348_ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__nand2_1
X_21379_ clknet_leaf_66_i_clk _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ net2117 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
Xhold990 _01429_ vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ net2219 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
X_15940_ _08955_ _08956_ _08965_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__or3_1
Xhold3081 rbzero.pov.ready_buffer\[11\] vssd1 vssd1 vccd1 vccd1 net3605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3092 _03642_ vssd1 vssd1 vccd1 vccd1 net3616 sky130_fd_sc_hd__dlygate4sd3_1
X_15871_ _08938_ _08945_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__nand2_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2380 _01485_ vssd1 vssd1 vccd1 vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
X_17610_ _10597_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__xnor2_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2391 _03549_ vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
X_14822_ _07562_ _07571_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ net4666 rbzero.wall_tracer.rayAddendX\[1\] vssd1 vssd1 vccd1 vccd1 _02602_
+ sky130_fd_sc_hd__or2_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 _01325_ vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _09593_ _10539_ vssd1 vssd1 vccd1 vccd1 _10540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _07444_ _07805_ _07889_ _07903_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__o31a_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11965_ _05127_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03779_ clknet_0__03779_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03779_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13704_ _06851_ _06854_ _06715_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__clkbuf_4
X_17472_ _10469_ _10470_ vssd1 vssd1 vccd1 vccd1 _10471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ _07814_ _07833_ _07834_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__a21oi_2
X_11896_ _05064_ _05065_ _05004_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19211_ net5773 _03078_ _03105_ _03096_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16423_ _09493_ _09495_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_157_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _06676_ _06769_ _06770_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__or3_1
XFILLER_0_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net2041 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__04800_ clknet_0__04800_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04800_
+ sky130_fd_sc_hd__clkbuf_16
X_19142_ net6002 _03052_ _03063_ _03061_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__o211a_1
X_16354_ _09425_ _09426_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13566_ _06676_ _06687_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__xnor2_4
X_10778_ net2690 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ net3356 _08378_ _08379_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__mux2_1
X_12517_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _05218_ vssd1 vssd1 vccd1 vccd1 _05683_
+ sky130_fd_sc_hd__mux2_1
X_19073_ net6104 net2843 net2971 _03011_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__o211a_1
X_16285_ _08560_ _09216_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ _06589_ _06644_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18024_ _02072_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15236_ _08306_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12448_ net83 _05614_ net4006 vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15167_ net4334 _08144_ _08260_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _05483_ vssd1 vssd1 vccd1 vccd1 _05546_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _06881_ net531 _07268_ _06931_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19975_ rbzero.debug_overlay.facingX\[-8\] _03582_ vssd1 vssd1 vccd1 vccd1 _03584_
+ sky130_fd_sc_hd__or2_1
X_15098_ net6278 _08201_ vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14049_ _07171_ _07170_ _07169_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__a21oi_1
X_18926_ _02863_ _05391_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18857_ _05391_ _05396_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17808_ _01857_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__nand2_1
X_18788_ _02780_ _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17739_ _10597_ _01661_ _01659_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ net1689 _03212_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22420_ clknet_leaf_57_i_clk net4989 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7303 rbzero.wall_tracer.stepDistX\[-1\] vssd1 vssd1 vccd1 vccd1 net7827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7314 rbzero.wall_tracer.stepDistY\[-9\] vssd1 vssd1 vccd1 vccd1 net7838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22351_ net483 net1934 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6602 rbzero.tex_g1\[44\] vssd1 vssd1 vccd1 vccd1 net7126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6613 net2734 vssd1 vssd1 vccd1 vccd1 net7137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6624 rbzero.tex_r0\[32\] vssd1 vssd1 vccd1 vccd1 net7148 sky130_fd_sc_hd__dlygate4sd3_1
X_21302_ clknet_leaf_43_i_clk _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[5\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold6635 net2497 vssd1 vssd1 vccd1 vccd1 net7159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5901 net1372 vssd1 vssd1 vccd1 vccd1 net6425 sky130_fd_sc_hd__dlygate4sd3_1
X_22282_ net414 net2863 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
Xhold6646 _04224_ vssd1 vssd1 vccd1 vccd1 net7170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5912 rbzero.tex_r0\[14\] vssd1 vssd1 vccd1 vccd1 net6436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6657 net2602 vssd1 vssd1 vccd1 vccd1 net7181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5923 net1348 vssd1 vssd1 vccd1 vccd1 net6447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6668 rbzero.tex_r0\[50\] vssd1 vssd1 vccd1 vccd1 net7192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6679 net2169 vssd1 vssd1 vccd1 vccd1 net7203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5934 _04427_ vssd1 vssd1 vccd1 vccd1 net6458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold220 rbzero.pov.ready_buffer\[68\] vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
X_21233_ clknet_leaf_71_i_clk _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5945 net1386 vssd1 vssd1 vccd1 vccd1 net6469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5956 rbzero.tex_g1\[0\] vssd1 vssd1 vccd1 vccd1 net6480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 net5013 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5967 net1425 vssd1 vssd1 vccd1 vccd1 net6491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold242 net5027 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5978 net1478 vssd1 vssd1 vccd1 vccd1 net6502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 net5052 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 net5067 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5989 _04360_ vssd1 vssd1 vccd1 vccd1 net6513 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ _02488_ clknet_1_0__leaf__06092_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__and2_2
Xhold275 _03339_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold286 net5198 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 net5109 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
X_20115_ net4844 net4795 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21095_ net4936 net1886 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__or2_1
X_20046_ _03616_ net3176 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__or2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_104 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ net222 net2291 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ net2909 _04918_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__nand3_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ net2008 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__clkbuf_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _04843_ net4063 _04846_ _04726_ _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a221oi_1
X_13420_ _06433_ _06570_ _06569_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ net2572 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ net7582 _06160_ _06161_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__o31a_1
XFILLER_0_162_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _05464_ _05466_ _05469_ _05061_ net81 vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a221o_1
X_16070_ _09127_ _09144_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13282_ _06414_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__clkbuf_4
X_15021_ net7759 _08133_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12233_ net3241 _05374_ _05372_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1
+ vccd1 _05402_ sky130_fd_sc_hd__a22o_1
X_12164_ _04604_ net3910 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11115_ net7217 net6670 _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__mux2_1
X_12095_ rbzero.tex_r1\[11\] rbzero.tex_r1\[10\] _05263_ vssd1 vssd1 vccd1 vccd1 _05264_
+ sky130_fd_sc_hd__mux2_1
X_19760_ net6298 _03429_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__or2_1
X_16972_ _09968_ _09984_ vssd1 vssd1 vccd1 vccd1 _09986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15923_ _08989_ _08991_ _08990_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__a21o_1
X_11046_ net6878 net6618 _04392_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__mux2_1
X_18711_ net3195 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__clkbuf_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19691_ net6062 _03361_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__or2_1
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18642_ net4587 rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _02651_
+ sky130_fd_sc_hd__and2_1
X_15854_ _08869_ _08911_ _08928_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__nand3_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _07920_ _07950_ _07955_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__o21bai_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ net3838 _02586_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__or2_1
X_15785_ _08857_ _08858_ _08859_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__nand3_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12997_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__or2_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17524_ _10514_ _10522_ vssd1 vssd1 vccd1 vccd1 _10523_ sky130_fd_sc_hd__nand2_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ _07534_ _07524_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11948_ _05096_ _05116_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _06204_ _10454_ vssd1 vssd1 vccd1 vccd1 _10455_ sky130_fd_sc_hd__and2_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _07771_ _07778_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_200_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11879_ _05043_ _05045_ _05048_ _05010_ _04978_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a221o_1
X_16406_ _08584_ _09364_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ _06669_ _06693_ _06694_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__and3_1
X_17386_ _08873_ _09477_ vssd1 vssd1 vccd1 vccd1 _10386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _07747_ _07748_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19125_ net4683 _03052_ _03054_ _03048_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__o211a_1
X_16337_ net7407 _09410_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13549_ net538 _06687_ _06699_ _06692_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_153_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19056_ net5838 _03009_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__or2_1
X_16268_ _09338_ _09340_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5208 rbzero.map_overlay.i_mapdy\[5\] vssd1 vssd1 vccd1 vccd1 net5732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5219 net1593 vssd1 vssd1 vccd1 vccd1 net5743 sky130_fd_sc_hd__dlygate4sd3_1
X_18007_ _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15219_ net3507 _04818_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__nor2_2
Xhold4507 _00863_ vssd1 vssd1 vccd1 vccd1 net5031 sky130_fd_sc_hd__dlygate4sd3_1
X_16199_ _09271_ _09272_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4518 net805 vssd1 vssd1 vccd1 vccd1 net5042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4529 net777 vssd1 vssd1 vccd1 vccd1 net5053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3806 net1539 vssd1 vssd1 vccd1 vccd1 net4330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3817 net7735 vssd1 vssd1 vccd1 vccd1 net4341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3828 net7800 vssd1 vssd1 vccd1 vccd1 net4352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19958_ net3081 _03485_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__nor2_1
X_18909_ net4459 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__inv_2
X_19889_ net3921 _03511_ _03476_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__a21o_1
X_21920_ clknet_leaf_93_i_clk net1338 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_21851_ clknet_leaf_98_i_clk net4643 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20802_ clknet_1_1__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__buf_1
X_21782_ clknet_leaf_31_i_clk net3963 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20815__238 clknet_1_1__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__inv_2
XFILLER_0_92_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7100 rbzero.spi_registers.texadd3\[12\] vssd1 vssd1 vccd1 vccd1 net7624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7111 rbzero.traced_texa\[-3\] vssd1 vssd1 vccd1 vccd1 net7635 sky130_fd_sc_hd__dlygate4sd3_1
X_22403_ net155 net1042 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7122 rbzero.spi_registers.texadd2\[0\] vssd1 vssd1 vccd1 vccd1 net7646 sky130_fd_sc_hd__dlygate4sd3_1
X_20595_ net3312 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__clkbuf_1
Xhold7133 rbzero.spi_registers.texadd2\[6\] vssd1 vssd1 vccd1 vccd1 net7657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7144 rbzero.spi_registers.texadd2\[13\] vssd1 vssd1 vccd1 vccd1 net7668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6410 net2430 vssd1 vssd1 vccd1 vccd1 net6934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7155 rbzero.row_render.texu\[0\] vssd1 vssd1 vccd1 vccd1 net7679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6421 _04279_ vssd1 vssd1 vccd1 vccd1 net6945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22334_ net466 net1734 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6432 net2051 vssd1 vssd1 vccd1 vccd1 net6956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6443 _04440_ vssd1 vssd1 vccd1 vccd1 net6967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7188 net4189 vssd1 vssd1 vccd1 vccd1 net7712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6454 net2608 vssd1 vssd1 vccd1 vccd1 net6978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7199 rbzero.row_render.size\[5\] vssd1 vssd1 vccd1 vccd1 net7723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6465 _04318_ vssd1 vssd1 vccd1 vccd1 net6989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5720 rbzero.spi_registers.buf_sky\[1\] vssd1 vssd1 vccd1 vccd1 net6244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22265_ net397 net2312 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
Xhold6476 net2302 vssd1 vssd1 vccd1 vccd1 net7000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5731 rbzero.spi_registers.buf_texadd2\[9\] vssd1 vssd1 vccd1 vccd1 net6255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5742 _03949_ vssd1 vssd1 vccd1 vccd1 net6266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6487 rbzero.tex_g0\[60\] vssd1 vssd1 vccd1 vccd1 net7011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6498 net2547 vssd1 vssd1 vccd1 vccd1 net7022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5753 _00816_ vssd1 vssd1 vccd1 vccd1 net6277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21216_ clknet_leaf_75_i_clk net4734 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\]
+ sky130_fd_sc_hd__dfxtp_4
Xhold5764 rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 net6288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5775 rbzero.spi_registers.buf_texadd1\[0\] vssd1 vssd1 vccd1 vccd1 net6299 sky130_fd_sc_hd__dlygate4sd3_1
X_20709__143 clknet_1_0__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__inv_2
X_22196_ net328 net1940 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
Xhold5786 _02749_ vssd1 vssd1 vccd1 vccd1 net6310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5797 rbzero.pov.ss_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6321 sky130_fd_sc_hd__dlygate4sd3_1
X_21147_ net4030 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__clkbuf_1
X_21078_ _04069_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3_1
X_20029_ net3859 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_1
X_12920_ _04160_ _04718_ _04727_ _04777_ _06046_ _06052_ vssd1 vssd1 vccd1 vccd1 _06077_
+ sky130_fd_sc_hd__mux4_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _05207_ net29 net28 vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__and3_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _04966_ _04965_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__and2b_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _08596_ _08597_ _08613_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ net4095 _05897_ _05902_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__o22a_2
XFILLER_0_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ _06923_ _07467_ _07468_ _07090_ _07624_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__a221oi_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _04897_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20755__185 clknet_1_1__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__inv_2
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _10132_ _10134_ _10240_ vssd1 vssd1 vccd1 vccd1 _10241_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _07533_ _07599_ _07601_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nand3_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ net3853 net4052 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13403_ _06549_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__xnor2_2
X_10615_ net2263 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17171_ net3565 _09305_ vssd1 vssd1 vccd1 vccd1 _10173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14383_ _06957_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11595_ rbzero.spi_registers.texadd0\[2\] _04680_ _04765_ _04766_ _04159_ vssd1 vssd1
+ vccd1 vccd1 _04767_ sky130_fd_sc_hd__o221a_1
X_16122_ _09195_ _09196_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13334_ _06433_ _06482_ _06483_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_150_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16053_ _08493_ _09096_ _09095_ _09097_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__a2bb2o_1
X_13265_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ net7457 _08140_ _08142_ net7436 _08143_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__a221o_2
X_12216_ rbzero.debug_overlay.facingY\[-4\] _05383_ _05384_ rbzero.debug_overlay.facingY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__a22o_1
X_13196_ net2839 _06229_ _06190_ net2864 vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19812_ net6033 _03426_ net2874 _03454_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__o211a_1
X_12147_ _04790_ net4059 _05194_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__or3b_1
X_20920__333 clknet_1_0__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__inv_2
XFILLER_0_198_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19743_ net3109 _03407_ net2021 _03413_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__o211a_1
X_12078_ _05245_ _05246_ _05002_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__mux2_1
X_16955_ net4922 _09968_ vssd1 vssd1 vccd1 vccd1 _09971_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ _04243_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__clkbuf_4
X_15906_ _08949_ _08950_ _08967_ _08980_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19674_ net6588 _03375_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__or2_1
X_16886_ net4344 _09934_ _09936_ _08137_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15837_ _08898_ _08906_ _08905_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__a21o_1
X_18625_ _04633_ _02634_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15768_ _08841_ _08842_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__xnor2_1
X_18556_ _02561_ _02562_ _02563_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__o21ai_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17507_ _10385_ _10397_ _10395_ vssd1 vssd1 vccd1 vccd1 _10506_ sky130_fd_sc_hd__a21o_1
X_14719_ _07855_ _07856_ _07869_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18487_ _02495_ _02507_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15699_ _08769_ _08773_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17438_ _10253_ _10314_ _10313_ vssd1 vssd1 vccd1 vccd1 _10438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_26 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 _10205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_48 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ _10366_ _10367_ vssd1 vssd1 vccd1 vccd1 _10369_ sky130_fd_sc_hd__and2_1
XANTENNA_59 _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19108_ net5808 _03037_ _03044_ _03022_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20380_ _03791_ net3190 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5005 net1152 vssd1 vssd1 vccd1 vccd1 net5529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5016 net1294 vssd1 vssd1 vccd1 vccd1 net5540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19039_ net3941 _02988_ _03001_ _02993_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__o211a_1
Xhold5027 net1204 vssd1 vssd1 vccd1 vccd1 net5551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5038 net1123 vssd1 vssd1 vccd1 vccd1 net5562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4304 _06256_ vssd1 vssd1 vccd1 vccd1 net4828 sky130_fd_sc_hd__clkbuf_4
Xhold5049 _01037_ vssd1 vssd1 vccd1 vccd1 net5573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4315 _03757_ vssd1 vssd1 vccd1 vccd1 net4839 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22050_ clknet_leaf_90_i_clk net3368 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4326 net1282 vssd1 vssd1 vccd1 vccd1 net4850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4337 net1187 vssd1 vssd1 vccd1 vccd1 net4861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3603 net7625 vssd1 vssd1 vccd1 vccd1 net4127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4348 _00613_ vssd1 vssd1 vccd1 vccd1 net4872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3614 net681 vssd1 vssd1 vccd1 vccd1 net4138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4359 rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net4883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3625 net7634 vssd1 vssd1 vccd1 vccd1 net4149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3636 net7643 vssd1 vssd1 vccd1 vccd1 net4160 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2902 net7540 vssd1 vssd1 vccd1 vccd1 net3426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3647 _00773_ vssd1 vssd1 vccd1 vccd1 net4171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2913 _03897_ vssd1 vssd1 vccd1 vccd1 net3437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3658 net7497 vssd1 vssd1 vccd1 vccd1 net4182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2924 rbzero.pov.ready_buffer\[19\] vssd1 vssd1 vccd1 vccd1 net3448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3669 net1085 vssd1 vssd1 vccd1 vccd1 net4193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2935 _00602_ vssd1 vssd1 vccd1 vccd1 net3459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2946 net4569 vssd1 vssd1 vccd1 vccd1 net3470 sky130_fd_sc_hd__buf_1
X_20895__310 clknet_1_0__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__inv_2
Xhold2957 _02902_ vssd1 vssd1 vccd1 vccd1 net3481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2968 net4578 vssd1 vssd1 vccd1 vccd1 net3492 sky130_fd_sc_hd__buf_1
XFILLER_0_208_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2979 net4567 vssd1 vssd1 vccd1 vccd1 net3503 sky130_fd_sc_hd__buf_1
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21903_ clknet_leaf_93_i_clk net1371 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_21834_ clknet_leaf_88_i_clk net3771 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21765_ clknet_leaf_20_i_clk net1746 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21696_ clknet_leaf_2_i_clk net970 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20647_ _03977_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_101_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ net6353 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20578_ net1013 net3679 _03911_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__mux2_1
Xhold6240 net2149 vssd1 vssd1 vccd1 vccd1 net6764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6251 rbzero.tex_b1\[33\] vssd1 vssd1 vccd1 vccd1 net6775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22317_ net449 net1666 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold6262 net2328 vssd1 vssd1 vccd1 vccd1 net6786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6273 rbzero.tex_b0\[4\] vssd1 vssd1 vccd1 vccd1 net6797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6284 net2482 vssd1 vssd1 vccd1 vccd1 net6808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6295 _04187_ vssd1 vssd1 vccd1 vccd1 net6819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5550 rbzero.spi_registers.spi_buffer\[21\] vssd1 vssd1 vccd1 vccd1 net6074 sky130_fd_sc_hd__dlygate4sd3_1
X_13050_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__buf_4
Xhold5561 _02578_ vssd1 vssd1 vccd1 vccd1 net6085 sky130_fd_sc_hd__dlygate4sd3_1
X_22248_ net380 net2767 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5572 rbzero.debug_overlay.playerY\[-6\] vssd1 vssd1 vccd1 vccd1 net6096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ net4004 _05158_ _05159_ net4041 _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a221o_1
Xhold4860 _01078_ vssd1 vssd1 vccd1 vccd1 net5384 sky130_fd_sc_hd__dlygate4sd3_1
X_22179_ net311 net2667 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4871 net1066 vssd1 vssd1 vccd1 vccd1 net5395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4882 net1000 vssd1 vssd1 vccd1 vccd1 net5406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4893 net1050 vssd1 vssd1 vccd1 vccd1 net5417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ _09696_ vssd1 vssd1 vccd1 vccd1 _09810_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13952_ _07057_ _07058_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__xor2_2
XFILLER_0_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12903_ net38 net39 vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16671_ _09739_ _09741_ vssd1 vssd1 vccd1 vccd1 _09742_ sky130_fd_sc_hd__xnor2_2
X_13883_ net3408 _06898_ _06796_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_201_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15622_ _08655_ _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18410_ _02438_ _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19390_ net4194 _03198_ net1116 _03207_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _05969_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or2_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _02375_ _02378_ _01870_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a21o_1
X_15553_ _08379_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__buf_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ net3937 _05904_ _05905_ net3930 _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _07652_ _07653_ _07654_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nand3_1
X_18272_ _10259_ _10172_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__nor2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ net2802 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__inv_2
X_15484_ _08347_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__clkbuf_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12696_ net53 _05844_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ _10223_ vssd1 vssd1 vccd1 vccd1 _10224_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ _07550_ _07556_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__xnor2_1
X_11647_ net2 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_4
X_17154_ _09064_ _09364_ vssd1 vssd1 vccd1 vccd1 _10156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_4
X_14366_ _07515_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__nand2_1
Xinput46 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_4
X_11578_ _04671_ _04654_ _04669_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput57 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_4
X_16105_ _08945_ _09179_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold808 net6456 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _06466_ _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__nor2_1
X_17085_ _09669_ _09786_ _09787_ vssd1 vssd1 vccd1 vccd1 _10087_ sky130_fd_sc_hd__o21ai_4
Xhold819 net3341 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14297_ _06737_ _07366_ _07000_ _06611_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__o211a_1
X_16036_ _09102_ _09110_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__nand2_1
X_13248_ _06180_ _06182_ _06198_ _06395_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _06310_ _06313_ _06315_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a21oi_1
Xhold2209 _01540_ vssd1 vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1508 _01132_ vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_80_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17987_ _01802_ _09375_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__nor2_1
Xhold1519 net5807 vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__clkbuf_2
X_19726_ net614 _03407_ net4258 _03400_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__o211a_1
X_16938_ _06222_ _09294_ vssd1 vssd1 vccd1 vccd1 _09956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19657_ net6730 _03362_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16869_ net3993 _09925_ _09928_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18608_ net3242 net4493 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_95_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19588_ net3949 _03327_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18539_ _04623_ _09930_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21550_ clknet_leaf_3_i_clk net4250 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20501_ net3440 net1228 _03867_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__mux2_1
X_21481_ clknet_leaf_21_i_clk net2981 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20432_ _03814_ net3292 vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20927__339 clknet_1_0__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__inv_2
XFILLER_0_125_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20363_ net1587 net3268 _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4101 rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 net4625 sky130_fd_sc_hd__dlygate4sd3_1
X_22102_ net234 net2438 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4112 _01027_ vssd1 vssd1 vccd1 vccd1 net4636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4123 net846 vssd1 vssd1 vccd1 vccd1 net4647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4134 _04144_ vssd1 vssd1 vccd1 vccd1 net4658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4145 _00583_ vssd1 vssd1 vccd1 vccd1 net4669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3400 _00618_ vssd1 vssd1 vccd1 vccd1 net3924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4156 _01609_ vssd1 vssd1 vccd1 vccd1 net4680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22033_ clknet_leaf_96_i_clk net3560 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3411 _00631_ vssd1 vssd1 vccd1 vccd1 net3935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3422 _02987_ vssd1 vssd1 vccd1 vccd1 net3946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4167 _02582_ vssd1 vssd1 vccd1 vccd1 net4691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4178 _01602_ vssd1 vssd1 vccd1 vccd1 net4702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3433 net3180 vssd1 vssd1 vccd1 vccd1 net3957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3444 rbzero.spi_registers.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 net3968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4189 net7451 vssd1 vssd1 vccd1 vccd1 net4713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2710 _02406_ vssd1 vssd1 vccd1 vccd1 net3234 sky130_fd_sc_hd__buf_1
Xhold3455 _09917_ vssd1 vssd1 vccd1 vccd1 net3979 sky130_fd_sc_hd__buf_2
Xhold2721 _01014_ vssd1 vssd1 vccd1 vccd1 net3245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3466 _00474_ vssd1 vssd1 vccd1 vccd1 net3990 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_48_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2732 _03243_ vssd1 vssd1 vccd1 vccd1 net3256 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3477 net5956 vssd1 vssd1 vccd1 vccd1 net4001 sky130_fd_sc_hd__buf_2
Xhold3488 _00477_ vssd1 vssd1 vccd1 vccd1 net4012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2743 _00620_ vssd1 vssd1 vccd1 vccd1 net3267 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2754 _01223_ vssd1 vssd1 vccd1 vccd1 net3278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3499 _03964_ vssd1 vssd1 vccd1 vccd1 net4023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2765 _01229_ vssd1 vssd1 vccd1 vccd1 net3289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2776 rbzero.pov.ready_buffer\[42\] vssd1 vssd1 vccd1 vccd1 net3300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2787 _03941_ vssd1 vssd1 vccd1 vccd1 net3311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2798 rbzero.pov.ready_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net3322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ net5775 net1488 _04310_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20672__109 clknet_1_1__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__inv_2
XFILLER_0_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire81 _04977_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
X_21817_ clknet_leaf_91_i_clk net4366 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _04983_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__or2_1
X_21748_ clknet_leaf_0_i_clk net1786 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11501_ rbzero.texu_hot\[5\] _04649_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _05456_ vssd1 vssd1 vccd1 vccd1 _05647_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21679_ clknet_leaf_44_i_clk net5081 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdy\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_14220_ _07365_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ net4052 _04599_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ _07254_ _07257_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__xor2_1
X_11363_ net2431 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
X_20867__286 clknet_1_1__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__inv_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6070 net1485 vssd1 vssd1 vccd1 vccd1 net6594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _06214_ net3621 _06225_ _06257_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and4b_1
XFILLER_0_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6081 _04284_ vssd1 vssd1 vccd1 vccd1 net6605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6092 net1739 vssd1 vssd1 vccd1 vccd1 net6616 sky130_fd_sc_hd__dlygate4sd3_1
X_14082_ _07211_ _07213_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__nor2_1
X_11294_ net1907 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
Xhold5380 net2176 vssd1 vssd1 vccd1 vccd1 net5904 sky130_fd_sc_hd__dlygate4sd3_1
X_17910_ _01762_ _01852_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a21oi_1
X_13033_ _06185_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__and2_1
Xhold5391 _04210_ vssd1 vssd1 vccd1 vccd1 net5915 sky130_fd_sc_hd__dlygate4sd3_1
X_18890_ net6102 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4690 net1229 vssd1 vssd1 vccd1 vccd1 net5214 sky130_fd_sc_hd__dlygate4sd3_1
X_17841_ _01802_ _01778_ _01801_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__or3_1
X_17772_ _01799_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__xnor2_1
X_14984_ _08126_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__clkbuf_1
X_19511_ net5402 _03274_ _03281_ _03280_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__o211a_1
X_16723_ _09671_ _09688_ _09686_ vssd1 vssd1 vccd1 vccd1 _09793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13935_ _07053_ _07055_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__xor2_2
XFILLER_0_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16654_ _09719_ _09724_ vssd1 vssd1 vccd1 vccd1 _09725_ sky130_fd_sc_hd__xnor2_1
X_19442_ net5291 _03224_ _03236_ _03233_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__o211a_1
X_13866_ _06970_ _06859_ _07015_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15605_ _08652_ _08656_ _08679_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12817_ _05825_ _05957_ _05958_ net3964 vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a22o_1
X_16585_ _09535_ _09557_ _09655_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_187_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19373_ net4205 _03185_ net1407 _03194_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__o211a_1
X_13797_ _06937_ _06947_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18324_ _02363_ _02361_ _02362_ _06205_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15536_ _08320_ _08606_ _08607_ _08610_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__a31o_4
XFILLER_0_155_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ net53 _05895_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nand2_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18255_ _02181_ _02196_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15467_ _06210_ _08540_ _08541_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_182_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12679_ reg_gpout\[0\] clknet_1_0__leaf__05840_ _05204_ vssd1 vssd1 vccd1 vccd1 _05841_
+ sky130_fd_sc_hd__mux2_2
X_17206_ _10207_ net3578 net4903 vssd1 vssd1 vccd1 vccd1 _10208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418_ _07519_ _07488_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18186_ _02205_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15398_ net4288 net4358 _08434_ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__or3_4
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17137_ _08872_ _09216_ vssd1 vssd1 vccd1 vccd1 _10139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14349_ _07498_ _07497_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__or2b_1
XFILLER_0_64_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03775_ clknet_0__03775_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03775_
+ sky130_fd_sc_hd__clkbuf_16
Xhold605 _01635_ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _01312_ vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 net5526 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 net5584 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17068_ _10019_ _09769_ vssd1 vssd1 vccd1 vccd1 _10072_ sky130_fd_sc_hd__nand2_1
Xhold649 _03978_ vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
X_16019_ _08454_ _08632_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2006 net7013 vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 net7672 vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2028 _01376_ vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 net5912 vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 net6629 vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 _01285_ vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1327 net6671 vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1338 rbzero.spi_registers.buf_texadd3\[20\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1349 _00929_ vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19709_ _03294_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21602_ clknet_leaf_102_i_clk net5506 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21533_ clknet_leaf_36_i_clk net1570 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21464_ clknet_leaf_30_i_clk net3943 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20415_ net3347 net1105 _03801_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21395_ clknet_leaf_61_i_clk _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20277_ net3514 _03756_ _03767_ _03761_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3230 _03928_ vssd1 vssd1 vccd1 vccd1 net3754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3241 _03852_ vssd1 vssd1 vccd1 vccd1 net3765 sky130_fd_sc_hd__dlygate4sd3_1
X_22016_ clknet_leaf_98_i_clk net3687 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3252 _03868_ vssd1 vssd1 vccd1 vccd1 net3776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3263 _03595_ vssd1 vssd1 vccd1 vccd1 net3787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3274 _00584_ vssd1 vssd1 vccd1 vccd1 net3798 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3285 _03645_ vssd1 vssd1 vccd1 vccd1 net3809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2540 net5685 vssd1 vssd1 vccd1 vccd1 net3064 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2551 _02493_ vssd1 vssd1 vccd1 vccd1 net3075 sky130_fd_sc_hd__buf_2
Xhold3296 _01178_ vssd1 vssd1 vccd1 vccd1 net3820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2562 net4872 vssd1 vssd1 vccd1 vccd1 net3086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 _03010_ vssd1 vssd1 vccd1 vccd1 net3097 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2584 net6145 vssd1 vssd1 vccd1 vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1850 _04215_ vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2595 _00813_ vssd1 vssd1 vccd1 vccd1 net3119 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1861 net7065 vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1872 net2707 vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _04598_ _05135_ _05133_ net4041 _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__o221a_1
Xhold1883 _01569_ vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1894 net7242 vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ _06865_ _06867_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__nor2_1
X_10932_ net2831 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ _06606_ _06801_ _06621_ _06619_ _06687_ _06677_ vssd1 vssd1 vccd1 vccd1 _06802_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10863_ net6824 net2292 _04299_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20873__290 clknet_1_1__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__inv_2
X_12602_ _05035_ _05762_ _05766_ _05023_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _09333_ _09343_ _09341_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13582_ _06613_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__buf_4
X_10794_ net6936 net6704 _04266_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _08346_ _08353_ _08366_ _08373_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ reg_rgb\[22\] _05698_ _05204_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__mux2_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _02086_ _02087_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _08307_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__buf_4
X_12464_ _05069_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_91 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_91/HI o_rgb[1] sky130_fd_sc_hd__conb_1
X_14203_ _07353_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__buf_2
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ net2371 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15183_ _08270_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
X_12395_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _05483_ vssd1 vssd1 vccd1 vccd1 _05562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14134_ _07279_ _07284_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__xnor2_1
X_11346_ net2052 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
X_19991_ net3337 _03578_ net4645 _03550_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14065_ _07175_ _07215_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__nor2_1
X_18942_ _02864_ net4634 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nand2_1
X_11277_ net2437 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13016_ _06122_ _06140_ _06141_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18873_ _09943_ net4722 _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__or3_1
XFILLER_0_207_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ _01795_ _01872_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17755_ _01804_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__nand2_1
X_14967_ _07991_ _08007_ _08036_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16706_ _09773_ _09775_ _08633_ vssd1 vssd1 vccd1 vccd1 _09777_ sky130_fd_sc_hd__a21o_1
X_13918_ _07066_ _07067_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__and2b_1
X_17686_ _10340_ _10564_ _01737_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14898_ _08033_ _08045_ _08047_ vssd1 vssd1 vccd1 vccd1 _08048_ sky130_fd_sc_hd__a21o_2
XFILLER_0_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19425_ net2352 _03224_ net5862 _03220_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__o211a_1
X_16637_ _09705_ _09706_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__and2_1
X_13849_ net530 vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19356_ net5758 _03185_ _03188_ _03181_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__o211a_1
X_16568_ _09530_ _09639_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__05994_ clknet_0__05994_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__05994_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ _02346_ _02349_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15519_ _04646_ _06535_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__nand2_1
X_16499_ _08471_ _08588_ _08565_ _08516_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__o22ai_1
X_19287_ net5267 _03146_ _03149_ _03142_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18238_ _02189_ _02194_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__or2_1
Xhold6806 _03671_ vssd1 vssd1 vccd1 vccd1 net7330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6817 _03605_ vssd1 vssd1 vccd1 vccd1 net7341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6828 gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 net7352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6839 rbzero.color_sky\[2\] vssd1 vssd1 vccd1 vccd1 net7363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18169_ _02214_ _02215_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold402 net5137 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold413 net5254 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
X_20200_ net5533 _03717_ _03724_ _03722_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__o211a_1
Xhold424 net5357 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
X_21180_ net4951 net65 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold435 net5183 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 net7339 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold457 net5366 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 net5303 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
X_20131_ net3737 _03676_ _03685_ _03683_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold479 net5288 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20062_ _05393_ _03614_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _03378_ vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 rbzero.spi_registers.buf_texadd2\[19\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _03377_ vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 net6619 vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1146 net6070 vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1157 net6583 vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 net6587 vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1179 net6299 vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21516_ clknet_leaf_37_i_clk net5658 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21447_ clknet_leaf_47_i_clk net4000 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ net5870 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12180_ _04604_ net3910 _05344_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nor3_1
X_21378_ clknet_leaf_63_i_clk _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11131_ net6980 net6656 _04437_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__mux2_1
Xhold980 net4652 vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__buf_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold991 net6526 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net6940 net6449 _04404_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
Xhold3060 net5474 vssd1 vssd1 vccd1 vccd1 net3584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3071 net6116 vssd1 vssd1 vccd1 vccd1 net3595 sky130_fd_sc_hd__dlygate4sd3_1
X_15870_ _08943_ _08944_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__nor2b_4
Xhold3082 net3543 vssd1 vssd1 vccd1 vccd1 net3606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3093 _03643_ vssd1 vssd1 vccd1 vccd1 net3617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2370 _00979_ vssd1 vssd1 vccd1 vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _07638_ _07640_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__and2_1
Xhold2381 net6004 vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlymetal6s2s_1
X_20678__115 clknet_1_0__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__inv_2
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2392 net4359 vssd1 vssd1 vccd1 vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1680 _04575_ vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1691 net7009 vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _10174_ vssd1 vssd1 vccd1 vccd1 _10539_ sky130_fd_sc_hd__buf_2
X_14752_ _07887_ _07888_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__nand2_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ net2955 _05126_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03778_ clknet_0__03778_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03778_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13703_ _06800_ _06852_ _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__o21a_1
X_17471_ _10372_ _10467_ _10468_ vssd1 vssd1 vccd1 vccd1 _10470_ sky130_fd_sc_hd__and3_1
X_10915_ _04168_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14683_ _07815_ _07832_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__nor2_1
X_11895_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _05037_ vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19210_ net5247 _03079_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__or2_1
X_16422_ _09365_ _09493_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__or3_1
X_13634_ _06676_ _06776_ _06777_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and3_1
X_10846_ net7069 net7058 _04288_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16353_ _09250_ _08490_ vssd1 vssd1 vccd1 vccd1 _09426_ sky130_fd_sc_hd__and2b_1
X_19141_ net5371 _03053_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__or2_1
X_13565_ _06589_ _06715_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__nand2_2
X_10777_ net7193 net6489 _04255_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__mux2_1
X_15304_ _08304_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__buf_4
XFILLER_0_212_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _04993_ _05681_ _04999_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__o21a_1
X_19072_ net2970 _03009_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__or2_1
X_16284_ _08587_ _08582_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13496_ _06565_ _06587_ _06633_ _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15235_ _08309_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__buf_2
X_18023_ _02071_ net4599 _01749_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12447_ net4909 _04817_ _04820_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o22a_1
X_15166_ _08261_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12378_ _05261_ _05542_ _05544_ _05000_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14117_ net542 vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__inv_2
X_11329_ net2317 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19974_ net3695 _03578_ net4631 _03550_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__o211a_1
X_15097_ net3417 net3221 _08191_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14048_ _07171_ _07169_ _07170_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__and3_1
X_18925_ _02903_ _02904_ net4817 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nand3_2
XFILLER_0_197_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18856_ _05391_ _05396_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17807_ _01756_ _01757_ _01856_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18787_ net4459 rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02781_
+ sky130_fd_sc_hd__nand2_1
X_15999_ _09067_ _09073_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _01777_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ _01718_ _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19408_ net5605 _03211_ _03217_ _03207_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20680_ clknet_1_1__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__buf_1
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ net5594 _03172_ _03178_ _03168_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7304 net4361 vssd1 vssd1 vccd1 vccd1 net7828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7315 rbzero.wall_tracer.stepDistY\[-1\] vssd1 vssd1 vccd1 vccd1 net7839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22350_ net482 net1955 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6603 net2461 vssd1 vssd1 vccd1 vccd1 net7127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6614 _04583_ vssd1 vssd1 vccd1 vccd1 net7138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6625 net2641 vssd1 vssd1 vccd1 vccd1 net7149 sky130_fd_sc_hd__dlygate4sd3_1
X_21301_ clknet_leaf_41_i_clk _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22281_ net413 net2498 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
Xhold6636 rbzero.tex_r1\[54\] vssd1 vssd1 vccd1 vccd1 net7160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5902 _04478_ vssd1 vssd1 vccd1 vccd1 net6426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6647 net2729 vssd1 vssd1 vccd1 vccd1 net7171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6658 rbzero.tex_g1\[27\] vssd1 vssd1 vccd1 vccd1 net7182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5913 net1258 vssd1 vssd1 vccd1 vccd1 net6437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6669 net2689 vssd1 vssd1 vccd1 vccd1 net7193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5924 rbzero.tex_g0\[42\] vssd1 vssd1 vccd1 vccd1 net6448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5935 net1333 vssd1 vssd1 vccd1 vccd1 net6459 sky130_fd_sc_hd__dlygate4sd3_1
X_21232_ clknet_leaf_59_i_clk _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold210 _03482_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5946 _04547_ vssd1 vssd1 vccd1 vccd1 net6470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _03506_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 net5015 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5957 net1501 vssd1 vssd1 vccd1 vccd1 net6481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5968 rbzero.tex_b1\[32\] vssd1 vssd1 vccd1 vccd1 net6492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 net4606 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5979 rbzero.tex_b1\[26\] vssd1 vssd1 vccd1 vccd1 net6503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 net5054 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 net5069 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _04138_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__buf_1
Xhold276 net5122 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 net5105 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20114_ net4968 _03670_ _03673_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a21oi_1
Xhold298 net5111 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
X_21094_ _04018_ _04084_ _04086_ _04017_ net4701 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a32o_1
X_20045_ net6237 net3175 _03580_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__mux2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20980__7 clknet_1_0__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_105 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21996_ net221 net2162 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ net6359 net6852 _04214_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__mux2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ net3897 net4358 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ net7153 net7161 _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ net3262 net7582 rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _06501_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _05467_ _05468_ _05068_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13281_ _06172_ _06173_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__o21ai_1
X_22479_ clknet_leaf_67_i_clk net665 vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15020_ net7478 _08147_ vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__and2_1
X_12232_ net4772 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12163_ _04812_ net3909 vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ _04403_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__clkbuf_8
X_16971_ _09968_ _09984_ vssd1 vssd1 vccd1 vccd1 _09985_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18710_ net7146 _02713_ _02714_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ _08947_ _08993_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__xnor2_2
X_11045_ net1951 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ net4322 _03359_ net1701 _03384_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__o211a_1
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ net4587 net6237 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__nor2_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _08907_ _08912_ _08926_ _08927_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__a31o_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _07930_ _07933_ _07952_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__a21oi_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ net4476 net4446 _05403_ _02545_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__o31a_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _08449_ _08433_ _08456_ _08424_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__o22ai_2
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _06111_ _06149_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__xnor2_2
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17523_ _10519_ _10521_ vssd1 vssd1 vccd1 vccd1 _10522_ sky130_fd_sc_hd__xor2_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11947_ _05105_ net3378 _05095_ _04909_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _07858_ _07885_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__xnor2_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _10449_ _10453_ vssd1 vssd1 vccd1 vccd1 _10454_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14666_ _07816_ _07807_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__xnor2_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _05046_ _05047_ _05019_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16405_ _09086_ _09477_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__nor2_1
X_13617_ _06616_ _06688_ _06767_ _06677_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__a211o_1
X_10829_ net6712 net6403 _04277_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__mux2_1
X_17385_ _10382_ _10384_ vssd1 vssd1 vccd1 vccd1 _10385_ sky130_fd_sc_hd__xnor2_2
X_14597_ _06990_ _07359_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20732__164 clknet_1_0__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__inv_2
X_19124_ net3864 _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__or2_1
X_16336_ _09408_ _09409_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13548_ _06697_ _06698_ _06519_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16267_ _09338_ _09340_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19055_ net5838 net2843 net3097 _03011_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13479_ _06565_ _06587_ _06554_ _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__and4_1
Xhold5209 net1506 vssd1 vssd1 vccd1 vccd1 net5733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18006_ _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__nor2_1
X_15218_ net4088 _08201_ _06387_ _08239_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o211a_1
X_16198_ _09271_ _09272_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4508 net704 vssd1 vssd1 vccd1 vccd1 net5032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4519 _00726_ vssd1 vssd1 vccd1 vccd1 net5043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ net4571 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3807 net7906 vssd1 vssd1 vccd1 vccd1 net4331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3818 net2959 vssd1 vssd1 vccd1 vccd1 net4342 sky130_fd_sc_hd__buf_1
XFILLER_0_26_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3829 net3057 vssd1 vssd1 vccd1 vccd1 net4353 sky130_fd_sc_hd__buf_1
X_19957_ _03483_ _03568_ _03529_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18908_ _02863_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__inv_2
X_19888_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _02807_ _02808_ _05396_ _02787_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_175_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21850_ clknet_leaf_81_i_clk net4731 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21781_ clknet_leaf_30_i_clk _00950_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__04009_ clknet_0__04009_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04009_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22402_ net154 net2068 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
Xhold7101 rbzero.spi_registers.texadd0\[14\] vssd1 vssd1 vccd1 vccd1 net7625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7112 rbzero.spi_registers.texadd2\[19\] vssd1 vssd1 vccd1 vccd1 net7636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7123 rbzero.pov.ready_buffer\[35\] vssd1 vssd1 vccd1 vccd1 net7647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7134 rbzero.spi_registers.buf_texadd2\[20\] vssd1 vssd1 vccd1 vccd1 net7658 sky130_fd_sc_hd__dlygate4sd3_1
X_20594_ _03924_ net3311 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__and2_1
Xhold6400 net2313 vssd1 vssd1 vccd1 vccd1 net6924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7145 rbzero.spi_registers.buf_texadd2\[10\] vssd1 vssd1 vccd1 vccd1 net7669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6411 rbzero.tex_r0\[42\] vssd1 vssd1 vccd1 vccd1 net6935 sky130_fd_sc_hd__dlygate4sd3_1
X_22333_ net465 net1354 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
Xhold6422 net2446 vssd1 vssd1 vccd1 vccd1 net6946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6433 rbzero.tex_g1\[7\] vssd1 vssd1 vccd1 vccd1 net6957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_i_clk sky130_fd_sc_hd__clkbuf_8
Xhold6444 net1936 vssd1 vssd1 vccd1 vccd1 net6968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5710 rbzero.spi_registers.spi_buffer\[11\] vssd1 vssd1 vccd1 vccd1 net6234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6455 rbzero.tex_g0\[10\] vssd1 vssd1 vccd1 vccd1 net6979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22264_ net396 net2676 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
Xhold6466 net2058 vssd1 vssd1 vccd1 vccd1 net6990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5721 net1595 vssd1 vssd1 vccd1 vccd1 net6245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6477 rbzero.tex_b1\[7\] vssd1 vssd1 vccd1 vccd1 net7001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5732 net1806 vssd1 vssd1 vccd1 vccd1 net6256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6488 net2131 vssd1 vssd1 vccd1 vccd1 net7012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5743 _01252_ vssd1 vssd1 vccd1 vccd1 net6267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6499 _04375_ vssd1 vssd1 vccd1 vccd1 net7023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5754 net695 vssd1 vssd1 vccd1 vccd1 net6278 sky130_fd_sc_hd__clkbuf_2
Xhold5765 rbzero.spi_registers.buf_leak\[3\] vssd1 vssd1 vccd1 vccd1 net6289 sky130_fd_sc_hd__dlygate4sd3_1
X_21215_ clknet_leaf_74_i_clk net4949 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22195_ net327 net1958 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
Xhold5776 net1703 vssd1 vssd1 vccd1 vccd1 net6300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5787 rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 net6311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5798 net624 vssd1 vssd1 vccd1 vccd1 net6322 sky130_fd_sc_hd__dlygate4sd3_1
X_21146_ _08195_ net4029 vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__and2_1
X_21077_ _04069_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20028_ _03616_ net3858 vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12850_ net28 net29 vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net3026 _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nor2_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05916_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__or2_2
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21979_ net204 net2401 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _07622_ _07626_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__xnor2_4
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _04898_ _04599_ _04900_ _04164_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o221a_1
XFILLER_0_178_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ _07533_ _07599_ _07601_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__a21o_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11663_ net4059 net4387 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _06539_ _06550_ _06541_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a21oi_2
X_17170_ _09873_ _09738_ _09305_ vssd1 vssd1 vccd1 vccd1 _10172_ sky130_fd_sc_hd__a21o_1
X_10614_ net6902 net7026 _04170_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14382_ _06957_ _07532_ _07463_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__or3_2
XFILLER_0_187_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ rbzero.spi_registers.texadd3\[2\] _04640_ _04642_ rbzero.spi_registers.texadd2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _08411_ _08498_ vssd1 vssd1 vccd1 vccd1 _09196_ sky130_fd_sc_hd__nor2_1
X_13333_ _06140_ _06157_ net7582 vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _09089_ _09126_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ rbzero.wall_tracer.visualWallDist\[-8\] _06165_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__mux2_2
X_15003_ _06734_ _08072_ net3457 vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12215_ _05350_ _05359_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__nor2_2
X_13195_ _04868_ net3984 _06185_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19811_ net2873 _03428_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ net4001 _04831_ _04164_ _04600_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__or4_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19742_ net6784 _03408_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__or2_1
X_12077_ rbzero.tex_r1\[43\] rbzero.tex_r1\[42\] _05071_ vssd1 vssd1 vccd1 vccd1 _05246_
+ sky130_fd_sc_hd__mux2_1
X_16954_ net5969 _09966_ _09965_ _09970_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11028_ net7000 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__clkbuf_1
X_15905_ _08978_ _08979_ vssd1 vssd1 vccd1 vccd1 _08980_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19673_ net3038 _03374_ net1626 _03371_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16885_ net4611 _09934_ _09936_ net7437 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ _02621_ _02633_ _02632_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a21o_1
X_15836_ _08855_ _08856_ _08867_ _08868_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__a22o_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18555_ net4476 _02560_ _04623_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a21oi_1
X_15767_ _08367_ _08393_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__nor2_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _06130_ _06131_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__a21bo_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17506_ _10472_ _10504_ vssd1 vssd1 vccd1 vccd1 _10505_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14718_ _07858_ _07867_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__a21o_1
X_18486_ net3925 net3960 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nor2_1
X_15698_ _08770_ _08772_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__xor2_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17437_ _10375_ _10436_ vssd1 vssd1 vccd1 vccd1 _10437_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ _07797_ _07798_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__xnor2_1
XANTENNA_16 _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _10205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _10366_ _10367_ vssd1 vssd1 vccd1 vccd1 _10368_ sky130_fd_sc_hd__nor2_1
XANTENNA_49 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19107_ net5110 _03040_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__or2_1
X_16319_ _09323_ _09392_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17299_ _08755_ _09870_ vssd1 vssd1 vccd1 vccd1 _10300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5006 rbzero.pov.spi_buffer\[10\] vssd1 vssd1 vccd1 vccd1 net5530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5017 _01054_ vssd1 vssd1 vccd1 vccd1 net5541 sky130_fd_sc_hd__dlygate4sd3_1
X_19038_ net3934 _02990_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__or2_1
Xhold5028 _01041_ vssd1 vssd1 vccd1 vccd1 net5552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5039 _00822_ vssd1 vssd1 vccd1 vccd1 net5563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4305 _08245_ vssd1 vssd1 vccd1 vccd1 net4829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4316 _03764_ vssd1 vssd1 vccd1 vccd1 net4840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4327 _03760_ vssd1 vssd1 vccd1 vccd1 net4851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4338 _01109_ vssd1 vssd1 vccd1 vccd1 net4862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4349 net3086 vssd1 vssd1 vccd1 vccd1 net4873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3604 _00720_ vssd1 vssd1 vccd1 vccd1 net4128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3615 net7491 vssd1 vssd1 vccd1 vccd1 net4139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3626 _00718_ vssd1 vssd1 vccd1 vccd1 net4150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3637 _00516_ vssd1 vssd1 vccd1 vccd1 net4161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2903 rbzero.pov.ready_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net3427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3648 net1134 vssd1 vssd1 vccd1 vccd1 net4172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3659 net1010 vssd1 vssd1 vccd1 vccd1 net4183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2914 _01226_ vssd1 vssd1 vccd1 vccd1 net3438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2925 net1366 vssd1 vssd1 vccd1 vccd1 net3449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2936 net4539 vssd1 vssd1 vccd1 vccd1 net3460 sky130_fd_sc_hd__buf_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2947 net4565 vssd1 vssd1 vccd1 vccd1 net3471 sky130_fd_sc_hd__buf_1
Xhold2958 net4664 vssd1 vssd1 vccd1 vccd1 net3482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2969 net4555 vssd1 vssd1 vccd1 vccd1 net3493 sky130_fd_sc_hd__dlygate4sd3_1
X_21902_ clknet_leaf_93_i_clk net1315 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21833_ clknet_leaf_91_i_clk net4421 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21764_ clknet_leaf_25_i_clk net6174 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21695_ clknet_leaf_2_i_clk net800 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20646_ net46 _03026_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__and2_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20577_ net3672 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
Xhold6230 net2018 vssd1 vssd1 vccd1 vccd1 net6754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6241 _04468_ vssd1 vssd1 vccd1 vccd1 net6765 sky130_fd_sc_hd__dlygate4sd3_1
X_22316_ net448 net2904 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6252 net1809 vssd1 vssd1 vccd1 vccd1 net6776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6263 _04217_ vssd1 vssd1 vccd1 vccd1 net6787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6274 net1803 vssd1 vssd1 vccd1 vccd1 net6798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6285 rbzero.tex_b1\[8\] vssd1 vssd1 vccd1 vccd1 net6809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5540 _00898_ vssd1 vssd1 vccd1 vccd1 net6064 sky130_fd_sc_hd__dlygate4sd3_1
X_22247_ net379 net2526 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold6296 net2067 vssd1 vssd1 vccd1 vccd1 net6820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5551 rbzero.spi_registers.buf_texadd2\[22\] vssd1 vssd1 vccd1 vccd1 net6075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5562 net3238 vssd1 vssd1 vccd1 vccd1 net6086 sky130_fd_sc_hd__dlygate4sd3_1
X_20904__318 clknet_1_0__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__inv_2
Xhold5573 net2942 vssd1 vssd1 vccd1 vccd1 net6097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5584 _02796_ vssd1 vssd1 vccd1 vccd1 net6108 sky130_fd_sc_hd__dlygate4sd3_1
X_12000_ net2955 _04598_ _05159_ net4041 _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__o221a_1
Xhold4850 rbzero.spi_registers.buf_othery\[4\] vssd1 vssd1 vccd1 vccd1 net5374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5595 _02817_ vssd1 vssd1 vccd1 vccd1 net6119 sky130_fd_sc_hd__dlygate4sd3_1
X_22178_ net310 net1852 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold4861 net1285 vssd1 vssd1 vccd1 vccd1 net5385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4872 _00721_ vssd1 vssd1 vccd1 vccd1 net5396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4883 _00826_ vssd1 vssd1 vccd1 vccd1 net5407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4894 _00722_ vssd1 vssd1 vccd1 vccd1 net5418 sky130_fd_sc_hd__dlygate4sd3_1
X_21129_ _04114_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__nor2_1
X_13951_ _07099_ _07100_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12902_ _06048_ net36 _06054_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a31o_2
X_16670_ _09740_ _09608_ _08632_ vssd1 vssd1 vccd1 vccd1 _09741_ sky130_fd_sc_hd__a21oi_1
X_13882_ net554 _06896_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15621_ _08680_ _08694_ _08695_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ net27 _05984_ _05991_ _05944_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a22o_2
XFILLER_0_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18340_ _02375_ _02378_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__nor2_1
X_15552_ _08581_ _08626_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__nor2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _04802_ _05895_ _05903_ net4002 vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14503_ _07444_ _07400_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11715_ _04801_ _04883_ net2789 _04881_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__o221a_1
X_15483_ _08387_ _08557_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__or2_1
X_18271_ _01802_ _09863_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__nor2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _05201_ _05844_ _05852_ net73 _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_204_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17222_ _09328_ _09538_ vssd1 vssd1 vccd1 vccd1 _10223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14434_ _07546_ _07560_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__xnor2_2
X_11646_ _04802_ _04808_ _04809_ net7362 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a211oi_2
Xinput14 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_2
XFILLER_0_182_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17153_ _09103_ _09483_ vssd1 vssd1 vccd1 vccd1 _10155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14365_ _07508_ _07513_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__xor2_1
Xinput25 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_2
Xinput36 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
X_11577_ _04727_ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
X_16104_ _08938_ _08996_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__nor2_2
X_13316_ net3786 net3043 vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nor2_1
X_17084_ _10076_ net3401 _10083_ _10084_ vssd1 vssd1 vccd1 vccd1 _10086_ sky130_fd_sc_hd__o211ai_1
Xhold809 net6458 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14296_ _07416_ _07424_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16035_ _09107_ _09109_ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _06399_ _06400_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20844__265 clknet_1_0__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__inv_2
XFILLER_0_202_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13178_ _06293_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nor2_1
X_12129_ _04164_ _04637_ _04603_ _04607_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__and4_1
X_17986_ _10259_ _09602_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__nor2_1
Xhold1509 rbzero.tex_b0\[63\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
X_19725_ net4257 _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16937_ _06213_ _09295_ _09954_ vssd1 vssd1 vccd1 vccd1 _09955_ sky130_fd_sc_hd__o21ai_1
X_19656_ net1727 _03360_ net1605 _03354_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__o211a_1
XFILLER_0_204_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16868_ net3993 _09925_ _09919_ vssd1 vssd1 vccd1 vccd1 _09928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__06044_ _06044_ vssd1 vssd1 vccd1 vccd1 clknet_0__06044_ sky130_fd_sc_hd__clkbuf_16
X_18607_ _02616_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__xnor2_1
X_15819_ _08892_ _08893_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__xor2_2
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19587_ net5087 _03325_ _03328_ _03314_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__o211a_1
X_16799_ _08188_ _09737_ _08633_ vssd1 vssd1 vccd1 vccd1 _09869_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18538_ _04632_ _02547_ _02548_ net6240 _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a32o_1
XFILLER_0_181_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20348__80 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18469_ net1212 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__clkbuf_1
X_20500_ net3303 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21480_ clknet_leaf_21_i_clk net2963 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20431_ net1440 net3291 _03823_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03989_ clknet_0__03989_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03989_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20362_ _03782_ net5467 _08276_ _03477_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22101_ net233 net2106 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4102 _02799_ vssd1 vssd1 vccd1 vccd1 net4626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4113 net732 vssd1 vssd1 vccd1 vccd1 net4637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4124 rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 net4648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4135 _01637_ vssd1 vssd1 vccd1 vccd1 net4659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3401 rbzero.spi_registers.spi_cmd\[3\] vssd1 vssd1 vccd1 vccd1 net3925 sky130_fd_sc_hd__buf_1
Xhold4146 net3604 vssd1 vssd1 vccd1 vccd1 net4670 sky130_fd_sc_hd__dlygate4sd3_1
X_22032_ clknet_leaf_96_i_clk net3550 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4157 net2159 vssd1 vssd1 vccd1 vccd1 net4681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3412 net6219 vssd1 vssd1 vccd1 vccd1 net3936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4168 _02585_ vssd1 vssd1 vccd1 vccd1 net4692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3423 _00632_ vssd1 vssd1 vccd1 vccd1 net3947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4179 net1365 vssd1 vssd1 vccd1 vccd1 net4703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3434 _02996_ vssd1 vssd1 vccd1 vccd1 net3958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3445 net3374 vssd1 vssd1 vccd1 vccd1 net3969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2700 _00428_ vssd1 vssd1 vccd1 vccd1 net3224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2711 _02416_ vssd1 vssd1 vccd1 vccd1 net3235 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3456 _04127_ vssd1 vssd1 vccd1 vccd1 net3980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3467 net6312 vssd1 vssd1 vccd1 vccd1 net3991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2733 _00802_ vssd1 vssd1 vccd1 vccd1 net3257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3478 _05829_ vssd1 vssd1 vccd1 vccd1 net4002 sky130_fd_sc_hd__buf_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2744 net5570 vssd1 vssd1 vccd1 vccd1 net3268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3489 net6329 vssd1 vssd1 vccd1 vccd1 net4013 sky130_fd_sc_hd__clkbuf_2
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2755 net7256 vssd1 vssd1 vccd1 vccd1 net3279 sky130_fd_sc_hd__clkbuf_4
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20984__11 clknet_1_0__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
Xhold2766 net5602 vssd1 vssd1 vccd1 vccd1 net3290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2777 net935 vssd1 vssd1 vccd1 vccd1 net3301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2788 _03942_ vssd1 vssd1 vccd1 vccd1 net3312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2799 net1251 vssd1 vssd1 vccd1 vccd1 net3323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21816_ clknet_leaf_91_i_clk net4633 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_211_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21747_ clknet_leaf_0_i_clk net1547 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11500_ _04654_ _04669_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a21o_1
X_12480_ _05248_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21678_ clknet_leaf_27_i_clk net5188 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdy\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ _04605_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__nor2_1
X_20629_ _05816_ _03032_ _03083_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _07258_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__xnor2_2
X_11362_ net6934 net6804 _04562_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6060 net1681 vssd1 vssd1 vccd1 vccd1 net6584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _06238_ _06251_ _06255_ net4828 vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__o211a_1
Xhold6071 _04467_ vssd1 vssd1 vccd1 vccd1 net6595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6082 net1665 vssd1 vssd1 vccd1 vccd1 net6606 sky130_fd_sc_hd__dlygate4sd3_1
X_14081_ _06862_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__buf_2
X_11293_ net6692 net6506 _04529_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__mux2_1
Xhold6093 rbzero.tex_g0\[49\] vssd1 vssd1 vccd1 vccd1 net6617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5370 _04328_ vssd1 vssd1 vccd1 vccd1 net5894 sky130_fd_sc_hd__dlygate4sd3_1
X_13032_ net6186 _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__nor2_1
Xhold5381 _04480_ vssd1 vssd1 vccd1 vccd1 net5905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5392 net2557 vssd1 vssd1 vccd1 vccd1 net5916 sky130_fd_sc_hd__dlygate4sd3_1
X_17840_ _10383_ _09312_ _01783_ _01781_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4680 rbzero.pov.spi_buffer\[46\] vssd1 vssd1 vccd1 vccd1 net5204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4691 rbzero.spi_registers.buf_mapdy\[2\] vssd1 vssd1 vccd1 vccd1 net5215 sky130_fd_sc_hd__dlygate4sd3_1
X_17771_ _01820_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__nand2_1
X_14983_ net3505 _08125_ _08027_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__mux2_1
X_19510_ net614 _03275_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__or2_1
X_16722_ _09787_ _09791_ vssd1 vssd1 vccd1 vccd1 _09792_ sky130_fd_sc_hd__and2_1
X_13934_ net3405 _07081_ _07084_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19441_ net2282 _03225_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__or2_1
X_16653_ _09722_ _09723_ vssd1 vssd1 vccd1 vccd1 _09724_ sky130_fd_sc_hd__xnor2_1
X_13865_ _06970_ _06858_ _07015_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15604_ _08670_ _08677_ _08678_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__a21boi_1
X_19372_ net1784 _03186_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__or2_1
X_12816_ net25 net26 _05971_ _05973_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__a32o_1
X_16584_ _09558_ _09533_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13796_ _06920_ _06938_ net565 _06946_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_158_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18323_ _02361_ _02362_ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _08609_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _05201_ _05895_ _05903_ net73 _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__a221oi_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18254_ _02298_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15466_ net3041 _08327_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__nand2_1
X_12678_ net4045 _05788_ _05794_ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__o22a_2
XFILLER_0_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17205_ _09987_ _10085_ net7824 _10206_ vssd1 vssd1 vccd1 vccd1 _10207_ sky130_fd_sc_hd__a31o_1
X_14417_ _07565_ _07567_ _07500_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21boi_2
X_11629_ clknet_leaf_66_i_clk vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__buf_1
X_18185_ _02207_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__xor2_1
X_15397_ _08433_ _08471_ vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17136_ _09839_ _09842_ vssd1 vssd1 vccd1 vccd1 _10138_ sky130_fd_sc_hd__or2b_1
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ _07497_ _07498_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__03774_ clknet_0__03774_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03774_
+ sky130_fd_sc_hd__clkbuf_16
Xhold606 net4886 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 net5753 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold628 net5528 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_20768__196 clknet_1_1__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__inv_2
X_17067_ net3399 _10067_ _10068_ _06205_ vssd1 vssd1 vccd1 vccd1 _10071_ sky130_fd_sc_hd__a31o_1
X_14279_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__inv_2
Xhold639 net5586 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16018_ _09048_ _09092_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _04550_ vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2018 _03267_ vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 net6274 vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _03367_ vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 net6673 vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1328 _01347_ vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
X_17969_ _02016_ _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nand2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1339 _03455_ vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
X_19708_ net6740 _03395_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_100_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19639_ _02491_ _02514_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21601_ clknet_leaf_102_i_clk net4207 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21532_ clknet_leaf_36_i_clk net1530 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21463_ clknet_leaf_30_i_clk net3947 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20414_ net3455 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21394_ clknet_leaf_61_i_clk _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20276_ net3679 net4839 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3220 net7341 vssd1 vssd1 vccd1 vccd1 net3744 sky130_fd_sc_hd__dlygate4sd3_1
X_22015_ clknet_leaf_98_i_clk net3320 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3231 _01240_ vssd1 vssd1 vccd1 vccd1 net3755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3242 _03853_ vssd1 vssd1 vccd1 vccd1 net3766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3253 _03869_ vssd1 vssd1 vccd1 vccd1 net3777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3264 _03596_ vssd1 vssd1 vccd1 vccd1 net3788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2530 net4535 vssd1 vssd1 vccd1 vccd1 net3054 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3275 net5636 vssd1 vssd1 vccd1 vccd1 net3799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2541 net7828 vssd1 vssd1 vccd1 vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3286 _01023_ vssd1 vssd1 vccd1 vccd1 net3810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2552 _03251_ vssd1 vssd1 vccd1 vccd1 net3076 sky130_fd_sc_hd__clkbuf_2
Xhold3297 net6154 vssd1 vssd1 vccd1 vccd1 net3821 sky130_fd_sc_hd__buf_2
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2563 rbzero.spi_registers.spi_buffer\[13\] vssd1 vssd1 vccd1 vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2574 _00638_ vssd1 vssd1 vccd1 vccd1 net3098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1840 net7154 vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2585 net2970 vssd1 vssd1 vccd1 vccd1 net3109 sky130_fd_sc_hd__clkbuf_2
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1851 _01546_ vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2596 net7813 vssd1 vssd1 vccd1 vccd1 net3120 sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ _04602_ _05137_ _05135_ _04598_ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a221o_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1862 net7067 vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 net5845 vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 net6983 vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10931_ net7101 net7288 _04333_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__mux2_1
Xhold1895 _04254_ vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ net6533 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__clkbuf_1
X_13650_ _06616_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12601_ _05003_ _05763_ _05765_ _05061_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__o211a_1
X_13581_ _06724_ _06717_ _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__and3_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ net6774 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__clkbuf_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20327__61 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
X_15320_ _08387_ _08394_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ net83 _05697_ net4044 vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12463_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _05219_ vssd1 vssd1 vccd1 vccd1 _05629_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ _08325_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20342__75 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
X_11414_ net6920 net5924 _04584_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__mux2_1
X_14202_ _07351_ _07352_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__nand2_2
XFILLER_0_22_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_92 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_92/HI o_rgb[2] sky130_fd_sc_hd__conb_1
X_15182_ net4530 _08181_ _08260_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__mux2_1
X_12394_ _05559_ _05560_ _05248_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__mux2_1
X_14133_ _07016_ _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__xnor2_1
X_11345_ net6956 net6535 _04551_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19990_ rbzero.debug_overlay.facingX\[-2\] _03582_ vssd1 vssd1 vccd1 vccd1 _03593_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_94_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14064_ _07173_ _07174_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__and2_1
X_18941_ _02864_ net4634 vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or2_1
X_11276_ net6780 net7020 _04514_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ _06115_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18872_ net4721 _02856_ _02858_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__and3_1
XFILLER_0_207_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _09447_ _09784_ _01774_ _01772_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17754_ _08634_ _08708_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14966_ _08063_ _08064_ net7891 vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20956__366 clknet_1_0__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__inv_2
X_16705_ _09773_ _09775_ vssd1 vssd1 vccd1 vccd1 _09776_ sky130_fd_sc_hd__nor2_1
X_13917_ _07066_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__xnor2_2
X_17685_ _10562_ _10563_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nor2_1
X_14897_ net6162 vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19424_ net5861 _03225_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__or2_1
X_16636_ _09705_ _09706_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13848_ _06880_ _06953_ _06959_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19355_ net2533 _03186_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or2_1
X_16567_ _09637_ _09638_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13779_ _06837_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18306_ _02347_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15518_ _08591_ _08592_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19286_ net2076 _03147_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16498_ _08470_ _08484_ _08550_ _08565_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_47_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _02189_ _02194_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__and2_1
X_15449_ _08512_ _08522_ _08523_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6807 _03672_ vssd1 vssd1 vccd1 vccd1 net7331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6829 rbzero.trace_state\[3\] vssd1 vssd1 vccd1 vccd1 net7353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18168_ _10383_ net7378 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold403 net3439 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ _10106_ _10120_ vssd1 vssd1 vccd1 vccd1 _10121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 net5256 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold425 net3387 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18099_ _02049_ _02116_ _02145_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold436 net5374 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold447 net5266 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20130_ net3817 _03679_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__or2_1
Xhold458 net5368 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 net5370 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20061_ net4615 _03613_ _03637_ _03636_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__o211a_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _00889_ vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 net1132 vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _00888_ vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 _01379_ vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 net6072 vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 _01424_ vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _03379_ vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21515_ clknet_leaf_36_i_clk net5712 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21446_ clknet_leaf_45_i_clk net3824 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21377_ clknet_leaf_63_i_clk _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11130_ net1751 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
Xhold970 net5445 vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 net4654 vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 net6528 vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net2266 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
X_20259_ net3488 net4839 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or2_1
Xhold3050 _03883_ vssd1 vssd1 vccd1 vccd1 net3574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3061 net1125 vssd1 vssd1 vccd1 vccd1 net3585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3072 _00582_ vssd1 vssd1 vccd1 vccd1 net3596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3083 _03808_ vssd1 vssd1 vccd1 vccd1 net3607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3094 _01022_ vssd1 vssd1 vccd1 vccd1 net3618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2360 net6221 vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _07691_ _07740_ _07742_ _07968_ _07970_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__a32o_2
Xhold2371 net5998 vssd1 vssd1 vccd1 vccd1 net2895 sky130_fd_sc_hd__buf_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2382 net6006 vssd1 vssd1 vccd1 vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2393 net6013 vssd1 vssd1 vccd1 vccd1 net2917 sky130_fd_sc_hd__buf_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1670 net5851 vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__buf_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1681 _01130_ vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _07886_ _07901_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__or2_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1692 _04589_ vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11963_ _05128_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nand2_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03777_ clknet_0__03777_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03777_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06800_ _06802_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_212_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10914_ net2254 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__clkbuf_1
X_17470_ _10372_ _10467_ _10468_ vssd1 vssd1 vccd1 vccd1 _10469_ sky130_fd_sc_hd__a21oi_2
X_11894_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _05037_ vssd1 vssd1 vccd1 vccd1 _05064_
+ sky130_fd_sc_hd__mux2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _07815_ _07832_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__xor2_2
XFILLER_0_157_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _09369_ _09370_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10845_ net2560 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13633_ _06677_ _06782_ _06783_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19140_ net5918 _03052_ _03062_ _03061_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16352_ _08454_ _08795_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10776_ net2849 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__clkbuf_1
X_13564_ net7431 _06714_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__nand2_2
XFILLER_0_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15303_ _08377_ net2942 _06178_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__mux2_1
X_12515_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _05456_ vssd1 vssd1 vccd1 vccd1 _05681_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19071_ net3109 net2843 _03019_ _03011_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16283_ _09349_ _09356_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__xnor2_2
X_13495_ _06531_ _06645_ _06595_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__and3b_1
XFILLER_0_212_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18022_ net7799 _01979_ _02070_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ _08299_ _08302_ _08308_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__a21oi_2
X_12446_ _05189_ _05608_ _05610_ net4065 _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o32a_1
XFILLER_0_125_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12377_ _04993_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__or2_1
X_15165_ net4362 _08137_ _08260_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11328_ net7179 net7014 _04540_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14116_ _06957_ _06987_ _06988_ _06991_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__a2bb2o_1
X_19973_ rbzero.debug_overlay.facingX\[-9\] _03582_ vssd1 vssd1 vccd1 vccd1 _03583_
+ sky130_fd_sc_hd__or2_1
X_15096_ _08190_ net3201 net6254 _08215_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ _02903_ _02904_ net4817 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11259_ net2881 net6862 _04503_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__mux2_1
X_14047_ _07192_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18855_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _01756_ _01757_ _01856_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__nand3_1
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18786_ net4459 rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02780_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15998_ _09041_ _09071_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17737_ _01786_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__nor2_1
X_14949_ _08092_ _08094_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17668_ _10538_ _10547_ _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19407_ net2070 _03212_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__or2_1
X_16619_ _09660_ _09689_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_175_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _10358_ _10487_ _10489_ vssd1 vssd1 vccd1 vccd1 _10597_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19338_ net1909 _03173_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7316 rbzero.wall_tracer.stepDistX\[-6\] vssd1 vssd1 vccd1 vccd1 net7840 sky130_fd_sc_hd__dlygate4sd3_1
X_20306__42 clknet_1_0__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19269_ net5681 _03132_ _03138_ _03128_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6604 rbzero.tex_g1\[6\] vssd1 vssd1 vccd1 vccd1 net7128 sky130_fd_sc_hd__dlygate4sd3_1
X_21300_ clknet_leaf_43_i_clk _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.texu_hot\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6615 net2735 vssd1 vssd1 vccd1 vccd1 net7139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22280_ net412 net2454 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
Xhold6626 _04280_ vssd1 vssd1 vccd1 vccd1 net7150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6637 net2571 vssd1 vssd1 vccd1 vccd1 net7161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5903 net1373 vssd1 vssd1 vccd1 vccd1 net6427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6648 rbzero.tex_r0\[38\] vssd1 vssd1 vccd1 vccd1 net7172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5914 _04300_ vssd1 vssd1 vccd1 vccd1 net6438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6659 net2490 vssd1 vssd1 vccd1 vccd1 net7183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 net4440 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
X_21231_ clknet_leaf_71_i_clk _00400_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
X_20321__56 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
Xhold5925 net1191 vssd1 vssd1 vccd1 vccd1 net6449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 net4336 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5936 rbzero.tex_b0\[6\] vssd1 vssd1 vccd1 vccd1 net6460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5947 net1387 vssd1 vssd1 vccd1 vccd1 net6471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 net6156 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5958 _04385_ vssd1 vssd1 vccd1 vccd1 net6482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 net7492 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 net4608 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5969 net1397 vssd1 vssd1 vccd1 vccd1 net6493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 net4982 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ _02488_ clknet_1_0__leaf__06044_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__and2_2
XFILLER_0_141_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 net5090 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 net5131 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
X_20113_ net4968 _03670_ _03661_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21ai_1
Xhold288 net5107 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 rbzero.spi_registers.buf_mapdx\[3\] vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
X_21093_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20044_ net3840 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939__350 clknet_1_1__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__inv_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ net220 net2615 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ clknet_1_0__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__buf_1
XFILLER_0_139_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _04169_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12300_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _05218_ vssd1 vssd1 vccd1 vccd1 _05468_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__buf_2
XFILLER_0_162_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22478_ clknet_leaf_77_i_clk net1184 vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ net4708 _05371_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__a21oi_1
X_21429_ clknet_leaf_43_i_clk net3036 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20684__120 clknet_1_0__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__inv_2
XFILLER_0_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12162_ net3908 _04811_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ net2718 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12093_ _05070_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__clkbuf_8
X_16970_ net5420 _09983_ vssd1 vssd1 vccd1 vccd1 _09984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15921_ _08994_ _08995_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__and2_1
X_11044_ net6932 net6878 _04392_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _02645_ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _08913_ _08925_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__and2b_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 net7299 vssd1 vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _07920_ _07950_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ net4691 _02581_ _02580_ _02574_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a211o_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _08444_ _08493_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__nor2_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _06147_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__xnor2_2
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _10520_ _09477_ _10387_ _10390_ vssd1 vssd1 vccd1 vccd1 _10521_ sky130_fd_sc_hd__o31a_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _07868_ _07867_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__and2b_1
X_11946_ _05107_ _05114_ _05115_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__mux2_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _10204_ _10451_ _10452_ vssd1 vssd1 vccd1 vccd1 _10453_ sky130_fd_sc_hd__o21a_4
XFILLER_0_188_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14665_ _07808_ _07803_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__nand2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _04988_ vssd1 vssd1 vccd1 vccd1 _05047_
+ sky130_fd_sc_hd__mux2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16404_ _09222_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _06697_ _06698_ _06614_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10828_ net2852 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__clkbuf_1
X_17384_ _10383_ _08708_ vssd1 vssd1 vccd1 vccd1 _10384_ sky130_fd_sc_hd__nor2_1
X_14596_ _07746_ _07744_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19123_ _03039_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__buf_2
XFILLER_0_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16335_ _09278_ _09292_ _09407_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__and3_1
X_13547_ _06694_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__buf_4
X_10759_ net1473 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__clkbuf_1
X_19054_ _02992_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__clkbuf_4
X_16266_ _09195_ _09196_ _09339_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _06612_ _06552_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nor2_1
X_18005_ _01935_ _01947_ _01945_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15217_ net4087 vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__buf_4
X_12429_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _04994_ vssd1 vssd1 vccd1 vccd1 _05596_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16197_ _08943_ _08836_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4509 rbzero.spi_registers.buf_texadd0\[21\] vssd1 vssd1 vccd1 vccd1 net5033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15148_ net4570 _08059_ _08249_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3808 net3042 vssd1 vssd1 vccd1 vccd1 net4332 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3819 net3551 vssd1 vssd1 vccd1 vccd1 net4343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15079_ rbzero.wall_tracer.visualWallDist\[-8\] _08201_ vssd1 vssd1 vccd1 vccd1 _08204_
+ sky130_fd_sc_hd__or2_1
X_19956_ net3279 _03564_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18907_ net4662 _02883_ _02890_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__nand3_1
X_19887_ net3921 _03511_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__or2_1
X_18838_ net1580 _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18769_ net4438 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21780_ clknet_leaf_30_i_clk net3154 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__04008_ clknet_0__04008_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04008_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22401_ net153 net2471 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7113 rbzero.traced_texa\[5\] vssd1 vssd1 vccd1 vccd1 net7637 sky130_fd_sc_hd__dlygate4sd3_1
X_20593_ net3310 net1508 net3250 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__mux2_1
Xhold7124 rbzero.traced_texa\[4\] vssd1 vssd1 vccd1 vccd1 net7648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7135 rbzero.spi_registers.buf_texadd3\[10\] vssd1 vssd1 vccd1 vccd1 net7659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6401 rbzero.tex_b1\[20\] vssd1 vssd1 vccd1 vccd1 net6925 sky130_fd_sc_hd__dlygate4sd3_1
X_22332_ net464 net2306 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
Xhold7146 rbzero.row_render.texu\[3\] vssd1 vssd1 vccd1 vccd1 net7670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6412 net2421 vssd1 vssd1 vccd1 vccd1 net6936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6423 rbzero.tex_b0\[23\] vssd1 vssd1 vccd1 vccd1 net6947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6434 net2514 vssd1 vssd1 vccd1 vccd1 net6958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6445 rbzero.tex_b0\[18\] vssd1 vssd1 vccd1 vccd1 net6969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5700 rbzero.spi_registers.spi_buffer\[5\] vssd1 vssd1 vccd1 vccd1 net6224 sky130_fd_sc_hd__dlygate4sd3_1
X_22263_ net395 net1063 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
Xhold6456 net2116 vssd1 vssd1 vccd1 vccd1 net6980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5711 rbzero.spi_registers.buf_texadd2\[5\] vssd1 vssd1 vccd1 vccd1 net6235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6467 rbzero.tex_r0\[11\] vssd1 vssd1 vccd1 vccd1 net6991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5722 _03244_ vssd1 vssd1 vccd1 vccd1 net6246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5733 rbzero.spi_registers.buf_texadd1\[5\] vssd1 vssd1 vccd1 vccd1 net6257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6478 net2653 vssd1 vssd1 vccd1 vccd1 net7002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6489 rbzero.tex_b0\[43\] vssd1 vssd1 vccd1 vccd1 net7013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5744 rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 net6268 sky130_fd_sc_hd__dlygate4sd3_1
X_21214_ _03502_ net1048 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__nor2_1
Xhold5755 _08217_ vssd1 vssd1 vccd1 vccd1 net6279 sky130_fd_sc_hd__dlygate4sd3_1
X_22194_ net326 net2026 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
Xhold5766 net1735 vssd1 vssd1 vccd1 vccd1 net6290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5777 rbzero.spi_registers.buf_floor\[0\] vssd1 vssd1 vccd1 vccd1 net6301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5788 gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 net6312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5799 rbzero.pov.sclk_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6323 sky130_fd_sc_hd__dlygate4sd3_1
X_21145_ net4028 net4027 net3981 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux2_1
Xwire1 _02826_ vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__buf_1
XFILLER_0_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21076_ _04064_ _04067_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__nand2_1
X_20027_ net3857 net3764 _03594_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11800_ _04912_ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__xnor2_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ net21 _05931_ _05939_ _05893_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a22o_2
X_21978_ net203 net2583 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer70 _06846_ vssd1 vssd1 vccd1 vccd1 net3370 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ net4345 _04600_ _04606_ net2774 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__o22a_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20716__149 clknet_1_1__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__inv_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14450_ _07531_ _07600_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__or2_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _04831_ net3917 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _06547_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__xor2_4
XFILLER_0_187_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10613_ net2648 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14381_ _06955_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__buf_2
X_11593_ rbzero.spi_registers.texadd1\[2\] _04644_ _04709_ vssd1 vssd1 vccd1 vccd1
+ _04765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16120_ _09193_ _09194_ vssd1 vssd1 vccd1 vccd1 _09195_ sky130_fd_sc_hd__xnor2_1
X_13332_ net6281 _06430_ _06414_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__o21a_1
X_16051_ _09100_ _09099_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13263_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _08093_ _08111_ _08128_ _08141_ _08069_ net7759 vssd1 vssd1 vccd1 vccd1 _08142_
+ sky130_fd_sc_hd__mux4_2
X_12214_ _05367_ _05359_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__nor2_2
XFILLER_0_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6990 net4233 vssd1 vssd1 vccd1 vccd1 net7514 sky130_fd_sc_hd__dlygate4sd3_1
X_13194_ net2925 vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__inv_2
X_19810_ net6047 _03426_ net2283 _03454_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__o211a_1
X_12145_ _05310_ _05312_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ rbzero.tex_r1\[41\] rbzero.tex_r1\[40\] _05071_ vssd1 vssd1 vccd1 vccd1 _05245_
+ sky130_fd_sc_hd__mux2_1
X_19741_ net6029 _03407_ net1645 _03413_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__o211a_1
X_16953_ _09967_ _09969_ vssd1 vssd1 vccd1 vccd1 _09970_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ net6998 net2439 _04310_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15904_ _08951_ _08966_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__xor2_1
X_19672_ net6562 _03375_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16884_ net4284 _09934_ _09936_ _08125_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18623_ _02613_ _02619_ _02607_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__o21ai_1
X_15835_ _08871_ _08883_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__xnor2_2
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18554_ net4476 net4446 _05403_ net4424 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__or4_1
X_15766_ _08347_ _08373_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__or2_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12978_ _06132_ _06094_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__or2b_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _10502_ _10503_ vssd1 vssd1 vccd1 vccd1 _10504_ sky130_fd_sc_hd__nand2_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ _07859_ _07860_ _07866_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__and3_1
XFILLER_0_185_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11929_ net4303 net4271 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nand2_1
X_18485_ net3889 _02505_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15697_ _08686_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__nand2_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ _10433_ _10435_ vssd1 vssd1 vccd1 vccd1 _10436_ sky130_fd_sc_hd__xor2_2
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14648_ _07797_ _07798_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17367_ _10235_ _10243_ _10241_ vssd1 vssd1 vccd1 vccd1 _10367_ sky130_fd_sc_hd__a21oi_1
XANTENNA_39 _10329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ _07676_ _07722_ _07725_ _07727_ _07729_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_67_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19106_ net6014 _03037_ _03043_ _03022_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__o211a_1
X_16318_ _09389_ _09391_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17298_ _09096_ _10168_ vssd1 vssd1 vccd1 vccd1 _10299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19037_ net3940 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__buf_4
Xhold5007 _01046_ vssd1 vssd1 vccd1 vccd1 net5531 sky130_fd_sc_hd__dlygate4sd3_1
X_16249_ _09259_ _09322_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5018 net1295 vssd1 vssd1 vccd1 vccd1 net5542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5029 rbzero.pov.spi_buffer\[11\] vssd1 vssd1 vccd1 vccd1 net5553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4306 _00434_ vssd1 vssd1 vccd1 vccd1 net4830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4317 _01101_ vssd1 vssd1 vccd1 vccd1 net4841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4328 _01098_ vssd1 vssd1 vccd1 vccd1 net4852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4339 net1188 vssd1 vssd1 vccd1 vccd1 net4863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3605 net608 vssd1 vssd1 vccd1 vccd1 net4129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3616 net757 vssd1 vssd1 vccd1 vccd1 net4140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3627 net611 vssd1 vssd1 vccd1 vccd1 net4151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3638 net672 vssd1 vssd1 vccd1 vccd1 net4162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2904 net740 vssd1 vssd1 vccd1 vccd1 net3428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3649 net7641 vssd1 vssd1 vccd1 vccd1 net4173 sky130_fd_sc_hd__buf_1
Xhold2915 rbzero.pov.ready_buffer\[43\] vssd1 vssd1 vccd1 vccd1 net3439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2926 _03826_ vssd1 vssd1 vccd1 vccd1 net3450 sky130_fd_sc_hd__dlygate4sd3_1
X_19939_ _03553_ _03554_ _03476_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2937 net4925 vssd1 vssd1 vccd1 vccd1 net3461 sky130_fd_sc_hd__dlygate4sd3_1
X_20821__244 clknet_1_0__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__inv_2
Xhold2948 net4557 vssd1 vssd1 vccd1 vccd1 net3472 sky130_fd_sc_hd__buf_1
Xhold2959 rbzero.pov.ready_buffer\[58\] vssd1 vssd1 vccd1 vccd1 net3483 sky130_fd_sc_hd__buf_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21901_ clknet_leaf_94_i_clk net1511 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21832_ clknet_leaf_96_i_clk net4415 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21763_ clknet_leaf_25_i_clk net6166 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21694_ clknet_leaf_3_i_clk net5032 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20645_ net3937 _03974_ _03976_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ _03924_ net3671 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6220 net1759 vssd1 vssd1 vccd1 vccd1 net6744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6231 rbzero.tex_g0\[4\] vssd1 vssd1 vccd1 vccd1 net6755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6242 net2150 vssd1 vssd1 vccd1 vccd1 net6766 sky130_fd_sc_hd__dlygate4sd3_1
X_22315_ net447 net2853 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold6253 rbzero.tex_g1\[4\] vssd1 vssd1 vccd1 vccd1 net6777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6264 net2329 vssd1 vssd1 vccd1 vccd1 net6788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6275 _04593_ vssd1 vssd1 vccd1 vccd1 net6799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5530 rbzero.spi_registers.buf_texadd2\[21\] vssd1 vssd1 vccd1 vccd1 net6054 sky130_fd_sc_hd__dlygate4sd3_1
X_22246_ net378 net2640 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold6286 net2605 vssd1 vssd1 vccd1 vccd1 net6810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5541 rbzero.spi_registers.buf_texadd2\[17\] vssd1 vssd1 vccd1 vccd1 net6065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5552 net2354 vssd1 vssd1 vccd1 vccd1 net6076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6297 rbzero.tex_b0\[31\] vssd1 vssd1 vccd1 vccd1 net6821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5574 net3222 vssd1 vssd1 vccd1 vccd1 net6098 sky130_fd_sc_hd__clkbuf_4
Xhold5585 net3458 vssd1 vssd1 vccd1 vccd1 net6109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4840 net1052 vssd1 vssd1 vccd1 vccd1 net5364 sky130_fd_sc_hd__dlygate4sd3_1
X_22177_ net309 net1937 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold5596 net3726 vssd1 vssd1 vccd1 vccd1 net6120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4851 net960 vssd1 vssd1 vccd1 vccd1 net5375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4862 rbzero.pov.spi_buffer\[41\] vssd1 vssd1 vccd1 vccd1 net5386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4873 rbzero.spi_registers.texadd3\[2\] vssd1 vssd1 vccd1 vccd1 net5397 sky130_fd_sc_hd__dlygate4sd3_1
X_21128_ net4133 net4740 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__and2_1
Xhold4884 net1001 vssd1 vssd1 vccd1 vccd1 net5408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4895 rbzero.wall_tracer.mapX\[10\] vssd1 vssd1 vccd1 vccd1 net5419 sky130_fd_sc_hd__dlygate4sd3_1
X_13950_ _07098_ _07086_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__and2b_1
X_21059_ _04053_ _04056_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__xnor2_1
X_20796__221 clknet_1_1__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__inv_2
X_12901_ _06055_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__o21ba_2
X_13881_ _06864_ _06966_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__nor2_2
XFILLER_0_193_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15620_ _08652_ _08656_ _08679_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__or3_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12832_ _05986_ _05987_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a21o_2
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15551_ _08625_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__clkbuf_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _05825_ _05904_ _05905_ net3965 vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14502_ _07438_ _07532_ net586 _07466_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _01812_ _01711_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__nor2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ net4033 net2879 vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__xnor2_1
X_15482_ net3171 _08312_ _08556_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__a21boi_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ net52 _05853_ _05854_ net51 vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17221_ _10148_ _10127_ vssd1 vssd1 vccd1 vccd1 _10222_ sky130_fd_sc_hd__or2b_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _07583_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ net4004 _04814_ net3992 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17152_ _09862_ _09867_ _10153_ vssd1 vssd1 vccd1 vccd1 _10154_ sky130_fd_sc_hd__a21bo_1
Xinput15 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_2
X_14364_ _07514_ _07487_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__xnor2_1
X_11576_ _04714_ _04678_ _04745_ _04747_ _04160_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o311a_1
Xinput26 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_2
Xinput37 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_4
X_16103_ _09174_ _09177_ _08995_ _09175_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__a2bb2o_2
Xinput48 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
X_13315_ net3786 net3043 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17083_ _10083_ _10084_ _10076_ net3401 vssd1 vssd1 vccd1 vccd1 _10085_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295_ _07428_ _07430_ _07426_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _09108_ _08874_ _09106_ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13246_ net4887 _06396_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13177_ _06288_ _06289_ _06332_ _06278_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12128_ _04892_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__inv_2
X_17985_ _01942_ _01936_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__or2b_1
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12059_ _05002_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__or2_1
X_19724_ _03394_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__buf_2
X_16936_ _09952_ _09953_ vssd1 vssd1 vccd1 vccd1 _09954_ sky130_fd_sc_hd__nand2_1
X_19655_ net6258 _03362_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__or2_1
X_16867_ net4056 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15818_ _08367_ _08410_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__nor2_1
X_18606_ net4667 _02606_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19586_ net1571 _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or2_1
X_16798_ _09862_ _09867_ vssd1 vssd1 vccd1 vccd1 _09868_ sky130_fd_sc_hd__xor2_1
X_18537_ _02549_ net6239 _08246_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15749_ _08459_ _08447_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ net7205 _02488_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17419_ _09138_ _09139_ _10168_ _10174_ vssd1 vssd1 vccd1 vccd1 _10419_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18399_ _02430_ net4487 _02411_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20430_ net3354 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03988_ clknet_0__03988_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03988_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20361_ net6176 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__buf_4
XFILLER_0_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22100_ net232 net1876 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4103 _02802_ vssd1 vssd1 vccd1 vccd1 net4627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4114 net7797 vssd1 vssd1 vccd1 vccd1 net4638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4125 net2776 vssd1 vssd1 vccd1 vccd1 net4649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4136 net716 vssd1 vssd1 vccd1 vccd1 net4660 sky130_fd_sc_hd__dlygate4sd3_1
X_22031_ clknet_leaf_96_i_clk net3846 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3402 _03466_ vssd1 vssd1 vccd1 vccd1 net3926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4147 rbzero.spi_registers.buf_texadd1\[20\] vssd1 vssd1 vccd1 vccd1 net4671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3413 _05828_ vssd1 vssd1 vccd1 vccd1 net3937 sky130_fd_sc_hd__buf_4
XFILLER_0_12_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4158 rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 net4682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3424 rbzero.spi_registers.spi_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net3948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4169 _00581_ vssd1 vssd1 vccd1 vccd1 net4693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3435 _00630_ vssd1 vssd1 vccd1 vccd1 net3959 sky130_fd_sc_hd__dlygate4sd3_1
X_20291__28 clknet_1_1__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
Xhold3446 _02519_ vssd1 vssd1 vccd1 vccd1 net3970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2701 rbzero.pov.spi_counter\[0\] vssd1 vssd1 vccd1 vccd1 net3225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 _02422_ vssd1 vssd1 vccd1 vccd1 net3236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3457 _04128_ vssd1 vssd1 vccd1 vccd1 net3981 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2723 net6088 vssd1 vssd1 vccd1 vccd1 net3247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3468 net3975 vssd1 vssd1 vccd1 vccd1 net3992 sky130_fd_sc_hd__clkbuf_4
Xhold2734 rbzero.pov.ready_buffer\[61\] vssd1 vssd1 vccd1 vccd1 net3258 sky130_fd_sc_hd__buf_1
Xhold3479 _01261_ vssd1 vssd1 vccd1 vccd1 net4003 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2745 _03783_ vssd1 vssd1 vccd1 vccd1 net3269 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2756 _02744_ vssd1 vssd1 vccd1 vccd1 net3280 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2767 net1272 vssd1 vssd1 vccd1 vccd1 net3291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2778 _03876_ vssd1 vssd1 vccd1 vccd1 net3302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2789 _01247_ vssd1 vssd1 vccd1 vccd1 net3313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21815_ clknet_leaf_9_i_clk net3955 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21746_ clknet_leaf_0_i_clk net1565 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21677_ clknet_leaf_16_i_clk net5016 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdy\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ net3908 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__inv_2
XFILLER_0_191_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20628_ _05299_ net3898 _03965_ _08276_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11361_ net6834 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20559_ net3258 net1282 _03911_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6050 net1641 vssd1 vssd1 vccd1 vccd1 net6574 sky130_fd_sc_hd__dlygate4sd3_1
X_13100_ net7770 vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__inv_2
Xhold6061 rbzero.spi_registers.buf_texadd1\[11\] vssd1 vssd1 vccd1 vccd1 net6585 sky130_fd_sc_hd__dlygate4sd3_1
X_11292_ net2416 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
Xhold6072 net1486 vssd1 vssd1 vccd1 vccd1 net6596 sky130_fd_sc_hd__dlygate4sd3_1
X_14080_ _07189_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6083 rbzero.spi_registers.buf_texadd1\[3\] vssd1 vssd1 vccd1 vccd1 net6607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6094 net1658 vssd1 vssd1 vccd1 vccd1 net6618 sky130_fd_sc_hd__dlygate4sd3_1
X_20657__96 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__inv_2
Xhold5360 _00704_ vssd1 vssd1 vccd1 vccd1 net5884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5371 net2633 vssd1 vssd1 vccd1 vccd1 net5895 sky130_fd_sc_hd__dlygate4sd3_1
X_13031_ _06186_ _06178_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nor2_1
X_22229_ net361 net1981 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold5382 net2177 vssd1 vssd1 vccd1 vccd1 net5906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5393 rbzero.map_overlay.i_mapdy\[0\] vssd1 vssd1 vccd1 vccd1 net5917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4670 _01080_ vssd1 vssd1 vccd1 vccd1 net5194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4681 net1375 vssd1 vssd1 vccd1 vccd1 net5205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4692 net841 vssd1 vssd1 vccd1 vccd1 net5216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17770_ _01706_ _01800_ _01819_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__nand3_1
Xhold3980 _01600_ vssd1 vssd1 vccd1 vccd1 net4504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3991 _03601_ vssd1 vssd1 vccd1 vccd1 net4515 sky130_fd_sc_hd__dlygate4sd3_1
X_14982_ net7439 _08124_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16721_ _09788_ _09789_ net7378 _08326_ vssd1 vssd1 vccd1 vccd1 _09791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13933_ _06862_ _06867_ _07082_ _07083_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19440_ net4979 _03224_ _03235_ _03233_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__o211a_1
X_16652_ _08684_ _08582_ vssd1 vssd1 vccd1 vccd1 _09723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13864_ _06876_ _06867_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15603_ _08657_ _08659_ _08669_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__nand3_1
X_19371_ net4208 _03185_ net1215 _03194_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__o211a_1
X_12815_ _04760_ _04603_ _04637_ _04165_ net22 net23 vssd1 vssd1 vccd1 vccd1 _05974_
+ sky130_fd_sc_hd__mux4_1
X_16583_ _09531_ _09635_ _09634_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__a21o_2
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13795_ _06891_ _06943_ _06944_ _06945_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18322_ _02353_ _02354_ _02355_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__o21ai_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _08319_ _08608_ _08297_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__o21a_4
XFILLER_0_167_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12746_ net52 _05904_ _05905_ net51 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _09231_ _09310_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__or2_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15465_ net3210 _08305_ _08536_ _08539_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__a22o_4
X_20850__270 clknet_1_1__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__inv_2
X_12677_ _05784_ _05804_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a21o_2
XFILLER_0_155_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17204_ _06204_ _10205_ vssd1 vssd1 vccd1 vccd1 _10206_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14416_ _07502_ _07566_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__nand2_2
X_18184_ _02216_ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11628_ _04799_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_2
X_15396_ _08470_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__buf_2
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17135_ _09840_ _09841_ vssd1 vssd1 vccd1 vccd1 _10137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _07082_ _07467_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03773_ clknet_0__03773_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03773_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11559_ _04691_ _04694_ _04695_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a21o_1
Xhold607 net4888 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _03076_ vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold629 net6406 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ _10067_ _10068_ net3399 vssd1 vssd1 vccd1 vccd1 _10070_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14278_ _07374_ _07383_ _07381_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _09091_ _08664_ _09020_ _09050_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13229_ _06203_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__or2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _01152_ vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 net6272 vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _00881_ vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 net6675 vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17968_ _01932_ _01988_ _02015_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__nand3_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1329 net6687 vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
X_19707_ _02996_ _03393_ net1788 _03384_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__o211a_1
X_16919_ net4176 _09941_ _09942_ net6146 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899_ _01823_ _01843_ _01841_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a21oi_1
X_19638_ net5038 net798 _03356_ _03354_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19569_ net3093 _03304_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20933__345 clknet_1_1__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__inv_2
XFILLER_0_193_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21600_ clknet_leaf_102_i_clk net4210 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21531_ clknet_leaf_36_i_clk net1651 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21462_ clknet_leaf_30_i_clk net3935 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20413_ _03814_ net3454 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21393_ clknet_leaf_60_i_clk _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20344_ clknet_1_1__leaf__03773_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__buf_1
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20275_ net3679 _03756_ _03766_ _03761_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3210 _03923_ vssd1 vssd1 vccd1 vccd1 net3734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22014_ clknet_leaf_97_i_clk net3588 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3221 _03606_ vssd1 vssd1 vccd1 vccd1 net3745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3232 rbzero.pov.ready_buffer\[22\] vssd1 vssd1 vccd1 vccd1 net3756 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3243 _01206_ vssd1 vssd1 vccd1 vccd1 net3767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3254 _01213_ vssd1 vssd1 vccd1 vccd1 net3778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2520 _02701_ vssd1 vssd1 vccd1 vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3265 _00993_ vssd1 vssd1 vccd1 vccd1 net3789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3276 net1306 vssd1 vssd1 vccd1 vccd1 net3800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2531 _08225_ vssd1 vssd1 vccd1 vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2542 net4928 vssd1 vssd1 vccd1 vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3287 net4847 vssd1 vssd1 vccd1 vccd1 net3811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2553 _03252_ vssd1 vssd1 vccd1 vccd1 net3077 sky130_fd_sc_hd__buf_2
Xhold3298 _02945_ vssd1 vssd1 vccd1 vccd1 net3822 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 net697 vssd1 vssd1 vccd1 vccd1 net3088 sky130_fd_sc_hd__clkbuf_4
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2575 rbzero.spi_registers.spi_buffer\[15\] vssd1 vssd1 vccd1 vccd1 net3099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 net6075 vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1841 _01575_ vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2586 _00646_ vssd1 vssd1 vccd1 vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1852 net6865 vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 _04618_ vssd1 vssd1 vccd1 vccd1 net3121 sky130_fd_sc_hd__clkbuf_1
Xhold1863 _01463_ vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1874 _01440_ vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ net6754 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__clkbuf_1
Xhold1885 _04590_ vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1896 _01513_ vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10861_ net6531 net2107 _04299_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ _05068_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__or2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13580_ _06421_ _06695_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ net6772 net2421 _04266_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _05189_ _05692_ _05695_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__o211a_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21729_ clknet_leaf_21_i_clk net1714 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _08299_ _08323_ _08324_ _08312_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__a211o_2
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ _05062_ _05623_ _05625_ _05627_ _04979_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ _07307_ _07350_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__nand2_1
X_11413_ net6800 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _08269_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_93 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_93/HI o_rgb[3] sky130_fd_sc_hd__conb_1
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12393_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _05456_ vssd1 vssd1 vccd1 vccd1 _05560_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14132_ _07281_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__and2_1
X_11344_ net6748 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14063_ _07211_ _07213_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__and2_1
X_18940_ _02903_ _02909_ _02921_ _08246_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a31o_1
X_11275_ net6339 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
Xhold5190 net1585 vssd1 vssd1 vccd1 vccd1 net5714 sky130_fd_sc_hd__dlygate4sd3_1
X_13014_ _06095_ _06104_ _06108_ _06105_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18871_ net4721 _02856_ _02858_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a21oi_1
X_17822_ _01797_ _01763_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17753_ _01801_ _01803_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__xnor2_1
X_14965_ _08006_ _08061_ _06664_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__a21o_1
X_16704_ net7407 _09774_ vssd1 vssd1 vccd1 vccd1 _09775_ sky130_fd_sc_hd__xnor2_1
X_13916_ _06981_ _06983_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__xor2_2
XFILLER_0_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17684_ _10469_ _01735_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ _06626_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__clkbuf_1
X_16635_ _08564_ _08717_ _09572_ _09570_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__o31a_1
X_19423_ net5578 _03224_ _03226_ _03220_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _06956_ _06958_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _09414_ _09512_ _09510_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__a21oi_4
X_19354_ net5736 _03185_ _03187_ _03181_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__o211a_1
X_13778_ _06826_ _06888_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__xor2_2
XFILLER_0_58_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18305_ net4687 net4455 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__nand2_1
X_15517_ _08152_ _08575_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12729_ _05865_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__or2_2
X_19285_ net5306 _03146_ _03148_ _03142_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__o211a_1
X_16497_ _09567_ _09568_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _02181_ _02281_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15448_ _08513_ _08521_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6819 _03599_ vssd1 vssd1 vccd1 vccd1 net7343 sky130_fd_sc_hd__dlygate4sd3_1
X_18167_ _02212_ _02213_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ _08298_ _08452_ _08453_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17118_ _10118_ _10119_ vssd1 vssd1 vccd1 vccd1 _10120_ sky130_fd_sc_hd__nor2_1
Xhold404 net4408 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18098_ _02049_ _02116_ _02145_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a21oi_1
Xhold415 net5317 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 net4495 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 net5376 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold448 net5268 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ _10019_ _09521_ vssd1 vssd1 vccd1 vccd1 _10055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold459 net5290 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20060_ net4438 _03614_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 net6563 vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _03419_ vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 net5772 vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__buf_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1137 net6232 vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1148 net6073 vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 net6879 vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21514_ clknet_leaf_36_i_clk net4199 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21445_ clknet_leaf_86_i_clk net3020 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21376_ clknet_leaf_63_i_clk _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 net4848 vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 net7754 vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net7095 net6940 _04404_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__mux2_1
Xhold982 net5732 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__buf_1
Xhold993 _01406_ vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
X_20258_ net4838 vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__buf_1
Xhold3040 _01034_ vssd1 vssd1 vccd1 vccd1 net3564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3051 _03884_ vssd1 vssd1 vccd1 vccd1 net3575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3062 _03802_ vssd1 vssd1 vccd1 vccd1 net3586 sky130_fd_sc_hd__dlygate4sd3_1
X_20189_ _03678_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__clkbuf_2
Xhold3073 net5766 vssd1 vssd1 vccd1 vccd1 net3597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3084 _03809_ vssd1 vssd1 vccd1 vccd1 net3608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2350 _03458_ vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3095 net5698 vssd1 vssd1 vccd1 vccd1 net3619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2361 net6223 vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2372 net6000 vssd1 vssd1 vccd1 vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2383 net5490 vssd1 vssd1 vccd1 vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 net6015 vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1660 _01291_ vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1671 net5853 vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_14750_ _07891_ _07899_ _07900_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1682 net6789 vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ net3040 _05127_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__nand2_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1693 _01117_ vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03776_ clknet_0__03776_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03776_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _06591_ _06627_ _06603_ _06600_ _06677_ _06688_ vssd1 vssd1 vccd1 vccd1 _06852_
+ sky130_fd_sc_hd__mux4_1
X_10913_ net2253 net7075 _04321_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__mux2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _07817_ _07830_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__a21oi_2
X_11893_ _05055_ _05057_ _05060_ _05062_ _05030_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a221o_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ _09227_ _09371_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13632_ _06773_ _06774_ _06677_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__a21oi_1
X_10844_ net7221 net7069 _04288_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16351_ _09327_ _09331_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13563_ _06657_ _06658_ _06713_ _06661_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__a22o_2
X_10775_ net7292 net7193 _04255_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15302_ _08375_ _08376_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12514_ _05229_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or2_1
X_19070_ net6029 _03009_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__or2_1
X_16282_ _09350_ _09355_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__xnor2_2
X_13494_ _06485_ _06555_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18021_ _02067_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ net4310 _08305_ _08307_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__a21o_1
X_12445_ net4093 _05318_ _05611_ _05309_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_23_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ net4933 vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__buf_4
X_12376_ rbzero.tex_g1\[57\] rbzero.tex_g1\[56\] _05483_ vssd1 vssd1 vccd1 vccd1 _05543_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14115_ _07264_ _07265_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__xor2_1
X_11327_ net6726 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20962__371 clknet_1_0__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__inv_2
X_19972_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__buf_2
XFILLER_0_61_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ _08195_ vssd1 vssd1 vccd1 vccd1 _08215_ sky130_fd_sc_hd__buf_2
XFILLER_0_197_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ _06862_ _06990_ _07196_ _07194_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o31ai_1
X_18923_ _02879_ _02880_ _02905_ net4816 net4758 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a311o_1
X_11258_ net2585 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18854_ net6069 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__clkbuf_1
X_11189_ net2201 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17805_ _10581_ _01855_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__xnor2_1
X_15997_ _09041_ _09071_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__or2_1
X_18785_ _02769_ _02770_ _02771_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17736_ _01779_ _01680_ _01785_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14948_ _08070_ _08093_ _08069_ vssd1 vssd1 vccd1 vccd1 _08094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17667_ _10545_ _10546_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nor2_1
X_14879_ net7908 _07998_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19406_ net5536 _03211_ _03216_ _03207_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__o211a_1
X_16618_ _09671_ _09688_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__xor2_2
XFILLER_0_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17598_ _10594_ _10595_ vssd1 vssd1 vccd1 vccd1 _10596_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16549_ _09592_ _09620_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19337_ net4191 _03172_ net1084 _03168_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19268_ net5161 _03133_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6605 net2599 vssd1 vssd1 vccd1 vccd1 net7129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6616 rbzero.tex_r1\[34\] vssd1 vssd1 vccd1 vccd1 net7140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18219_ net4577 _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__xor2_1
X_19199_ net2975 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
Xhold6627 net2642 vssd1 vssd1 vccd1 vccd1 net7151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6638 rbzero.tex_r0\[36\] vssd1 vssd1 vccd1 vccd1 net7162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5904 rbzero.tex_b0\[40\] vssd1 vssd1 vccd1 vccd1 net6428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6649 net2307 vssd1 vssd1 vccd1 vccd1 net7173 sky130_fd_sc_hd__dlygate4sd3_1
X_21230_ clknet_leaf_52_i_clk _00399_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold5915 net1259 vssd1 vssd1 vccd1 vccd1 net6439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5926 _04411_ vssd1 vssd1 vccd1 vccd1 net6450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 net3523 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5937 net1357 vssd1 vssd1 vccd1 vccd1 net6461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 net4990 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold223 rbzero.pov.ready_buffer\[56\] vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5948 rbzero.tex_b1\[0\] vssd1 vssd1 vccd1 vccd1 net6472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5959 net1502 vssd1 vssd1 vccd1 vccd1 net6483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 net5060 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ _04137_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__buf_1
Xhold245 net5071 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 net4984 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 net5092 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20112_ net3563 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
Xhold278 net5133 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21092_ _04081_ _04082_ _04083_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold289 net5021 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20043_ _03616_ net3839 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__or2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ net219 net2148 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20790__216 clknet_1_1__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__inv_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22477_ clknet_leaf_77_i_clk net655 vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
X_12230_ _05391_ _05381_ _05392_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a211o_1
X_21428_ clknet_leaf_44_i_clk net3282 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12161_ net4037 net4009 net3761 vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__or3_1
X_21359_ clknet_leaf_58_i_clk _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11112_ net7255 net7217 _04426_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
X_12092_ _05229_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__clkbuf_8
Xhold790 net3411 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ _08890_ _08937_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__xor2_2
X_11043_ net6385 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15851_ _08913_ _08925_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__xnor2_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2180 _01539_ vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2191 _04311_ vssd1 vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
X_14802_ _07952_ _07930_ _07933_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15782_ _08405_ _08422_ _08432_ _08455_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__or4_1
X_18570_ net7586 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__inv_2
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _06148_ _06149_ _06119_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1490 net597 vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
X_17521_ _08873_ vssd1 vssd1 vccd1 vccd1 _10520_ sky130_fd_sc_hd__clkbuf_4
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _07851_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__xor2_1
X_11945_ net3378 _05095_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__or2_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _10327_ _10450_ _10325_ vssd1 vssd1 vccd1 vccd1 _10452_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ _07768_ _07781_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__xnor2_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _04988_ vssd1 vssd1 vccd1 vccd1 _05046_
+ sky130_fd_sc_hd__mux2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _08587_ _09216_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ _06732_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__nand2_1
X_10827_ net7262 net6712 _04277_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__mux2_1
X_17383_ _08548_ vssd1 vssd1 vccd1 vccd1 _10383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14595_ _07534_ _07399_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16334_ _09278_ _09292_ _09407_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19122_ _03036_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__buf_2
X_13546_ _06693_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__buf_2
X_10758_ net2101 net7121 _04244_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19053_ net3096 _03009_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__or2_1
X_16265_ _08529_ _08471_ _09193_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13477_ _06600_ _06597_ _06588_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__and4b_2
X_10689_ net7209 net2855 _04203_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18004_ _02031_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__xnor2_1
X_15216_ net3511 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__clkbuf_1
X_12428_ _05593_ _05594_ _04993_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__mux2_1
X_16196_ _09268_ _09270_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15147_ net4580 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
X_12359_ net7322 net1027 _05120_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3809 net7822 vssd1 vssd1 vccd1 vccd1 net4333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15078_ net4528 net4499 _08191_ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__mux2_1
X_19955_ net6213 _03532_ net748 _03519_ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ _07135_ net551 vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__xor2_1
X_18906_ net4662 _02883_ net7580 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a21o_1
X_19886_ net6182 _03475_ net676 _03496_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__o211a_1
X_18837_ net3807 _05393_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ _02760_ net4551 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17719_ _01768_ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18699_ _02702_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__04007_ clknet_0__04007_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04007_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22400_ net152 net2407 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
Xhold7103 _02843_ vssd1 vssd1 vccd1 vccd1 net7627 sky130_fd_sc_hd__dlygate4sd3_1
X_20592_ net3526 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7114 rbzero.pov.ready_buffer\[28\] vssd1 vssd1 vccd1 vccd1 net7638 sky130_fd_sc_hd__dlygate4sd3_1
X_20969__377 clknet_1_1__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__inv_2
XFILLER_0_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7125 rbzero.spi_registers.texadd2\[23\] vssd1 vssd1 vccd1 vccd1 net7649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22331_ net463 net2423 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7136 rbzero.spi_registers.texadd2\[12\] vssd1 vssd1 vccd1 vccd1 net7660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6402 net2166 vssd1 vssd1 vccd1 vccd1 net6926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7147 rbzero.row_render.texu\[1\] vssd1 vssd1 vccd1 vccd1 net7671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6413 rbzero.tex_b1\[14\] vssd1 vssd1 vccd1 vccd1 net6937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6424 net2030 vssd1 vssd1 vccd1 vccd1 net6948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6435 _04379_ vssd1 vssd1 vccd1 vccd1 net6959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5701 net1726 vssd1 vssd1 vccd1 vccd1 net6225 sky130_fd_sc_hd__dlygate4sd3_1
X_22262_ net394 net2739 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
Xhold6446 net2511 vssd1 vssd1 vccd1 vccd1 net6970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6457 rbzero.tex_g1\[26\] vssd1 vssd1 vccd1 vccd1 net6981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5712 net1883 vssd1 vssd1 vccd1 vccd1 net6236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6468 net2143 vssd1 vssd1 vccd1 vccd1 net6992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5723 _00803_ vssd1 vssd1 vccd1 vccd1 net6247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6479 rbzero.tex_r0\[60\] vssd1 vssd1 vccd1 vccd1 net7003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5734 net1604 vssd1 vssd1 vccd1 vccd1 net6258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5745 rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 net6269 sky130_fd_sc_hd__dlygate4sd3_1
X_21213_ net6341 net4959 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__xnor2_1
X_22193_ net325 net635 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold5756 _00422_ vssd1 vssd1 vccd1 vccd1 net6280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5767 _03270_ vssd1 vssd1 vccd1 vccd1 net6291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5778 net1534 vssd1 vssd1 vccd1 vccd1 net6302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5789 net3991 vssd1 vssd1 vccd1 vccd1 net6313 sky130_fd_sc_hd__dlygate4sd3_1
X_21144_ net3402 net2982 _04626_ net3980 _08200_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a41o_1
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21075_ net4167 net4503 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__04800_ clknet_0__04800_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04800_
+ sky130_fd_sc_hd__clkbuf_16
X_20026_ _04241_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ net202 net2075 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer60 _06781_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer71 _06868_ vssd1 vssd1 vccd1 vccd1 net3405 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ net1185 _04899_ net3620 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o21a_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ net6330 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__buf_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _06549_ _06539_ _06550_ _06541_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__a31o_1
X_10612_ net7026 net2686 _04170_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ _07529_ _07530_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11592_ rbzero.spi_registers.texadd0\[3\] _04680_ _04762_ _04763_ _04724_ vssd1 vssd1
+ vccd1 vccd1 _04764_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13331_ _06465_ _06468_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16050_ _09111_ _09124_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20297__34 clknet_1_0__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
X_13262_ _06393_ _06412_ _06413_ _06394_ net5510 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ _07989_ _07993_ _06690_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__mux2_4
X_12213_ _05360_ _05376_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__nor2_2
X_13193_ net2677 _06219_ _06196_ net2823 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _05194_ _04599_ _04602_ _04801_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19740_ net6066 _03408_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__or2_1
X_12075_ _04999_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__clkbuf_8
X_16952_ net2807 _09968_ net4877 vssd1 vssd1 vccd1 vccd1 _09969_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_194_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11026_ net2132 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__clkbuf_1
X_15903_ _08974_ _08977_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__xnor2_1
X_19671_ net3022 _03374_ net1648 _03371_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__o211a_1
X_16883_ net6023 _09934_ _09936_ _08117_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18622_ _02630_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15834_ _08898_ _08907_ _08908_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__a21oi_2
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20773__200 clknet_1_1__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__inv_2
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ net6080 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__clkbuf_1
X_15765_ _08387_ _08411_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__nor2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _06094_ _06130_ _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a31o_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _10399_ _10473_ _10501_ vssd1 vssd1 vccd1 vccd1 _10503_ sky130_fd_sc_hd__nand3_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ _05008_ _05002_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__or3_1
X_14716_ _07859_ _07860_ _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__a21o_1
X_15696_ _08683_ _08685_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__or2_1
X_18484_ net3925 net3960 _02495_ _02499_ _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__o311a_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _10279_ _10309_ _10434_ vssd1 vssd1 vccd1 vccd1 _10435_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14647_ _07532_ _07358_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11859_ _04979_ _05001_ _05011_ _05024_ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__o311a_1
XFILLER_0_185_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _10356_ _10365_ vssd1 vssd1 vccd1 vccd1 _10366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14578_ _07728_ _07725_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19105_ net5562 _03040_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__or2_1
X_16317_ _09206_ _09241_ _09390_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__a21oi_1
X_13529_ _06612_ _06565_ _06587_ _06679_ _06579_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__a311o_1
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17297_ _09870_ _10169_ vssd1 vssd1 vccd1 vccd1 _10298_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ _09320_ _09321_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19036_ net3934 _02988_ _02999_ _02993_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__o211a_1
Xhold5008 rbzero.pov.spi_buffer\[34\] vssd1 vssd1 vccd1 vccd1 net5532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5019 rbzero.pov.spi_buffer\[24\] vssd1 vssd1 vccd1 vccd1 net5543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16179_ _08310_ _08795_ _09251_ _08326_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__o22a_1
Xhold4307 net2961 vssd1 vssd1 vccd1 vccd1 net4831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4318 net1356 vssd1 vssd1 vccd1 vccd1 net4842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4329 rbzero.pov.spi_buffer\[60\] vssd1 vssd1 vccd1 vccd1 net4853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3606 net7633 vssd1 vssd1 vccd1 vccd1 net4130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3617 net7471 vssd1 vssd1 vccd1 vccd1 net4141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3628 rbzero.traced_texa\[-4\] vssd1 vssd1 vccd1 vccd1 net4152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3639 net7501 vssd1 vssd1 vccd1 vccd1 net4163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2905 _03796_ vssd1 vssd1 vccd1 vccd1 net3429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2916 net927 vssd1 vssd1 vccd1 vccd1 net3440 sky130_fd_sc_hd__dlygate4sd3_1
X_19938_ net3917 _08473_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nand2_1
Xhold2927 _03827_ vssd1 vssd1 vccd1 vccd1 net3451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2938 net3283 vssd1 vssd1 vccd1 vccd1 net3462 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2949 net7551 vssd1 vssd1 vccd1 vccd1 net3473 sky130_fd_sc_hd__dlygate4sd3_1
X_19869_ net1013 _03470_ _03480_ _08481_ _03475_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o221a_1
X_21900_ clknet_leaf_95_i_clk net1434 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21831_ clknet_leaf_87_i_clk net3658 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21762_ clknet_leaf_24_i_clk net1966 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20713_ clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__buf_1
X_21693_ clknet_leaf_25_i_clk net5393 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20644_ net3979 net4017 _03974_ net3937 _04597_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20575_ net2999 net3670 _03911_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__mux2_1
Xhold6210 net1948 vssd1 vssd1 vccd1 vccd1 net6734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6221 rbzero.tex_b0\[37\] vssd1 vssd1 vccd1 vccd1 net6745 sky130_fd_sc_hd__dlygate4sd3_1
X_22314_ net446 net2056 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold6232 net2349 vssd1 vssd1 vccd1 vccd1 net6756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6243 rbzero.tex_g1\[13\] vssd1 vssd1 vccd1 vccd1 net6767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6254 net1979 vssd1 vssd1 vccd1 vccd1 net6778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5520 _03390_ vssd1 vssd1 vccd1 vccd1 net6044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6265 rbzero.tex_b1\[34\] vssd1 vssd1 vccd1 vccd1 net6789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22245_ net377 net2242 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold6276 net1804 vssd1 vssd1 vccd1 vccd1 net6800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5531 net1574 vssd1 vssd1 vccd1 vccd1 net6055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6287 _04519_ vssd1 vssd1 vccd1 vccd1 net6811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5542 net1644 vssd1 vssd1 vccd1 vccd1 net6066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6298 net1894 vssd1 vssd1 vccd1 vccd1 net6822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5553 _03422_ vssd1 vssd1 vccd1 vccd1 net6077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5564 _02786_ vssd1 vssd1 vccd1 vccd1 net6088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4830 _00714_ vssd1 vssd1 vccd1 vccd1 net5354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5575 _08232_ vssd1 vssd1 vccd1 vccd1 net6099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4841 _00729_ vssd1 vssd1 vccd1 vccd1 net5365 sky130_fd_sc_hd__dlygate4sd3_1
X_22176_ net308 net2273 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold5586 rbzero.spi_registers.buf_texadd3\[19\] vssd1 vssd1 vccd1 vccd1 net6110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4852 _00829_ vssd1 vssd1 vccd1 vccd1 net5376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4863 net1318 vssd1 vssd1 vccd1 vccd1 net5387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4874 net1056 vssd1 vssd1 vccd1 vccd1 net5398 sky130_fd_sc_hd__dlygate4sd3_1
X_21127_ net4133 net4740 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__nor2_1
Xhold4885 rbzero.pov.spi_buffer\[7\] vssd1 vssd1 vccd1 vccd1 net5409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4896 net977 vssd1 vssd1 vccd1 vccd1 net5420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21058_ _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__and2b_1
XFILLER_0_191_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12900_ net37 net36 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or2_1
X_20009_ rbzero.debug_overlay.facingY\[-6\] net3743 _03594_ vssd1 vssd1 vccd1 vccd1
+ _03605_ sky130_fd_sc_hd__mux2_1
X_13880_ _07025_ _07030_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _05945_ _05988_ _05989_ _05957_ _05947_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a221o_2
XFILLER_0_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ net4335 _06210_ _08601_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__o21ai_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ net19 net20 _05918_ _05920_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a32o_1
XFILLER_0_189_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _06957_ _07532_ _07463_ _07438_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__or4_4
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ net2791 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__inv_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15481_ _08298_ _08554_ _08555_ _08307_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__a211o_4
XFILLER_0_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ net10 net11 vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__nor2b_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17220_ _10147_ _10129_ vssd1 vssd1 vccd1 vccd1 _10221_ sky130_fd_sc_hd__or2b_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _07581_ _07582_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__and2_1
X_11644_ net4009 net3761 net4052 net4037 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17151_ _08584_ _10152_ _09865_ vssd1 vssd1 vccd1 vccd1 _10153_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14363_ _07361_ _07403_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
X_11575_ _04718_ _04687_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__or3b_1
Xinput27 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dlymetal6s2s_1
X_16102_ _08995_ _09176_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_4
X_13314_ _06445_ _06459_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__a21o_1
X_17082_ net3578 net4334 vssd1 vssd1 vccd1 vccd1 _10084_ sky130_fd_sc_hd__nand2_1
Xinput49 i_test_uc2 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_165_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ _07362_ _07397_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _09103_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ net4887 _06179_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13176_ _06328_ _06331_ _06292_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a21oi_1
X_20805__229 clknet_1_1__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__inv_2
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ net4077 _05206_ _05213_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__o2bb2a_1
X_17984_ _01825_ _01941_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19723_ _03392_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12058_ rbzero.tex_r1\[61\] rbzero.tex_r1\[60\] _05071_ vssd1 vssd1 vccd1 vccd1 _05227_
+ sky130_fd_sc_hd__mux2_1
X_16935_ _06213_ _09294_ vssd1 vssd1 vccd1 vccd1 _09953_ sky130_fd_sc_hd__xnor2_1
X_11009_ net5879 net6778 _04377_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__mux2_1
X_19654_ _03000_ _03360_ net1830 _03354_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__o211a_1
X_16866_ _09925_ _09920_ net4055 vssd1 vssd1 vccd1 vccd1 _09927_ sky130_fd_sc_hd__and3b_1
XFILLER_0_137_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18605_ net4666 net3796 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__xor2_1
XFILLER_0_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15817_ _08347_ _08393_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19585_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__buf_2
X_16797_ _09865_ _09866_ vssd1 vssd1 vccd1 vccd1 _09867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18536_ _02549_ net6239 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__or2_1
X_15748_ _08808_ _08822_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__xor2_2
XFILLER_0_158_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18467_ _02489_ vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15679_ _08314_ _08546_ _08547_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17418_ _09138_ _10168_ _10174_ _09139_ vssd1 vssd1 vccd1 vccd1 _10418_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18398_ _02261_ _02428_ _02429_ _10455_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17349_ _10347_ _10348_ vssd1 vssd1 vccd1 vccd1 _10349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03987_ clknet_0__03987_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03987_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19019_ net6271 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__buf_1
Xhold4104 net7577 vssd1 vssd1 vccd1 vccd1 net4628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4115 net3793 vssd1 vssd1 vccd1 vccd1 net4639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4126 _01605_ vssd1 vssd1 vccd1 vccd1 net4650 sky130_fd_sc_hd__dlygate4sd3_1
X_22030_ clknet_leaf_96_i_clk net3731 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3403 _03467_ vssd1 vssd1 vccd1 vccd1 net3927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4148 net1700 vssd1 vssd1 vccd1 vccd1 net4672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4159 net3026 vssd1 vssd1 vccd1 vccd1 net4683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3414 _01263_ vssd1 vssd1 vccd1 vccd1 net3938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3425 net1607 vssd1 vssd1 vccd1 vccd1 net3949 sky130_fd_sc_hd__dlygate4sd3_1
X_20745__176 clknet_1_0__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__inv_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3436 net7314 vssd1 vssd1 vccd1 vccd1 net3960 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3447 net88 vssd1 vssd1 vccd1 vccd1 net3971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2702 _03654_ vssd1 vssd1 vccd1 vccd1 net3226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3458 _01614_ vssd1 vssd1 vccd1 vccd1 net3982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2724 _00601_ vssd1 vssd1 vccd1 vccd1 net3248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3469 _04163_ vssd1 vssd1 vccd1 vccd1 net3993 sky130_fd_sc_hd__buf_4
Xhold2735 _03918_ vssd1 vssd1 vccd1 vccd1 net3259 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2746 _03784_ vssd1 vssd1 vccd1 vccd1 net3270 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2757 _02745_ vssd1 vssd1 vccd1 vccd1 net3281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2768 _03830_ vssd1 vssd1 vccd1 vccd1 net3292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2779 _03877_ vssd1 vssd1 vccd1 vccd1 net3303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21814_ clknet_leaf_9_i_clk net3084 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21745_ clknet_leaf_0_i_clk net2096 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20910__324 clknet_1_1__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__inv_2
XFILLER_0_175_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21676_ clknet_leaf_14_i_clk net842 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdy\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20627_ _05299_ _09929_ _03031_ _03957_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ net6832 net2430 _04562_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__mux2_1
X_20558_ net3478 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6040 net1628 vssd1 vssd1 vccd1 vccd1 net6564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6051 _04406_ vssd1 vssd1 vccd1 vccd1 net6575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6062 net1647 vssd1 vssd1 vccd1 vccd1 net6586 sky130_fd_sc_hd__dlygate4sd3_1
X_11291_ net7087 net6692 _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__mux2_1
Xhold6073 rbzero.tex_b0\[9\] vssd1 vssd1 vccd1 vccd1 net6597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20489_ net3139 net3530 _03867_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6084 net1667 vssd1 vssd1 vccd1 vccd1 net6608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5350 net2465 vssd1 vssd1 vccd1 vccd1 net5874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6095 _04402_ vssd1 vssd1 vccd1 vccd1 net6619 sky130_fd_sc_hd__dlygate4sd3_1
X_13030_ net6185 vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__clkbuf_4
Xhold5361 rbzero.tex_r1\[3\] vssd1 vssd1 vccd1 vccd1 net5885 sky130_fd_sc_hd__dlygate4sd3_1
X_22228_ net360 net2099 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold5372 rbzero.tex_g1\[33\] vssd1 vssd1 vccd1 vccd1 net5896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5383 rbzero.map_overlay.i_otherx\[0\] vssd1 vssd1 vccd1 vccd1 net5907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5394 net2802 vssd1 vssd1 vccd1 vccd1 net5918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4660 net959 vssd1 vssd1 vccd1 vccd1 net5184 sky130_fd_sc_hd__dlygate4sd3_1
X_22159_ net291 net1520 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4671 net1291 vssd1 vssd1 vccd1 vccd1 net5195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4682 _01082_ vssd1 vssd1 vccd1 vccd1 net5206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4693 _00845_ vssd1 vssd1 vccd1 vccd1 net5217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3970 _03625_ vssd1 vssd1 vccd1 vccd1 net4494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3981 net1167 vssd1 vssd1 vccd1 vccd1 net4505 sky130_fd_sc_hd__dlygate4sd3_1
X_14981_ _08068_ _08123_ net6162 vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__a21oi_1
Xhold3992 _00997_ vssd1 vssd1 vccd1 vccd1 net4516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16720_ net7554 _06211_ _08314_ vssd1 vssd1 vccd1 vccd1 _09790_ sky130_fd_sc_hd__and3_1
X_13932_ _06865_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16651_ _09720_ _09721_ vssd1 vssd1 vccd1 vccd1 _09722_ sky130_fd_sc_hd__xnor2_1
X_13863_ _06876_ _06859_ _06875_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__or3_1
XFILLER_0_199_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15602_ _08675_ _08676_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__and2_1
X_12814_ net24 _05951_ _05972_ net26 vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19370_ net1214 _03186_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__or2_1
X_16582_ _09637_ _09638_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__nor2_2
X_13794_ _06887_ _06890_ _06889_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18321_ net4591 net4382 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12745_ net16 net17 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__nor2b_2
X_15533_ _06133_ _06570_ net4086 vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__mux2_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18252_ _01778_ _09310_ _02222_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__o31a_1
XFILLER_0_132_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _08304_ _08538_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__nor2_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12676_ _05815_ _05837_ net9 vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17203_ _10202_ _10204_ vssd1 vssd1 vccd1 vccd1 _10205_ sky130_fd_sc_hd__xor2_4
X_14415_ _07493_ _07564_ _07563_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__nand3_4
X_20885__301 clknet_1_1__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__inv_2
X_11627_ net73 _04793_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and3b_1
X_18183_ _02228_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__xor2_1
X_15395_ _08312_ _08466_ _08469_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_167_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17134_ _10134_ _10135_ vssd1 vssd1 vccd1 vccd1 _10136_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14346_ _07356_ _07439_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11558_ _04696_ _04697_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold608 net1637 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ _10058_ _10059_ net3398 vssd1 vssd1 vccd1 vccd1 _10069_ sky130_fd_sc_hd__o21ai_1
Xhold619 net4198 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14277_ _07426_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_204_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ rbzero.texu_hot\[1\] _04657_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__or2_1
X_16016_ _09090_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__clkbuf_4
X_13228_ net4917 net4900 vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _06314_ net3174 _06308_ net3233 vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a22o_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 net6201 vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 net5847 vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
X_17967_ _01932_ _01988_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a21o_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1319 _01479_ vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19706_ net6682 _03395_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16918_ net4160 _09941_ _09942_ net6150 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a22o_1
X_17898_ _01935_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__xnor2_1
X_19637_ net1613 _03326_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__or2_1
X_16849_ _04241_ net3979 vssd1 vssd1 vccd1 vccd1 _09918_ sky130_fd_sc_hd__or2_1
X_19568_ net5014 _03303_ _03316_ _03314_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__o211a_1
X_18519_ net4446 net4806 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19499_ _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21530_ clknet_leaf_27_i_clk net3131 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21461_ clknet_leaf_30_i_clk net3959 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20412_ net3453 net1162 _03801_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
X_21392_ clknet_leaf_61_i_clk _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20274_ net3670 net4839 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__or2_1
Xhold3200 _00413_ vssd1 vssd1 vccd1 vccd1 net3724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22013_ clknet_leaf_97_i_clk net3639 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3211 _01238_ vssd1 vssd1 vccd1 vccd1 net3735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3222 _00999_ vssd1 vssd1 vccd1 vccd1 net3746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3233 _03832_ vssd1 vssd1 vccd1 vccd1 net3757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2510 net6308 vssd1 vssd1 vccd1 vccd1 net3034 sky130_fd_sc_hd__buf_1
Xhold3255 net7767 vssd1 vssd1 vccd1 vccd1 net3779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2521 net4813 vssd1 vssd1 vccd1 vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3277 _03898_ vssd1 vssd1 vccd1 vccd1 net3801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2532 net4785 vssd1 vssd1 vccd1 vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3288 net1483 vssd1 vssd1 vccd1 vccd1 net3812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2543 _08216_ vssd1 vssd1 vccd1 vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2554 _03254_ vssd1 vssd1 vccd1 vccd1 net3078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3299 _02946_ vssd1 vssd1 vccd1 vccd1 net3823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1820 _04205_ vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 _00641_ vssd1 vssd1 vccd1 vccd1 net3089 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1831 net6077 vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2576 net1546 vssd1 vssd1 vccd1 vccd1 net3100 sky130_fd_sc_hd__clkbuf_4
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1842 rbzero.tex_r0\[63\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2587 rbzero.spi_registers.spi_buffer\[6\] vssd1 vssd1 vccd1 vccd1 net3111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1853 _04293_ vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 net4733 vssd1 vssd1 vccd1 vccd1 net3122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1864 net7650 vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__clkbuf_2
Xhold1875 net7029 vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1886 _01116_ vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1897 net6935 vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10860_ net2144 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ net6467 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__clkbuf_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ _04818_ net3535 net2 vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__o21ai_2
X_21728_ clknet_leaf_2_i_clk net1702 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _05261_ _05626_ _05244_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21659_ clknet_leaf_16_i_clk net5047 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_othery\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14200_ _07307_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__or2_4
X_11412_ net6798 net2370 _04584_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_1
X_15180_ net4639 _08177_ _08260_ vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__mux2_1
X_12392_ rbzero.tex_g1\[41\] rbzero.tex_g1\[40\] _05456_ vssd1 vssd1 vccd1 vccd1 _05559_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_94 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_94/HI o_rgb[4] sky130_fd_sc_hd__conb_1
XFILLER_0_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ _06895_ _06858_ _07280_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__o21ai_1
X_11343_ net6746 net2051 _04551_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14062_ _07209_ _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nor2_1
X_11274_ net2436 net6337 _04514_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20728__160 clknet_1_1__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__inv_2
Xhold5180 net1403 vssd1 vssd1 vccd1 vccd1 net5704 sky130_fd_sc_hd__dlygate4sd3_1
X_13013_ _06156_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__nor2_1
Xhold5191 _00752_ vssd1 vssd1 vccd1 vccd1 net5715 sky130_fd_sc_hd__dlygate4sd3_1
X_18870_ _02822_ _02833_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a21o_1
X_17821_ _01867_ _01868_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a21o_1
Xhold4490 net755 vssd1 vssd1 vccd1 vccd1 net5014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ _01802_ _01778_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__nor2_1
X_14964_ _08090_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__inv_2
X_16703_ _09645_ _09647_ _09644_ vssd1 vssd1 vccd1 vccd1 _09774_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13915_ _07060_ _07061_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17683_ _01732_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__xor2_1
X_14895_ net7568 _08039_ _08044_ _06589_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_18_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19422_ net1718 _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__or2_1
X_16634_ _09703_ _09704_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13846_ _06974_ _06975_ _06996_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19353_ net2455 _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__or2_1
X_16565_ _09531_ _09636_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13777_ _06926_ _06927_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ net2005 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18304_ net4687 net4455 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15516_ _08155_ vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12728_ net15 _05880_ _05888_ _05842_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a22o_2
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19284_ net1652 _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__or2_1
X_16496_ _09328_ _08707_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18235_ _02176_ _02200_ _02177_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o21ba_1
X_15447_ _08513_ _08521_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ net6 _05791_ _05820_ net8 vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6809 _03607_ vssd1 vssd1 vccd1 vccd1 net7333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18166_ _10383_ _09805_ _02120_ _02118_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__o31a_1
XFILLER_0_142_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ net3193 _08304_ _08307_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17117_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10119_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14329_ _07471_ _07439_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__nor2_1
Xhold405 rbzero.spi_registers.buf_mapdx\[4\] vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ _02128_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold416 net5319 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold427 net7647 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_141_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold438 net5359 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ _10050_ _10053_ vssd1 vssd1 vccd1 vccd1 _10054_ sky130_fd_sc_hd__xnor2_1
Xhold449 net5278 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 net6565 vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
X_18999_ net7355 _02967_ net3890 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__and3b_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _00920_ vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1127 net5774 vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1138 _03435_ vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 net4277 vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__buf_1
XFILLER_0_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21513_ clknet_leaf_36_i_clk net5515 vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21444_ clknet_leaf_86_i_clk net4873 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21375_ clknet_leaf_64_i_clk _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold950 _01517_ vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 net6593 vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 net4255 vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
X_20257_ net4845 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__clkbuf_4
Xhold983 net5734 vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 net6546 vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3030 net4612 vssd1 vssd1 vccd1 vccd1 net3554 sky130_fd_sc_hd__buf_1
X_11630__1 clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
Xhold3041 net4604 vssd1 vssd1 vccd1 vccd1 net3565 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3052 _01220_ vssd1 vssd1 vccd1 vccd1 net3576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3063 _03803_ vssd1 vssd1 vccd1 vccd1 net3587 sky130_fd_sc_hd__dlygate4sd3_1
X_20188_ _03675_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__clkbuf_4
Xhold3074 net1362 vssd1 vssd1 vccd1 vccd1 net3598 sky130_fd_sc_hd__buf_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 net5958 vssd1 vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3085 _01186_ vssd1 vssd1 vccd1 vccd1 net3609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 net6034 vssd1 vssd1 vccd1 vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3096 _04893_ vssd1 vssd1 vccd1 vccd1 net3620 sky130_fd_sc_hd__buf_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2362 _00600_ vssd1 vssd1 vccd1 vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2373 net7295 vssd1 vssd1 vccd1 vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2384 net5492 vssd1 vssd1 vccd1 vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1650 _04484_ vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2395 rbzero.wall_tracer.rayAddendX\[-4\] vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1661 net7053 vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ net2869 net2069 _05128_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1672 rbzero.tex_b1\[27\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1683 _04490_ vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 net6939 vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03775_ clknet_0__03775_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03775_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10912_ net7077 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__clkbuf_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _06421_ _06663_ _06713_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__and3_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _07818_ _07829_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__nor2_1
X_11892_ _05061_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__buf_4
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13631_ _06747_ _06748_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10843_ net6502 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__clkbuf_1
X_16350_ _09422_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__inv_2
X_13562_ _06675_ _06686_ _06667_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__a21o_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10774_ net7081 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__clkbuf_1
X_12513_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _05230_ vssd1 vssd1 vccd1 vccd1 _05679_
+ sky130_fd_sc_hd__mux2_1
X_15301_ net2942 _08354_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__nand2_1
X_16281_ _09353_ _09354_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _06638_ _06595_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18020_ _02067_ _02068_ _06205_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15232_ _08306_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__clkbuf_8
X_12444_ _04892_ _05319_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _08259_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__clkbuf_1
X_12375_ rbzero.tex_g1\[59\] rbzero.tex_g1\[58\] _05541_ vssd1 vssd1 vccd1 vccd1 _05542_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ _06737_ _06990_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nor2_1
X_11326_ net6724 net2316 _04540_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19971_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__clkbuf_4
X_15094_ net6253 _08201_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _07194_ _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nand2_1
X_18922_ rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\] _02854_
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o21a_1
X_11257_ net6862 net6938 _04503_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18853_ rbzero.wall_tracer.rayAddendY\[2\] _02841_ _02714_ vssd1 vssd1 vccd1 vccd1
+ _02842_ sky130_fd_sc_hd__mux2_1
X_11188_ net6387 net6842 _04470_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17804_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__xor2_1
X_18784_ net4640 _02768_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__or2_1
X_15996_ _09062_ _09069_ _09070_ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_59_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17735_ _01779_ _01680_ _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a21oi_1
X_14947_ _08037_ _08040_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__or2_1
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17666_ _01709_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14878_ _08028_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19405_ net1964 _03212_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__or2_1
X_16617_ _09686_ _09687_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13829_ _06965_ _06979_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__xnor2_2
X_17597_ _09328_ net7378 vssd1 vssd1 vccd1 vccd1 _10595_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19336_ net1083 _03173_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16548_ _09617_ _09619_ vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19267_ net5452 _03132_ _03137_ _03128_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__o211a_1
X_16479_ _09549_ _09550_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18218_ _02257_ _02259_ _02256_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a21bo_1
Xhold6606 _04380_ vssd1 vssd1 vccd1 vccd1 net7130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6617 net2568 vssd1 vssd1 vccd1 vccd1 net7141 sky130_fd_sc_hd__dlygate4sd3_1
X_19198_ _03088_ net2974 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6628 rbzero.tex_r1\[53\] vssd1 vssd1 vccd1 vccd1 net7152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6639 net2644 vssd1 vssd1 vccd1 vccd1 net7163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5905 net1196 vssd1 vssd1 vccd1 vccd1 net6429 sky130_fd_sc_hd__dlygate4sd3_1
X_18149_ _02188_ _02195_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__xnor2_1
Xhold5916 rbzero.tex_b1\[56\] vssd1 vssd1 vccd1 vccd1 net6440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 _03518_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5927 net1192 vssd1 vssd1 vccd1 vccd1 net6451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5938 _04591_ vssd1 vssd1 vccd1 vccd1 net6462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold213 net4992 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5949 net1480 vssd1 vssd1 vccd1 vccd1 net6473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _03567_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold235 net5062 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ _02488_ clknet_1_0__leaf__05994_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_2
Xhold246 net5073 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold257 net5033 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
X_20111_ _03670_ net3562 net7330 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__and3b_1
Xhold268 net5056 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold279 net4998 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21091_ _04081_ _04082_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20042_ net3838 net3453 _03594_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21993_ net218 net1740 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22476_ clknet_3_5_0_i_clk net1922 vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21427_ clknet_leaf_44_i_clk net3896 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_1
X_20312__47 clknet_1_0__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12160_ _04814_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__or2_2
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21358_ clknet_leaf_42_i_clk net5422 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11111_ net6718 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
X_12091_ _05235_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__or2_1
Xhold780 net7740 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
X_21289_ clknet_leaf_75_i_clk net4008 vssd1 vssd1 vccd1 vccd1 reg_rgb\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold791 net5688 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__05994_ clknet_0__05994_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__05994_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net6383 net1950 _04392_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__mux2_1
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _08914_ _08923_ _08924_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__a21bo_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2170 _01120_ vssd1 vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _07891_ _07951_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2181 net5943 vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__clkbuf_2
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 _01462_ vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _08821_ _08839_ _08854_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__a21o_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _06095_ _06104_ _06108_ _06115_ _06118_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__o41a_1
XFILLER_0_118_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1480 net6985 vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _10517_ _10518_ vssd1 vssd1 vccd1 vccd1 _10519_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _07874_ _07873_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__and2b_1
Xhold1491 _03445_ vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
X_11944_ net3014 _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__xnor2_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _10325_ _10202_ _10450_ vssd1 vssd1 vccd1 vccd1 _10451_ sky130_fd_sc_hd__or3b_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ _05003_ _05044_ _04999_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__o21a_1
X_14663_ _07811_ _07813_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__nor2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _09464_ _09474_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__xnor2_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ net2903 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__clkbuf_1
X_13614_ net7431 _06714_ net7433 vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__a21oi_4
X_17382_ _10378_ _10381_ vssd1 vssd1 vccd1 vccd1 _10382_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ _07534_ _07400_ _07744_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19121_ net5993 _03037_ _03051_ _03048_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__o211a_1
X_16333_ _09405_ _09406_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10757_ net2102 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__clkbuf_1
X_13545_ _06556_ _06595_ _06695_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__mux2_1
X_19052_ net2979 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__buf_2
X_16264_ _09336_ _09337_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _06503_ _06607_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_180_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10688_ net2779 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ _02032_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__xnor2_1
X_12427_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _05483_ vssd1 vssd1 vccd1 vccd1 _05594_
+ sky130_fd_sc_hd__mux2_1
X_15215_ _08195_ net3510 vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16195_ _08528_ _08835_ _09269_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12358_ _05117_ _05451_ _05525_ _04909_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a2bb2o_1
X_15146_ net4579 _08048_ _08249_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ net6614 net2799 _04529_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15077_ _08190_ _08199_ net6139 _01622_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__o211a_1
X_19954_ net747 _03485_ _03565_ _03566_ _03529_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o221a_1
X_12289_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14028_ _07165_ _07177_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__o21bai_1
X_18905_ _02854_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02890_
+ sky130_fd_sc_hd__xnor2_2
X_19885_ net675 _03477_ _03479_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a211o_1
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18836_ net3807 _05393_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__nor4_1
XFILLER_0_208_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18767_ net4550 _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__or2b_1
X_15979_ _09047_ _09053_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ _09562_ _09805_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__nor2_1
X_18698_ _02646_ net7146 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__or2_1
XFILLER_0_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04006_ clknet_0__04006_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04006_
+ sky130_fd_sc_hd__clkbuf_16
X_17649_ _09108_ _10406_ _10416_ _10174_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__or4_1
XFILLER_0_202_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19319_ net1859 _03160_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20591_ _03924_ net3525 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7104 rbzero.spi_registers.texadd1\[10\] vssd1 vssd1 vccd1 vccd1 net7628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7115 rbzero.wall_tracer.rayAddendX\[-5\] vssd1 vssd1 vccd1 vccd1 net7639 sky130_fd_sc_hd__dlygate4sd3_1
X_22330_ net462 net1679 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
Xhold7126 rbzero.wall_tracer.mapY\[6\] vssd1 vssd1 vccd1 vccd1 net7650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7137 rbzero.spi_registers.buf_texadd3\[7\] vssd1 vssd1 vccd1 vccd1 net7661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6403 rbzero.spi_registers.buf_texadd1\[14\] vssd1 vssd1 vccd1 vccd1 net6927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7148 rbzero.spi_registers.buf_leak\[0\] vssd1 vssd1 vccd1 vccd1 net7672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20668__106 clknet_1_1__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__inv_2
Xhold6414 net2584 vssd1 vssd1 vccd1 vccd1 net6938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6425 _04572_ vssd1 vssd1 vccd1 vccd1 net6949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22261_ net393 net2047 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold6436 net2515 vssd1 vssd1 vccd1 vccd1 net6960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6447 rbzero.tex_b1\[49\] vssd1 vssd1 vccd1 vccd1 net6971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5702 _00807_ vssd1 vssd1 vccd1 vccd1 net6226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6458 net1865 vssd1 vssd1 vccd1 vccd1 net6982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5713 rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 net6237 sky130_fd_sc_hd__buf_2
Xhold5724 net6311 vssd1 vssd1 vccd1 vccd1 net6248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6469 rbzero.tex_g0\[46\] vssd1 vssd1 vccd1 vccd1 net6993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21212_ net4959 net65 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5735 net673 vssd1 vssd1 vccd1 vccd1 net6259 sky130_fd_sc_hd__buf_2
X_22192_ net324 net2315 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold5746 rbzero.spi_registers.spi_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net6270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5757 net656 vssd1 vssd1 vccd1 vccd1 net6281 sky130_fd_sc_hd__clkbuf_2
Xhold5768 _00817_ vssd1 vssd1 vccd1 vccd1 net6292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5779 _03253_ vssd1 vssd1 vccd1 vccd1 net6303 sky130_fd_sc_hd__dlygate4sd3_1
X_21143_ _04627_ net3979 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21074_ net4167 net4503 vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__or2_1
X_20025_ net2887 _03613_ net4601 _03602_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ net201 net2053 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer50 _07078_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer61 _06945_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer72 _06846_ vssd1 vssd1 vccd1 vccd1 net3408 sky130_fd_sc_hd__clkbuf_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _04826_ _04599_ _04605_ net3995 _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a221o_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ net2687 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ rbzero.spi_registers.texadd3\[3\] _04640_ _04642_ rbzero.spi_registers.texadd2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ _04635_ _06479_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__nor3_4
XFILLER_0_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _06396_ _06411_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22459_ clknet_leaf_38_i_clk _01628_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12212_ _05341_ _05360_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__nor2_2
X_15000_ net7843 _07995_ _08061_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6970 net4410 vssd1 vssd1 vccd1 vccd1 net7494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13192_ net2905 _06244_ net4821 _04876_ net4914 vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__o221a_1
Xhold6992 _00499_ vssd1 vssd1 vccd1 vccd1 net7516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ _04836_ net4010 _04605_ net4014 _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12074_ _05235_ _05240_ _05242_ _05061_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__o211a_1
X_16951_ _09294_ vssd1 vssd1 vccd1 vccd1 _09968_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ net7012 net6998 _04310_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__mux2_1
X_15902_ _08975_ _08976_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__xnor2_1
X_19670_ net6586 _03375_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__or2_1
X_16882_ net4265 _09934_ _09936_ _08106_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a22o_1
X_18621_ net3242 net4493 _02629_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__o21ai_1
X_15833_ _08875_ _08878_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__xor2_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ rbzero.wall_tracer.rayAddendX\[-3\] _02567_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15764_ _08817_ _08818_ _08820_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__a21o_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ net3876 net3018 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__and2_1
X_17503_ _10399_ _10473_ _10501_ vssd1 vssd1 vccd1 vccd1 _10502_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _07861_ _07864_ _07865_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__a21bo_1
X_11927_ net3026 _04970_ _04985_ _04952_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__o211a_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _02497_ _02500_ _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a21o_1
X_15695_ _08762_ _08764_ _08761_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__a21bo_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _10307_ _10308_ vssd1 vssd1 vccd1 vccd1 _10434_ sky130_fd_sc_hd__nor2_1
X_14646_ _07534_ _07353_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__nor2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _05027_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10809_ net2846 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__clkbuf_1
X_17365_ _10363_ _10364_ vssd1 vssd1 vccd1 vccd1 _10365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 _05892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _04933_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nor2_1
X_14577_ _07676_ _07722_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19104_ net5944 _03037_ _03042_ _03022_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__o211a_1
X_16316_ _09238_ _09240_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13528_ _06579_ _06586_ _06581_ _06584_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and4bb_1
X_17296_ _10293_ _10296_ vssd1 vssd1 vccd1 vccd1 _10297_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19035_ _02996_ _02990_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__or2_1
X_16247_ _09203_ _09302_ _09319_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13459_ _06609_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__inv_2
Xhold5009 net1510 vssd1 vssd1 vccd1 vccd1 net5533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16178_ _08796_ _09252_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4308 rbzero.pov.spi_buffer\[63\] vssd1 vssd1 vccd1 vccd1 net4832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4319 rbzero.pov.ss_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net4843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15129_ _08195_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3607 _00508_ vssd1 vssd1 vccd1 vccd1 net4131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3618 net785 vssd1 vssd1 vccd1 vccd1 net4142 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_92_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold3629 net7619 vssd1 vssd1 vccd1 vccd1 net4153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2906 _03797_ vssd1 vssd1 vccd1 vccd1 net3430 sky130_fd_sc_hd__dlygate4sd3_1
X_19937_ net3917 _08473_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__or2_2
XFILLER_0_177_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20996__22 clknet_1_1__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2917 _03878_ vssd1 vssd1 vccd1 vccd1 net3441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2928 _01194_ vssd1 vssd1 vccd1 vccd1 net3452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2939 _08211_ vssd1 vssd1 vccd1 vccd1 net3463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19868_ net6199 _03475_ net3001 _03496_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18819_ _02807_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__xnor2_1
X_19799_ net6029 _03442_ net1845 _03441_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21830_ clknet_leaf_89_i_clk net3746 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21761_ clknet_leaf_23_i_clk net1663 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21692_ clknet_leaf_26_i_clk net5224 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20643_ net3930 _03972_ _03975_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20574_ net3754 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_45_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6200 net1753 vssd1 vssd1 vccd1 vccd1 net6724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6211 rbzero.tex_b1\[41\] vssd1 vssd1 vccd1 vccd1 net6735 sky130_fd_sc_hd__dlygate4sd3_1
X_22313_ net445 net1161 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6222 net2073 vssd1 vssd1 vccd1 vccd1 net6746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6233 rbzero.tex_b1\[18\] vssd1 vssd1 vccd1 vccd1 net6757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6244 net1741 vssd1 vssd1 vccd1 vccd1 net6768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6255 rbzero.tex_b1\[4\] vssd1 vssd1 vccd1 vccd1 net6779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5510 _00948_ vssd1 vssd1 vccd1 vccd1 net6034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6266 net2206 vssd1 vssd1 vccd1 vccd1 net6790 sky130_fd_sc_hd__dlygate4sd3_1
X_22244_ net376 net2359 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5521 _00900_ vssd1 vssd1 vccd1 vccd1 net6045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6277 rbzero.tex_g0\[53\] vssd1 vssd1 vccd1 vccd1 net6801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5532 _03421_ vssd1 vssd1 vccd1 vccd1 net6056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6288 net2606 vssd1 vssd1 vccd1 vccd1 net6812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6299 rbzero.tex_r0\[9\] vssd1 vssd1 vccd1 vccd1 net6823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5565 net3247 vssd1 vssd1 vccd1 vccd1 net6089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4820 net967 vssd1 vssd1 vccd1 vccd1 net5344 sky130_fd_sc_hd__dlygate4sd3_1
X_22175_ net307 net1987 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold4831 rbzero.color_sky\[5\] vssd1 vssd1 vccd1 vccd1 net5355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5587 net1631 vssd1 vssd1 vccd1 vccd1 net6111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4842 rbzero.spi_registers.buf_otherx\[1\] vssd1 vssd1 vccd1 vccd1 net5366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5598 _08197_ vssd1 vssd1 vccd1 vccd1 net6122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4853 net961 vssd1 vssd1 vccd1 vccd1 net5377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4864 _01077_ vssd1 vssd1 vccd1 vccd1 net5388 sky130_fd_sc_hd__dlygate4sd3_1
X_21126_ _04108_ _04109_ _04110_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4875 _00780_ vssd1 vssd1 vccd1 vccd1 net5399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4886 net1222 vssd1 vssd1 vccd1 vccd1 net5410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4897 _00527_ vssd1 vssd1 vccd1 vccd1 net5421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21057_ net4146 net4736 vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__nand2_1
X_20722__155 clknet_1_0__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__inv_2
X_20008_ net3831 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ net6357 _05945_ _05987_ net56 vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a22o_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _04760_ _04603_ _04637_ _04165_ net16 net17 vssd1 vssd1 vccd1 vccd1 _05921_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21959_ net184 net2658 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _07595_ _07650_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__or2_2
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _04821_ net2726 net2789 _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a22o_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ net11 net10 vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__and2_2
X_15480_ net3148 _08297_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__nor2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _07572_ _07580_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__or2_1
X_11643_ net3760 _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ _09732_ _09733_ vssd1 vssd1 vccd1 vccd1 _10152_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14362_ _07444_ _07509_ _07512_ net7757 vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__o211a_1
X_11574_ _04686_ _04684_ _04685_ _04645_ _04683_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a311o_1
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
X_16101_ _08994_ _09175_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__or2_1
Xinput28 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_4
Xinput39 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
X_13313_ _06446_ _06450_ _06451_ _06462_ _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a221o_1
X_17081_ net3578 net4334 vssd1 vssd1 vccd1 vccd1 _10083_ sky130_fd_sc_hd__or2_1
X_14293_ _06990_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__clkbuf_4
X_16032_ _09103_ _08874_ _09106_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__or3_2
X_13244_ net5706 _06394_ _06393_ _06398_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13175_ _06273_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__04009_ clknet_0__04009_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04009_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12126_ _05207_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__nor2_1
X_17983_ _01920_ _01930_ _01928_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19722_ net3096 _03393_ net1807 _03400_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__o211a_1
X_12057_ _05224_ _05225_ _05002_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__mux2_1
X_16934_ _06221_ _09295_ _09951_ vssd1 vssd1 vccd1 vccd1 _09952_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_205_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11008_ net2326 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__clkbuf_1
X_19653_ net6630 _03362_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__or2_1
X_16865_ _04777_ net3989 net4054 _04162_ vssd1 vssd1 vccd1 vccd1 _09926_ sky130_fd_sc_hd__a31o_1
X_20697__132 clknet_1_1__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__inv_2
X_18604_ _02579_ net4668 _02606_ net3603 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a31o_1
X_15816_ _08387_ _08432_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19584_ _02501_ net797 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or2_4
X_16796_ _09732_ _09733_ _08584_ vssd1 vssd1 vccd1 vccd1 _09866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18535_ _02550_ net6238 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__or2b_1
X_15747_ _08817_ _08821_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _06113_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18466_ net43 _02488_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__and2_1
X_15678_ _08548_ net4954 _08664_ _08540_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__or4b_2
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17417_ _09593_ _10416_ vssd1 vssd1 vccd1 vccd1 _10417_ sky130_fd_sc_hd__nor2_1
X_14629_ _07771_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__a21o_1
X_18397_ _02419_ _02427_ _02425_ _02426_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ _09091_ _09666_ vssd1 vssd1 vccd1 vccd1 _10348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03986_ clknet_0__03986_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03986_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ _09582_ _09477_ _10157_ vssd1 vssd1 vccd1 vccd1 _10280_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19018_ net5619 _02982_ _02985_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4105 net3134 vssd1 vssd1 vccd1 vccd1 net4629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4116 rbzero.debug_overlay.vplaneY\[-7\] vssd1 vssd1 vccd1 vccd1 net4640 sky130_fd_sc_hd__buf_2
XFILLER_0_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4127 net2777 vssd1 vssd1 vccd1 vccd1 net4651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4138 _02877_ vssd1 vssd1 vccd1 vccd1 net4662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3404 _00952_ vssd1 vssd1 vccd1 vccd1 net3928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4149 _03387_ vssd1 vssd1 vccd1 vccd1 net4673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3415 rbzero.spi_registers.spi_buffer\[4\] vssd1 vssd1 vccd1 vccd1 net3939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3426 _02994_ vssd1 vssd1 vccd1 vccd1 net3950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3437 _03464_ vssd1 vssd1 vccd1 vccd1 net3961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3448 _03459_ vssd1 vssd1 vccd1 vccd1 net3972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2703 _03656_ vssd1 vssd1 vccd1 vccd1 net3227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2714 net6085 vssd1 vssd1 vccd1 vccd1 net3238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3459 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 net3983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2725 net6175 vssd1 vssd1 vccd1 vccd1 net3249 sky130_fd_sc_hd__buf_1
Xhold2736 _03919_ vssd1 vssd1 vccd1 vccd1 net3260 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2747 _01175_ vssd1 vssd1 vccd1 vccd1 net3271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _00597_ vssd1 vssd1 vccd1 vccd1 net3282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2769 _03831_ vssd1 vssd1 vccd1 vccd1 net3293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21813_ clknet_leaf_10_i_clk net6215 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21744_ clknet_leaf_1_i_clk net617 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xwire85 net86 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
X_20339__72 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21675_ clknet_leaf_14_i_clk net5373 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdy\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20354__86 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__inv_2
XFILLER_0_4_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20626_ net4023 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20557_ _03902_ net3477 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6030 gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 net6554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6041 _04191_ vssd1 vssd1 vccd1 vccd1 net6565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6052 net1642 vssd1 vssd1 vccd1 vccd1 net6576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ _04403_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__clkbuf_4
X_20488_ net3777 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__clkbuf_1
Xhold6063 rbzero.spi_registers.buf_texadd1\[13\] vssd1 vssd1 vccd1 vccd1 net6587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6074 net1620 vssd1 vssd1 vccd1 vccd1 net6598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6085 rbzero.tex_g0\[37\] vssd1 vssd1 vccd1 vccd1 net6609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5340 net2353 vssd1 vssd1 vccd1 vccd1 net5864 sky130_fd_sc_hd__dlygate4sd3_1
X_22227_ net359 net2444 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold6096 net1659 vssd1 vssd1 vccd1 vccd1 net6620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5351 rbzero.map_overlay.i_othery\[3\] vssd1 vssd1 vccd1 vccd1 net5875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5362 net2393 vssd1 vssd1 vccd1 vccd1 net5886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5373 net1780 vssd1 vssd1 vccd1 vccd1 net5897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5384 net2677 vssd1 vssd1 vccd1 vccd1 net5908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4650 net5494 vssd1 vssd1 vccd1 vccd1 net5174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5395 _00672_ vssd1 vssd1 vccd1 vccd1 net5919 sky130_fd_sc_hd__dlygate4sd3_1
X_22158_ net290 net1834 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
Xhold4661 rbzero.spi_registers.buf_mapdy\[4\] vssd1 vssd1 vccd1 vccd1 net5185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4672 rbzero.spi_registers.buf_texadd0\[6\] vssd1 vssd1 vccd1 vccd1 net5196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4683 net1376 vssd1 vssd1 vccd1 vccd1 net5207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21109_ net4143 net4649 vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__nor2_1
Xhold4694 rbzero.pov.spi_buffer\[47\] vssd1 vssd1 vccd1 vccd1 net5218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3960 net7534 vssd1 vssd1 vccd1 vccd1 net4484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3971 _01010_ vssd1 vssd1 vccd1 vccd1 net4495 sky130_fd_sc_hd__dlygate4sd3_1
X_14980_ _08083_ _08122_ _08092_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__mux2_1
X_22089_ clknet_leaf_48_i_clk net4035 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold3982 net7522 vssd1 vssd1 vccd1 vccd1 net4506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3993 net714 vssd1 vssd1 vccd1 vccd1 net4517 sky130_fd_sc_hd__dlygate4sd3_1
X_13931_ _06866_ net567 vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _09103_ _09477_ vssd1 vssd1 vccd1 vccd1 _09721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13862_ _06969_ _06977_ _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15601_ _08673_ _08674_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__or2_1
X_12813_ net23 net24 net25 vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a21oi_1
X_16581_ _09518_ _09520_ _09640_ _09651_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__o31a_4
X_13793_ _06920_ _06938_ _06942_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__a21o_1
X_18320_ net4591 net4382 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15532_ _08152_ _08155_ _08160_ _08575_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__or4_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__and2_2
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18251_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__nand2_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _04646_ _06174_ _08294_ _08537_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05823_ _05836_ net6 vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__mux2_1
X_17202_ _09652_ _09779_ _09907_ _10203_ vssd1 vssd1 vccd1 vccd1 _10204_ sky130_fd_sc_hd__o31a_4
XFILLER_0_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14414_ _07493_ _07563_ _07564_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18182_ _02129_ _02139_ _02137_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11626_ _04614_ _04797_ _04613_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__o21ai_1
X_15394_ net3028 _08381_ _08468_ _06209_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__a211o_1
X_17133_ _10130_ _08708_ _10133_ vssd1 vssd1 vccd1 vccd1 _10135_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14345_ _07440_ _07441_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ _04696_ _04697_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17064_ net3417 net4714 vssd1 vssd1 vccd1 vccd1 _10068_ sky130_fd_sc_hd__nand2_1
Xhold609 _03202_ vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ _07371_ _07409_ _07425_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__and3_1
X_11488_ rbzero.texu_hot\[0\] _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_204_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16015_ _08430_ _08431_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ net4916 _06367_ _06381_ _06382_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ net3578 vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__inv_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _05069_ _05275_ _05277_ _05034_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__o211a_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _01999_ _02014_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__xnor2_1
X_13089_ net4912 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__inv_2
Xhold1309 net5849 vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16917_ net4143 _09941_ _09942_ net6148 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__a22o_1
X_19705_ net1608 _03393_ net1910 _03384_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__o211a_1
X_17897_ _01945_ _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19636_ net5095 net798 _03355_ _03354_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__o211a_1
X_16848_ net3978 vssd1 vssd1 vccd1 vccd1 _09917_ sky130_fd_sc_hd__clkbuf_1
X_19567_ net3050 _03305_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__or2_1
X_16779_ _09847_ _09848_ vssd1 vssd1 vccd1 vccd1 _09849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18518_ _02532_ _02535_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__and2_1
X_19498_ _02491_ _02495_ _03238_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__and3_1
XFILLER_0_201_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18449_ _02474_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21460_ clknet_leaf_30_i_clk net3951 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20751__181 clknet_1_0__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__inv_2
X_20411_ net3390 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21391_ clknet_leaf_52_i_clk _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20273_ net3670 _03756_ _03765_ _03761_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22012_ clknet_leaf_95_i_clk net3431 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3212 net5507 vssd1 vssd1 vccd1 vccd1 net3736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_105_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3223 net7359 vssd1 vssd1 vccd1 vccd1 net3747 sky130_fd_sc_hd__buf_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3234 _03833_ vssd1 vssd1 vccd1 vccd1 net3758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3245 net7335 vssd1 vssd1 vccd1 vccd1 net3769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2500 net6081 vssd1 vssd1 vccd1 vccd1 net3024 sky130_fd_sc_hd__clkbuf_2
Xhold2511 net6310 vssd1 vssd1 vccd1 vccd1 net3035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3256 net3691 vssd1 vssd1 vccd1 vccd1 net3780 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2522 net7480 vssd1 vssd1 vccd1 vccd1 net3046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3267 net6138 vssd1 vssd1 vccd1 vccd1 net3791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 net4352 vssd1 vssd1 vccd1 vccd1 net3057 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3278 _03899_ vssd1 vssd1 vccd1 vccd1 net3802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3289 _03925_ vssd1 vssd1 vccd1 vccd1 net3813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2544 net6280 vssd1 vssd1 vccd1 vccd1 net3068 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1810 net6903 vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 _03255_ vssd1 vssd1 vccd1 vccd1 net3079 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1821 _01555_ vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2566 rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 net3090 sky130_fd_sc_hd__clkbuf_2
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2577 _00643_ vssd1 vssd1 vccd1 vccd1 net3101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1832 _00923_ vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1843 net2337 vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2588 net2088 vssd1 vssd1 vccd1 vccd1 net3112 sky130_fd_sc_hd__clkbuf_4
Xhold1854 _01478_ vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2599 net3932 vssd1 vssd1 vccd1 vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1865 net4825 vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1876 _04555_ vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1887 rbzero.tex_b1\[23\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1898 _04269_ vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10790_ net6465 net2304 _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20834__256 clknet_1_1__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__inv_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21727_ clknet_leaf_2_i_clk net6106 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _05457_ vssd1 vssd1 vccd1 vccd1 _05626_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21658_ clknet_leaf_15_i_clk net5126 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_othery\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11411_ net2794 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12391_ _05177_ _05555_ _05557_ _05461_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20609_ _04162_ _04601_ net2987 _09924_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or4b_1
X_21589_ clknet_leaf_23_i_clk net5635 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xtop_ew_algofoogle_95 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_95/HI o_rgb[5] sky130_fd_sc_hd__conb_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ net2582 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
X_14130_ _06895_ _06858_ _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11273_ net2654 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
X_14061_ _07201_ _07208_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__and2_1
Xhold5170 _01087_ vssd1 vssd1 vccd1 vccd1 net5694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5181 rbzero.wall_tracer.mapY\[7\] vssd1 vssd1 vccd1 vccd1 net5705 sky130_fd_sc_hd__dlygate4sd3_1
X_13012_ _06158_ _06162_ _06163_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__or4_1
Xhold5192 net1586 vssd1 vssd1 vccd1 vccd1 net5716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4480 _00795_ vssd1 vssd1 vccd1 vccd1 net5004 sky130_fd_sc_hd__dlygate4sd3_1
X_17820_ _06204_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__buf_4
Xhold4491 _00846_ vssd1 vssd1 vccd1 vccd1 net5015 sky130_fd_sc_hd__dlygate4sd3_1
X_17751_ _08329_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__buf_2
Xhold3790 net7791 vssd1 vssd1 vccd1 vccd1 net4314 sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ _08107_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16702_ _09771_ _09772_ vssd1 vssd1 vccd1 vccd1 _09773_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__03989_ clknet_0__03989_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03989_
+ sky130_fd_sc_hd__clkbuf_16
X_13914_ net566 _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__or2b_1
X_17682_ _10471_ _10561_ _01733_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a21oi_1
X_14894_ _06678_ _08041_ _08043_ vssd1 vssd1 vccd1 vccd1 _08044_ sky130_fd_sc_hd__a21o_1
X_19421_ _03084_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__clkbuf_4
X_16633_ _08498_ _08565_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13845_ _06971_ _06976_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__and2b_1
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19352_ _03084_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__buf_2
X_16564_ _09634_ _09635_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ _06925_ _06915_ _06920_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__nand3_1
X_10988_ net6768 net6986 _04366_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18303_ _02334_ _02342_ _02340_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15515_ _08586_ _08589_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _05882_ _05883_ _05885_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a211o_2
XFILLER_0_85_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19283_ _03039_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__buf_2
X_16495_ _09564_ _09566_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__nand2_1
X_20318__53 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
XFILLER_0_155_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18234_ _02276_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__xnor2_1
X_15446_ _08515_ _08519_ _08520_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__o21a_1
X_12658_ net5 net6 net7 vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18165_ _02210_ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__xnor2_1
X_11609_ _04724_ _04663_ _04778_ _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a31o_1
X_15377_ _08074_ net7773 _08295_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__mux2_1
X_12589_ _05019_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14328_ _07367_ net558 vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18096_ _02142_ _02143_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__nor2_1
Xhold406 net636 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold417 net7629 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold428 net4444 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17047_ _10051_ _10052_ vssd1 vssd1 vccd1 vccd1 _10053_ sky130_fd_sc_hd__or2b_1
Xhold439 net5361 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14259_ net569 _07370_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ net3889 _02966_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or2_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _01567_ vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 net6573 vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1128 net6601 vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ _08849_ _09784_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__nor2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 _00930_ vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19619_ net5350 net799 net911 _03343_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__o211a_1
X_20891_ clknet_1_1__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__buf_1
XFILLER_0_177_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21512_ clknet_leaf_35_i_clk net1313 vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21443_ clknet_leaf_88_i_clk net3137 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21374_ clknet_leaf_61_i_clk _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold940 net6515 vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold951 net5645 vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 net6595 vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 net6534 vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
X_20256_ net3488 _03743_ _03755_ _03748_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__o211a_1
Xhold984 net4867 vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 _04460_ vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3020 _03621_ vssd1 vssd1 vccd1 vccd1 net3544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3031 net4598 vssd1 vssd1 vccd1 vccd1 net3555 sky130_fd_sc_hd__buf_1
Xhold3042 net4596 vssd1 vssd1 vccd1 vccd1 net3566 sky130_fd_sc_hd__buf_1
Xhold3053 net7558 vssd1 vssd1 vccd1 vccd1 net3577 sky130_fd_sc_hd__dlygate4sd3_1
X_20187_ net5175 _03704_ _03716_ _03709_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3064 _01183_ vssd1 vssd1 vccd1 vccd1 net3588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2330 rbzero.tex_r1\[26\] vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3075 _03905_ vssd1 vssd1 vccd1 vccd1 net3599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3086 rbzero.pov.ready_buffer\[47\] vssd1 vssd1 vccd1 vccd1 net3610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2341 net5960 vssd1 vssd1 vccd1 vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2352 net7285 vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3097 _06215_ vssd1 vssd1 vccd1 vccd1 net3621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2363 net7678 vssd1 vssd1 vccd1 vccd1 net2887 sky130_fd_sc_hd__buf_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2374 _04397_ vssd1 vssd1 vccd1 vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 _04312_ vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2385 net4743 vssd1 vssd1 vccd1 vccd1 net2909 sky130_fd_sc_hd__buf_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1651 _01306_ vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2396 net6242 vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1662 _04495_ vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ net2069 _05128_ net2869 vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a21oi_2
Xhold1673 net2119 vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03774_ clknet_0__03774_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03774_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1684 _01300_ vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ net7075 net2762 _04321_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__mux2_1
Xhold1695 _04410_ vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _05008_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13630_ _06660_ _06751_ _06764_ _06766_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__a221o_2
XFILLER_0_212_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10842_ net6500 net2559 _04288_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13561_ _06650_ _06654_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__nand2_1
X_10773_ net7079 net2848 _04255_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ net2942 _08354_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__or2_1
X_12512_ _05279_ _05675_ _05677_ _05244_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__o211a_1
X_16280_ _08684_ _08565_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__nor2_1
X_13492_ _06565_ _06642_ _06587_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ _04627_ _06207_ _04626_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__and3b_2
X_12443_ net4077 _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15162_ net4714 net7437 _08249_ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__mux2_1
X_12374_ _05483_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__buf_4
XFILLER_0_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ _06668_ _06955_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__nor2_1
X_11325_ net6471 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19970_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__buf_2
X_15093_ net3200 net3184 _08191_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11256_ net2867 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
X_14044_ _06865_ _06955_ _07193_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__o21ai_1
X_18921_ _02890_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11187_ net2545 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
X_18852_ _02835_ _02840_ _04632_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
X_17803_ _10583_ _01731_ _01729_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a21oi_1
X_18783_ net4640 _02768_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__nand2_1
X_15995_ _09042_ _09043_ _09061_ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__or3_1
XFILLER_0_207_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17734_ _01783_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__xor2_1
X_14946_ net7759 vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17665_ _01715_ _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__nor2_1
X_14877_ net4315 _08025_ _08027_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16616_ _09683_ _09685_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__and2_1
X_19404_ net5346 _03211_ _03215_ _03207_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13828_ _06968_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__xor2_2
X_20817__240 clknet_1_1__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__inv_2
XFILLER_0_203_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17596_ _10592_ _10593_ vssd1 vssd1 vccd1 vccd1 _10594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16547_ _09481_ _09497_ _09618_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__a21bo_1
X_19335_ net5724 _03172_ _03176_ _03168_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13759_ _06908_ net575 vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19266_ net5140 _03133_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__or2_1
X_16478_ _09311_ _09133_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__and2b_1
Xhold7319 _06663_ vssd1 vssd1 vccd1 vccd1 net7843 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18217_ _02263_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15429_ _08456_ _08470_ _08484_ _08493_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_54_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6607 net2600 vssd1 vssd1 vccd1 vccd1 net7131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ net2973 net7325 _03084_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6618 rbzero.tex_g0\[45\] vssd1 vssd1 vccd1 vccd1 net7142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6629 net2363 vssd1 vssd1 vccd1 vccd1 net7153 sky130_fd_sc_hd__dlygate4sd3_1
X_18148_ _02189_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__xor2_1
Xhold5906 _04554_ vssd1 vssd1 vccd1 vccd1 net6430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5917 net1267 vssd1 vssd1 vccd1 vccd1 net6441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5928 rbzero.tex_r1\[0\] vssd1 vssd1 vccd1 vccd1 net6452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold203 net6211 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 net7616 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_1
Xhold5939 net1358 vssd1 vssd1 vccd1 vccd1 net6463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18079_ _10257_ net7378 _02125_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a21oi_1
Xhold225 net6214 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 net6336 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold247 net5002 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ net2937 _03667_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__or2_1
Xhold258 net5035 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold269 net5058 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21090_ _04076_ _04079_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__nand2_1
X_20863__282 clknet_1_0__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__inv_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20041_ net3388 _03613_ net4494 _03602_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21992_ net217 net2801 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22475_ clknet_leaf_77_i_clk net661 vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21426_ clknet_leaf_44_i_clk net3806 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21357_ clknet_leaf_41_i_clk net5748 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11110_ net6716 net2717 _04426_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ rbzero.tex_r1\[9\] rbzero.tex_r1\[8\] _05219_ vssd1 vssd1 vccd1 vccd1 _05259_
+ sky130_fd_sc_hd__mux2_1
X_21288_ clknet_leaf_88_i_clk net4097 vssd1 vssd1 vccd1 vccd1 reg_rgb\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold770 net5539 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 net4304 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ net1898 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
Xhold792 net3567 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
X_20239_ net3435 _03743_ _03746_ _03735_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__o211a_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _01464_ vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2171 net7234 vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
X_14800_ _07900_ _07899_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__and2b_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 net5945 vssd1 vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
X_15780_ _08821_ _08839_ _08854_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__nand3_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2193 net7254 vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__nor2_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1470 _01560_ vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1481 _04371_ vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _07843_ net78 vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__xor2_2
XFILLER_0_197_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ net3378 net3218 _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and3_1
Xhold1492 _00936_ vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ _10213_ _10214_ _10323_ vssd1 vssd1 vccd1 vccd1 _10450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14662_ _07810_ _07809_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__and2b_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _05014_ vssd1 vssd1 vccd1 vccd1 _05044_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _09472_ _09473_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__or2b_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ _06752_ _06701_ _06756_ _06763_ _06589_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a221o_1
XFILLER_0_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10825_ net7309 net7262 _04277_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
X_17381_ _10259_ _08329_ _10379_ _10380_ vssd1 vssd1 vccd1 vccd1 _10381_ sky130_fd_sc_hd__or4_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ _06955_ _07353_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19120_ net5375 _03040_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__or2_1
X_16332_ _09403_ net7381 vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13544_ _06694_ _06693_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__nand2_4
X_10756_ net7004 net2101 _04244_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19051_ net2842 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__clkbuf_1
X_16263_ _08394_ _08498_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13475_ net7757 net3237 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__nand2_4
X_10687_ net2855 net7241 _04203_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18002_ _02049_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__nand2_1
X_15214_ _04692_ _08290_ net3509 vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__mux2_1
X_12426_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _05483_ vssd1 vssd1 vccd1 vccd1 _05593_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16194_ _08805_ _08834_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15145_ _08250_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _04975_ _05491_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11308_ net2147 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
X_15076_ rbzero.wall_tracer.visualWallDist\[-9\] _08201_ vssd1 vssd1 vccd1 vccd1 _08202_
+ sky130_fd_sc_hd__or2_1
X_19953_ net3893 _03560_ _03476_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a21o_1
X_12288_ _04987_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__clkbuf_8
X_14027_ _07133_ _07166_ _07176_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__and3_1
X_18904_ _02529_ net4759 net7599 net3445 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__a31o_1
X_11239_ net2413 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
X_19884_ _03511_ _03512_ _03476_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ net4459 net4640 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _09048_ _09050_ _09020_ _09052_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__o2bb2a_1
X_18766_ _05396_ net1091 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17717_ _10586_ _01765_ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__o21a_1
X_14929_ net7891 _08016_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18697_ _02646_ net7146 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__04005_ clknet_0__04005_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04005_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17648_ _09593_ _10539_ _10543_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17579_ _10458_ _10460_ vssd1 vssd1 vccd1 vccd1 _10577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19318_ net794 _03159_ net4215 _03155_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20590_ net3524 net1302 net3250 vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7105 rbzero.wall_tracer.rayAddendY\[-6\] vssd1 vssd1 vccd1 vccd1 net7629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7116 rbzero.wall_tracer.rayAddendY\[-5\] vssd1 vssd1 vccd1 vccd1 net7640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7127 rbzero.floor_leak\[1\] vssd1 vssd1 vccd1 vccd1 net7651 sky130_fd_sc_hd__dlygate4sd3_1
X_19249_ net603 _03120_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7138 rbzero.row_render.texu\[4\] vssd1 vssd1 vccd1 vccd1 net7662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7149 rbzero.spi_registers.texadd3\[14\] vssd1 vssd1 vccd1 vccd1 net7673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6404 net2593 vssd1 vssd1 vccd1 vccd1 net6928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6415 rbzero.tex_g0\[43\] vssd1 vssd1 vccd1 vccd1 net6939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22260_ net392 net1514 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
Xhold6426 net2031 vssd1 vssd1 vccd1 vccd1 net6950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6437 rbzero.tex_g0\[39\] vssd1 vssd1 vccd1 vccd1 net6961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6448 net2285 vssd1 vssd1 vccd1 vccd1 net6972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_182_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5703 net1792 vssd1 vssd1 vccd1 vccd1 net6227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6459 rbzero.tex_b0\[7\] vssd1 vssd1 vccd1 vccd1 net6983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5714 _02551_ vssd1 vssd1 vccd1 vccd1 net6238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21211_ _03502_ net1136 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5725 _06216_ vssd1 vssd1 vccd1 vccd1 net6249 sky130_fd_sc_hd__dlygate4sd3_1
X_22191_ net323 net2404 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5736 _08224_ vssd1 vssd1 vccd1 vccd1 net6260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5747 net1571 vssd1 vssd1 vccd1 vccd1 net6271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5758 _08221_ vssd1 vssd1 vccd1 vccd1 net6282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5769 rbzero.spi_registers.buf_leak\[4\] vssd1 vssd1 vccd1 vccd1 net6293 sky130_fd_sc_hd__dlygate4sd3_1
X_21142_ _04626_ _04818_ net4027 vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o21ai_1
X_21073_ _04018_ _04067_ _04068_ _04017_ net4546 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20024_ net4600 _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21975_ net200 net1499 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer40 _06973_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer51 _06909_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer62 _06884_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ clknet_1_0__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__buf_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ net2686 net51 _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11590_ rbzero.spi_registers.texadd1\[3\] _04644_ _04709_ vssd1 vssd1 vccd1 vccd1
+ _04762_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ _06396_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22458_ clknet_leaf_38_i_clk _01627_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ rbzero.debug_overlay.facingY\[-6\] _05378_ _05379_ rbzero.debug_overlay.facingY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a22o_1
X_21409_ clknet_leaf_79_i_clk net2921 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13191_ net2864 _06190_ net4913 net2536 vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22389_ net521 net2520 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold6982 _00502_ vssd1 vssd1 vccd1 vccd1 net7506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6993 net4252 vssd1 vssd1 vccd1 vccd1 net7517 sky130_fd_sc_hd__dlygate4sd3_1
X_12142_ net4033 _04599_ _04759_ _04831_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ _05068_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__or2_1
X_16950_ net5969 _09294_ vssd1 vssd1 vccd1 vccd1 _09967_ sky130_fd_sc_hd__xor2_1
XFILLER_0_159_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ net2672 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__clkbuf_1
X_15901_ _08902_ _08903_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16881_ net4278 _09934_ _09936_ _08096_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__a22o_1
X_15832_ _08905_ _08898_ _08906_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__nand3_2
X_18620_ net3242 net4476 _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _08823_ _08824_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__xnor2_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _04632_ _02559_ _02560_ _02565_ _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a32o_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ net3876 net3085 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__nand2_2
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _10485_ _10500_ vssd1 vssd1 vccd1 vccd1 _10501_ sky130_fd_sc_hd__xnor2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _07774_ _07354_ _07862_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__or3_1
XFILLER_0_185_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11926_ net3378 _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nand2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _02499_ _02502_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nand2_1
X_15694_ _08425_ _08445_ _08423_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__a21bo_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _10402_ _10432_ vssd1 vssd1 vccd1 vccd1 _10433_ sky130_fd_sc_hd__xnor2_2
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _07763_ _07787_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__xnor2_2
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _04971_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__or2_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10808_ net7290 net6407 _04266_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
X_17364_ _10258_ _10262_ _10362_ vssd1 vssd1 vccd1 vccd1 _10364_ sky130_fd_sc_hd__and3_1
X_14576_ _07700_ _07726_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__and2_2
X_11788_ _04938_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ _09348_ _09388_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19103_ net5367 _03040_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__or2_1
X_13527_ _06677_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__clkbuf_4
X_10739_ net2724 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__clkbuf_1
X_17295_ _10294_ _10295_ vssd1 vssd1 vccd1 vccd1 _10296_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19034_ net3933 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__buf_4
X_16246_ _09203_ _09302_ _09319_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20929__341 clknet_1_0__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__inv_2
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13458_ _06600_ _06603_ _06606_ _06608_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_24_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _05062_ _05571_ _05573_ _05575_ _05030_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a221o_1
X_16177_ _08310_ _09251_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ _06478_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4309 net1209 vssd1 vssd1 vccd1 vccd1 net4833 sky130_fd_sc_hd__dlygate4sd3_1
X_15128_ net6146 _08223_ vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3608 net696 vssd1 vssd1 vccd1 vccd1 net4132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3619 net7637 vssd1 vssd1 vccd1 vccd1 net4143 sky130_fd_sc_hd__dlygate4sd3_1
X_19936_ net4288 _03532_ net1019 _03519_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__a211o_1
X_15059_ net4332 _08188_ _08026_ vssd1 vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__mux2_1
Xhold2907 _01181_ vssd1 vssd1 vccd1 vccd1 net3431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2918 _03879_ vssd1 vssd1 vccd1 vccd1 net3442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2929 rbzero.pov.ready_buffer\[15\] vssd1 vssd1 vccd1 vccd1 net3453 sky130_fd_sc_hd__dlygate4sd3_1
X_19867_ _03478_ net3000 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18818_ _05396_ _02787_ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19798_ net6060 _03443_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__or2_1
X_20975__383 clknet_1_0__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__inv_2
X_18749_ net4821 _06396_ _06198_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20674__111 clknet_1_1__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__inv_2
XFILLER_0_204_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21760_ clknet_leaf_23_i_clk net1873 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21691_ clknet_leaf_26_i_clk net5203 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20642_ _03083_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20573_ _03924_ net3753 vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6201 _04548_ vssd1 vssd1 vccd1 vccd1 net6725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22312_ net444 net1779 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6212 net1856 vssd1 vssd1 vccd1 vccd1 net6736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6223 _04557_ vssd1 vssd1 vccd1 vccd1 net6747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6234 net1880 vssd1 vssd1 vccd1 vccd1 net6758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6245 rbzero.tex_g0\[29\] vssd1 vssd1 vccd1 vccd1 net6769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5500 gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 net6024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5511 net2875 vssd1 vssd1 vccd1 vccd1 net6035 sky130_fd_sc_hd__dlygate4sd3_1
X_22243_ net375 net1203 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold6256 net2104 vssd1 vssd1 vccd1 vccd1 net6780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6267 rbzero.tex_g0\[7\] vssd1 vssd1 vccd1 vccd1 net6791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5522 rbzero.spi_registers.spi_buffer\[22\] vssd1 vssd1 vccd1 vccd1 net6046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6278 net1897 vssd1 vssd1 vccd1 vccd1 net6802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5533 rbzero.spi_registers.spi_buffer\[16\] vssd1 vssd1 vccd1 vccd1 net6057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6289 rbzero.tex_b1\[52\] vssd1 vssd1 vccd1 vccd1 net6813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5544 _02842_ vssd1 vssd1 vccd1 vccd1 net6068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4810 net872 vssd1 vssd1 vccd1 vccd1 net5334 sky130_fd_sc_hd__buf_1
XFILLER_0_30_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5555 _02568_ vssd1 vssd1 vccd1 vccd1 net6079 sky130_fd_sc_hd__dlygate4sd3_1
X_22174_ net306 net1890 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold4821 rbzero.spi_registers.texadd3\[5\] vssd1 vssd1 vccd1 vccd1 net5345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4832 net947 vssd1 vssd1 vccd1 vccd1 net5356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5577 _02876_ vssd1 vssd1 vccd1 vccd1 net6101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4843 net981 vssd1 vssd1 vccd1 vccd1 net5367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5588 rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 net6112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4854 rbzero.traced_texa\[-7\] vssd1 vssd1 vccd1 vccd1 net5378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5599 net4524 vssd1 vssd1 vccd1 vccd1 net6123 sky130_fd_sc_hd__clkbuf_4
X_21125_ net4744 _04017_ _04014_ _04112_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a22o_1
Xhold4865 net1319 vssd1 vssd1 vccd1 vccd1 net5389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4876 net1057 vssd1 vssd1 vccd1 vccd1 net5400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4887 _01043_ vssd1 vssd1 vccd1 vccd1 net5411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4898 net978 vssd1 vssd1 vccd1 vccd1 net5422 sky130_fd_sc_hd__dlygate4sd3_1
X_21056_ net4146 net4736 vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_1
X_20007_ _03261_ net3830 vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ net18 _05899_ _05919_ net20 vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a22o_1
X_21958_ net183 net2513 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ net4059 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__inv_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ net11 net10 vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_167_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21889_ clknet_leaf_96_i_clk net1289 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _07572_ _07580_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11642_ net6025 net3989 vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14361_ _07491_ _07510_ _07511_ _07450_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ _04677_ _04650_ _04675_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and3_1
X_16100_ _09036_ _08997_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__nor2_1
Xinput18 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XFILLER_0_18_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__and2_1
Xinput29 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_4
X_17080_ _10082_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__clkbuf_1
X_14292_ _07404_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16031_ _09084_ _09104_ _09105_ vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _06395_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6790 rbzero.spi_registers.spi_cmd\[2\] vssd1 vssd1 vccd1 vccd1 net7314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ _06272_ net3852 _06282_ _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__04008_ clknet_0__04008_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04008_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _05255_ _05293_ _04975_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _02029_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__nor2_1
X_19721_ net6256 _03395_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__or2_1
X_12056_ rbzero.tex_r1\[59\] rbzero.tex_r1\[58\] _05077_ vssd1 vssd1 vccd1 vccd1 _05225_
+ sky130_fd_sc_hd__mux2_1
X_16933_ _06217_ _09950_ vssd1 vssd1 vccd1 vccd1 _09951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11007_ net6778 net7145 _04377_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux2_1
X_19652_ _02998_ _03360_ net1668 _03354_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__o211a_1
X_16864_ _04162_ _04812_ net4054 vssd1 vssd1 vccd1 vccd1 _09925_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _02613_ _02614_ rbzero.wall_tracer.rayAddendX\[1\] _09932_ vssd1 vssd1 vccd1
+ vccd1 _02615_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_205_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15815_ _08886_ _08889_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__xnor2_2
X_16795_ _09863_ _09864_ _08626_ vssd1 vssd1 vccd1 vccd1 _09865_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19583_ net798 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15746_ _08817_ _08818_ _08820_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__nand3_1
XFILLER_0_158_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18534_ net6237 net2919 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _05077_ vssd1 vssd1 vccd1 vccd1 _05079_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ _08667_ _08668_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__xnor2_2
X_18465_ _08274_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__buf_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ net34 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__clkbuf_4
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17416_ _10415_ vssd1 vssd1 vccd1 vccd1 _10416_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14628_ _07772_ _07777_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__and2b_1
X_18396_ _02425_ _02426_ _02419_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17347_ _10345_ _10346_ vssd1 vssd1 vccd1 vccd1 _10347_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14559_ _07705_ _07708_ _07709_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__a21boi_2
Xclkbuf_1_1__f__03985_ clknet_0__03985_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03985_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17278_ _10254_ _10278_ vssd1 vssd1 vccd1 vccd1 _10279_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16229_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__or2b_1
X_19017_ net5619 _02982_ _02967_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4117 _03639_ vssd1 vssd1 vccd1 vccd1 net4641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4128 rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 net4652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4139 _02892_ vssd1 vssd1 vccd1 vccd1 net4663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3405 net6040 vssd1 vssd1 vccd1 vccd1 net3929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3416 net3104 vssd1 vssd1 vccd1 vccd1 net3940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3427 _00629_ vssd1 vssd1 vccd1 vccd1 net3951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3438 _03465_ vssd1 vssd1 vccd1 vccd1 net3962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3449 _03462_ vssd1 vssd1 vccd1 vccd1 net3973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2704 _01029_ vssd1 vssd1 vccd1 vccd1 net3228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2715 _00580_ vssd1 vssd1 vccd1 vccd1 net3239 sky130_fd_sc_hd__dlygate4sd3_1
X_19919_ net3611 _03477_ _03532_ _03540_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a211o_1
Xhold2726 _03800_ vssd1 vssd1 vccd1 vccd1 net3250 sky130_fd_sc_hd__buf_4
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2737 _01236_ vssd1 vssd1 vccd1 vccd1 net3261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2748 net7372 vssd1 vssd1 vccd1 vccd1 net3272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2759 net4926 vssd1 vssd1 vccd1 vccd1 net3283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21812_ clknet_leaf_10_i_clk net4389 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21743_ clknet_leaf_1_i_clk net4238 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xwire86 _05442_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21674_ clknet_leaf_14_i_clk net808 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdy\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20625_ _02992_ _03962_ net4022 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__and3_1
XFILLER_0_191_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20556_ net1156 net3476 _03911_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6020 _04394_ vssd1 vssd1 vccd1 vccd1 net6544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6031 net1920 vssd1 vssd1 vccd1 vccd1 net6555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6042 net1629 vssd1 vssd1 vccd1 vccd1 net6566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6053 rbzero.tex_r0\[39\] vssd1 vssd1 vccd1 vccd1 net6577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20487_ _03858_ net3776 vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__and2_1
Xhold6064 net1692 vssd1 vssd1 vccd1 vccd1 net6588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5330 rbzero.tex_g1\[32\] vssd1 vssd1 vccd1 vccd1 net5854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6075 _04588_ vssd1 vssd1 vccd1 vccd1 net6599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5341 rbzero.tex_b1\[28\] vssd1 vssd1 vccd1 vccd1 net5865 sky130_fd_sc_hd__dlygate4sd3_1
X_22226_ net358 net1503 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold6086 net1877 vssd1 vssd1 vccd1 vccd1 net6610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6097 rbzero.spi_registers.buf_texadd1\[18\] vssd1 vssd1 vccd1 vccd1 net6621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5352 net2536 vssd1 vssd1 vccd1 vccd1 net5876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5363 _04237_ vssd1 vssd1 vccd1 vccd1 net5887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5374 _04350_ vssd1 vssd1 vccd1 vccd1 net5898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4640 rbzero.spi_registers.texadd0\[17\] vssd1 vssd1 vccd1 vccd1 net5164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5385 _00655_ vssd1 vssd1 vccd1 vccd1 net5909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4651 net1470 vssd1 vssd1 vccd1 vccd1 net5175 sky130_fd_sc_hd__dlygate4sd3_1
X_22157_ net289 net2142 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold5396 rbzero.tex_g0\[1\] vssd1 vssd1 vccd1 vccd1 net5920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4662 net882 vssd1 vssd1 vccd1 vccd1 net5186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4673 net809 vssd1 vssd1 vccd1 vccd1 net5197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4684 rbzero.pov.spi_buffer\[9\] vssd1 vssd1 vccd1 vccd1 net5208 sky130_fd_sc_hd__dlygate4sd3_1
X_21108_ _04093_ _04095_ _04094_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a21boi_1
Xhold3950 net7459 vssd1 vssd1 vccd1 vccd1 net4474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4695 net1324 vssd1 vssd1 vccd1 vccd1 net5219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3961 net3284 vssd1 vssd1 vccd1 vccd1 net4485 sky130_fd_sc_hd__dlygate4sd3_1
X_22088_ clknet_leaf_49_i_clk net3899 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold3972 net7453 vssd1 vssd1 vccd1 vccd1 net4496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3983 net3447 vssd1 vssd1 vccd1 vccd1 net4507 sky130_fd_sc_hd__buf_1
XFILLER_0_195_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3994 net7753 vssd1 vssd1 vccd1 vccd1 net4518 sky130_fd_sc_hd__dlygate4sd3_1
X_13930_ net557 _07072_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__o21ai_2
X_21039_ net985 net5424 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _06978_ _06968_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15600_ _08673_ _08674_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12812_ net4060 _05957_ _05958_ _05194_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__a221o_1
X_16580_ _09530_ _09516_ _09639_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__a21o_1
X_13792_ _06920_ _06938_ _06942_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__nand3_1
X_15531_ _08604_ _08591_ _08534_ _08605_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__a31o_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__nor2b_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _01802_ _09732_ _02182_ _02186_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__o31a_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_91_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _08300_ _06470_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__nand2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12674_ net8 _05832_ _05835_ _05821_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _09782_ _09780_ _09906_ vssd1 vssd1 vccd1 vccd1 _10203_ sky130_fd_sc_hd__a21o_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _07467_ _07500_ _07494_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__and3_1
X_18181_ _02217_ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _04727_ _04718_ _04794_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__o31a_1
X_20811__235 clknet_1_1__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__inv_2
XFILLER_0_167_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15393_ _08381_ _08467_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17132_ _10130_ _08708_ _10133_ vssd1 vssd1 vccd1 vccd1 _10134_ sky130_fd_sc_hd__or3_1
XFILLER_0_170_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ _07490_ _07494_ net7438 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__a21o_1
X_11556_ _04717_ _04721_ _04723_ _04725_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17063_ net3417 net4714 vssd1 vssd1 vccd1 vccd1 _10067_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14275_ _07371_ _07409_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__a21oi_1
X_11487_ rbzero.spi_registers.texadd3\[6\] rbzero.spi_registers.texadd1\[6\] rbzero.spi_registers.texadd0\[6\]
+ rbzero.spi_registers.texadd2\[6\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__mux4_1
X_16014_ _09084_ _09088_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__xnor2_1
X_13226_ _06257_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _06312_ net3200 _06309_ net3221 vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a2bb2o_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _05002_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or2_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17965_ _02012_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nor2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13088_ _06186_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__inv_2
X_19704_ net6568 _03395_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ net3014 _05103_ _05115_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a21oi_1
X_16916_ net4186 _09941_ _09942_ net6098 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17896_ _01833_ _01837_ _01944_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__and3_1
X_20892__307 clknet_1_0__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_44_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19635_ net2948 _03326_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__or2_1
X_16847_ _04760_ _04812_ _04852_ net3977 vssd1 vssd1 vccd1 vccd1 _09916_ sky130_fd_sc_hd__and4_1
X_19566_ net5216 _03303_ _03315_ _03314_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__o211a_1
X_16778_ _09831_ _09832_ _09846_ vssd1 vssd1 vccd1 vccd1 _09848_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18517_ net4425 net4657 _02532_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__nand3b_1
X_15729_ _08802_ _08803_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__nor2_2
X_19497_ net1727 _03265_ net5784 _03260_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18448_ _02473_ net4437 _02411_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18379_ net4429 net4451 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20410_ _03814_ net3389 vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__and2_1
X_20786__212 clknet_1_1__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__inv_2
X_21390_ clknet_leaf_53_i_clk _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03999_ _03999_ vssd1 vssd1 vccd1 vccd1 clknet_0__03999_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20272_ net3752 net4839 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22011_ clknet_leaf_98_i_clk net3192 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3202 net6119 vssd1 vssd1 vccd1 vccd1 net3726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3213 net1243 vssd1 vssd1 vccd1 vccd1 net3737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3224 _02968_ vssd1 vssd1 vccd1 vccd1 net3748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3235 _01197_ vssd1 vssd1 vccd1 vccd1 net3759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3246 _03612_ vssd1 vssd1 vccd1 vccd1 net3770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2501 _09285_ vssd1 vssd1 vccd1 vccd1 net3025 sky130_fd_sc_hd__buf_1
XFILLER_0_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2512 _00598_ vssd1 vssd1 vccd1 vccd1 net3036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3257 rbzero.pov.spi_buffer\[30\] vssd1 vssd1 vccd1 vccd1 net3781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3268 _00415_ vssd1 vssd1 vccd1 vccd1 net3792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 net7547 vssd1 vssd1 vccd1 vccd1 net3047 sky130_fd_sc_hd__buf_1
Xhold3279 _01227_ vssd1 vssd1 vccd1 vccd1 net3803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2534 net3741 vssd1 vssd1 vccd1 vccd1 net3058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1800 _01316_ vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2545 rbzero.spi_registers.spi_buffer\[14\] vssd1 vssd1 vccd1 vccd1 net3069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 _04326_ vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2556 _00809_ vssd1 vssd1 vccd1 vccd1 net3080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1822 net7134 vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2567 _02918_ vssd1 vssd1 vccd1 vccd1 net3091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1833 net7051 vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2578 net7795 vssd1 vssd1 vccd1 vccd1 net3102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _04245_ vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2589 _00634_ vssd1 vssd1 vccd1 vccd1 net3113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1855 net7005 vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1866 net6727 vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1877 _01148_ vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1888 net2179 vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1899 _01500_ vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21726_ clknet_leaf_2_i_clk net1731 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21657_ clknet_leaf_15_i_clk net5408 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_othery\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ net7264 net6798 _04584_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20608_ net4103 net6266 net4015 _03947_ _08276_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__o221a_1
X_12390_ _05019_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__or2_1
X_21588_ clknet_leaf_23_i_clk net5654 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_96 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_96/HI o_rgb[8] sky130_fd_sc_hd__conb_1
X_11341_ net6888 net6746 _04551_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20539_ net3288 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ _07196_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__xnor2_1
X_11272_ net6337 net7002 _04514_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5160 net3063 vssd1 vssd1 vccd1 vccd1 net5684 sky130_fd_sc_hd__buf_1
XFILLER_0_120_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13011_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\] _06165_
+ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__or4_1
X_22209_ net341 net2664 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
Xhold5171 rbzero.pov.ready_buffer\[21\] vssd1 vssd1 vccd1 vccd1 net5695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5182 net2768 vssd1 vssd1 vccd1 vccd1 net5706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5193 rbzero.spi_registers.buf_texadd2\[15\] vssd1 vssd1 vccd1 vccd1 net5717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4470 rbzero.spi_registers.texadd1\[8\] vssd1 vssd1 vccd1 vccd1 net4994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4481 net772 vssd1 vssd1 vccd1 vccd1 net5005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4492 net756 vssd1 vssd1 vccd1 vccd1 net5016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3780 _00496_ vssd1 vssd1 vccd1 vccd1 net4304 sky130_fd_sc_hd__dlygate4sd3_1
X_17750_ _10259_ _09231_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__or2_1
X_14962_ net4473 _08106_ _08027_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__mux2_1
Xhold3791 net3017 vssd1 vssd1 vccd1 vccd1 net4315 sky130_fd_sc_hd__buf_1
Xclkbuf_1_0__f__03988_ clknet_0__03988_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03988_
+ sky130_fd_sc_hd__clkbuf_16
X_16701_ _09769_ net3029 vssd1 vssd1 vccd1 vccd1 _09772_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13913_ _07041_ _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__and2_4
X_17681_ _10558_ _10560_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14893_ _08006_ _08042_ _06838_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__a21o_1
X_19420_ _03035_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__clkbuf_4
X_16632_ _09701_ _09702_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__and2_1
X_13844_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__xor2_1
XFILLER_0_187_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19351_ _03035_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__clkbuf_4
X_16563_ _09631_ _09633_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13775_ _06915_ _06920_ _06925_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10987_ net6638 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__clkbuf_1
X_18302_ _02345_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__clkbuf_1
X_15514_ _08587_ _08588_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__nor2_1
X_12726_ _05853_ _05886_ _05845_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16494_ _09565_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19282_ _03036_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ _08516_ _08501_ _08518_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__or3_1
X_18233_ _02277_ _02278_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12657_ _05816_ _05795_ _05799_ net4060 _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11608_ _04159_ _04660_ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18164_ _09486_ _10379_ net8017 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__or3b_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15376_ _06165_ _06418_ net4086 vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__mux2_1
X_12588_ rbzero.tex_b1\[3\] rbzero.tex_b1\[2\] _05483_ vssd1 vssd1 vccd1 vccd1 _05753_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17115_ _09809_ _09819_ _09817_ vssd1 vssd1 vccd1 vccd1 _10117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14327_ _07477_ _07476_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18095_ _02140_ _02141_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11539_ _04680_ _04708_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold407 net7316 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 net4803 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ net3462 net4716 vssd1 vssd1 vccd1 vccd1 _10052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14258_ _07373_ _07384_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__or2b_1
Xhold429 net5597 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ _06222_ _06186_ _06183_ _06196_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__and4_1
X_14189_ _07279_ _07284_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__nand2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ net3889 _02966_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__and2_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 net6110 vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 net6575 vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ _01995_ _01996_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__nand2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 _03364_ vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
X_17879_ _01925_ _01927_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19618_ net910 _03340_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19549_ net5132 _03303_ _03306_ _03295_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21511_ clknet_leaf_44_i_clk net1055 vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21442_ clknet_leaf_86_i_clk net4820 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21373_ clknet_leaf_62_i_clk _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold930 net6454 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 net6517 vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold952 net5647 vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _01321_ vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
X_20255_ net5588 _03744_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__or2_1
Xhold974 net6536 vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3010 net4025 vssd1 vssd1 vccd1 vccd1 net3534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 net4869 vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 _01328_ vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3021 _03622_ vssd1 vssd1 vccd1 vccd1 net3545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3032 rbzero.pov.spi_buffer\[27\] vssd1 vssd1 vccd1 vccd1 net3556 sky130_fd_sc_hd__dlygate4sd3_1
X_20186_ net3651 _03705_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or2_1
Xhold3043 net5790 vssd1 vssd1 vccd1 vccd1 net3567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3054 net3186 vssd1 vssd1 vccd1 vccd1 net3578 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3065 net5611 vssd1 vssd1 vccd1 vccd1 net3589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2320 _00644_ vssd1 vssd1 vccd1 vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2331 net2778 vssd1 vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
X_20840__261 clknet_1_0__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__inv_2
Xhold3076 _03906_ vssd1 vssd1 vccd1 vccd1 net3600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2342 net7252 vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3087 net2922 vssd1 vssd1 vccd1 vccd1 net3611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2353 _04374_ vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3098 _06258_ vssd1 vssd1 vccd1 vccd1 net3622 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2364 net4602 vssd1 vssd1 vccd1 vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2375 _01384_ vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1630 _01559_ vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 _01461_ vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 net4745 vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1652 net5903 vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2397 _00578_ vssd1 vssd1 vccd1 vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1663 _01296_ vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1674 _04498_ vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03773_ clknet_0__03773_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03773_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1685 net6929 vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
X_10910_ net7231 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1696 _01373_ vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _05058_ _05059_ _04984_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__mux2_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ net2377 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xsplit34 _07464_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _06657_ _06702_ _06706_ _06710_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a31o_1
X_10772_ net6654 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ _05229_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21709_ clknet_leaf_19_i_clk net1654 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _06633_ _06637_ _06640_ _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ net788 net7327 _05120_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15161_ _08258_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__clkbuf_1
X_12373_ _05261_ _05537_ _05539_ _05244_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14112_ _06995_ _07006_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__nand2_1
X_11324_ net6469 net1753 _04540_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _08190_ net3463 net6204 _01622_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__o211a_1
X_14043_ _06864_ _07193_ _06970_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__or3_1
X_18920_ _02863_ net3090 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__or2_1
X_11255_ net6938 net7253 _04503_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_1
X_20923__336 clknet_1_0__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__inv_2
X_18851_ _02824_ _02839_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__xnor2_1
X_11186_ net6842 net7215 _04470_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17802_ _01762_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__xnor2_1
X_18782_ net2885 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__clkbuf_1
X_15994_ _09067_ _09068_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17733_ _10383_ _09312_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__nor2_1
X_14945_ _06664_ _08089_ _08090_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_203_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _10301_ _01710_ _01714_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__and3_1
X_14876_ _08026_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__buf_4
X_19403_ net1661 _03212_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__or2_1
X_16615_ _09683_ _09685_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_212_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13827_ _06969_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__xnor2_2
X_17595_ _10590_ _10591_ vssd1 vssd1 vccd1 vccd1 _10593_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19334_ net1548 _03173_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or2_1
X_16546_ _09496_ _09492_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13758_ _06892_ _06901_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12709_ _04760_ _04603_ _04637_ _04165_ net10 net11 vssd1 vssd1 vccd1 vccd1 _05870_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_183_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19265_ net5165 _03132_ _03136_ _03128_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__o211a_1
X_16477_ _09545_ _09546_ _09548_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__o21a_1
X_13689_ _06759_ _06753_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__nor2_1
Xhold7309 rbzero.wall_tracer.stepDistY\[4\] vssd1 vssd1 vccd1 vccd1 net7833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ _02262_ net3780 _01749_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_2
X_15428_ _08455_ _08470_ _08483_ _08493_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__or4_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19196_ net5330 _03078_ _03095_ _03096_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__o211a_1
Xhold6608 rbzero.tex_g1\[23\] vssd1 vssd1 vccd1 vccd1 net7132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6619 net2538 vssd1 vssd1 vccd1 vccd1 net7143 sky130_fd_sc_hd__dlygate4sd3_1
X_18147_ _02192_ _02193_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__xnor2_2
X_15359_ net4063 _08412_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__or2_1
Xhold5907 net1197 vssd1 vssd1 vccd1 vccd1 net6431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5918 _04466_ vssd1 vssd1 vccd1 vccd1 net6442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5929 net1453 vssd1 vssd1 vccd1 vccd1 net6453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 net6332 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold215 net4623 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold226 rbzero.tex_g0\[2\] vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _10257_ net7378 _02125_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__and3_1
Xhold237 net6338 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold248 net5004 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _10019_ _09276_ vssd1 vssd1 vccd1 vccd1 _10037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold259 net5037 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ net4493 _03614_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20898__313 clknet_1_1__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__inv_2
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21991_ net216 net1817 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20870__287 clknet_1_1__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__inv_2
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22474_ clknet_leaf_80_i_clk net4804 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21425_ clknet_leaf_43_i_clk net3884 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21356_ clknet_leaf_42_i_clk net4924 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold760 net5382 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
X_21287_ clknet_leaf_70_i_clk _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold771 net5541 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 net3799 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net6802 net6383 _04392_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__mux2_1
X_20764__192 clknet_1_1__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__inv_2
X_20238_ net3342 _03744_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__or2_1
Xhold793 _01093_ vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ net5591 _03705_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__or2_1
Xhold2150 net7226 vssd1 vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 rbzero.tex_r1\[63\] vssd1 vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2172 net7236 vssd1 vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2183 rbzero.tex_g1\[45\] vssd1 vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _06109_ _06110_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__nand2_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _04436_ vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1460 _01393_ vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1471 net6877 vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
X_11942_ _05108_ _05109_ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__o21ba_1
X_14730_ _07877_ _07880_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__nand2_1
Xhold1482 _01408_ vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1493 net6751 vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _07766_ _07784_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__xnor2_2
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11873_ _04983_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__or2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _09466_ _09471_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__or2_1
X_13612_ _06743_ _06758_ _06761_ _06762_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__o31a_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ net6606 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__clkbuf_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _10380_ sky130_fd_sc_hd__nand2_2
X_14592_ _07714_ _07737_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__xnor2_4
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16331_ _09403_ net7381 vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13543_ _06681_ _06683_ _06624_ _06685_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__and4b_2
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ net1954 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16262_ _09334_ _09335_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__nand2_1
X_19050_ net3096 _02988_ _03007_ _02993_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13474_ net3538 net3237 vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__and2_2
X_10686_ net5916 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18001_ _02033_ _02034_ _02048_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _08289_ net1008 _06258_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__mux2_1
X_12425_ _05177_ _05589_ _05591_ _05461_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16193_ _08802_ _09267_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15144_ net4566 _08025_ _08249_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12356_ _04975_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__nand2_1
X_20847__267 clknet_1_1__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__inv_2
XFILLER_0_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ net6846 net6614 _04529_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19952_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__inv_2
X_15075_ _08200_ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__buf_2
XFILLER_0_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12287_ _05069_ _05452_ _05454_ _05034_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__o211a_1
X_14026_ _07133_ _07166_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__a21oi_1
X_18903_ _02887_ _02888_ rbzero.wall_tracer.rayAddendY\[5\] _09932_ vssd1 vssd1 vccd1
+ vccd1 _02889_ sky130_fd_sc_hd__a2bb2o_1
X_11238_ net6539 net2412 _04492_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__mux2_1
X_19883_ net3995 _03503_ net4090 vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o21ai_1
X_18834_ net4459 net4640 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__nor2_1
X_11169_ net1485 net6441 _04459_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18765_ net4549 net1091 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__nor2_1
X_15977_ _09051_ _08755_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ _10130_ _09420_ _01766_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__or3_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14928_ _08075_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__clkbuf_1
X_18696_ _02579_ net4812 _02692_ net3044 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__a31o_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04004_ clknet_0__04004_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04004_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17647_ _10533_ _10535_ _10532_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14859_ net7908 _08009_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17578_ net7374 _10575_ vssd1 vssd1 vccd1 vccd1 _10576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_212_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19317_ net4214 _03160_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16529_ net3143 _08628_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19248_ net5172 _03119_ _03126_ _03115_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__o211a_1
Xhold7117 rbzero.traced_texa\[-1\] vssd1 vssd1 vccd1 vccd1 net7641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7128 rbzero.pov.ready_buffer\[13\] vssd1 vssd1 vccd1 vccd1 net7652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7139 rbzero.spi_registers.texadd2\[11\] vssd1 vssd1 vccd1 vccd1 net7663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6405 rbzero.tex_g1\[43\] vssd1 vssd1 vccd1 vccd1 net6929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6416 net2218 vssd1 vssd1 vccd1 vccd1 net6940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6427 rbzero.tex_b0\[17\] vssd1 vssd1 vccd1 vccd1 net6951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19179_ _03083_ net3145 vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__or2_1
Xhold6438 net1812 vssd1 vssd1 vccd1 vccd1 net6962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6449 _04474_ vssd1 vssd1 vccd1 vccd1 net6973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5704 rbzero.spi_registers.buf_sky\[3\] vssd1 vssd1 vccd1 vccd1 net6228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5715 _02552_ vssd1 vssd1 vccd1 vccd1 net6239 sky130_fd_sc_hd__dlygate4sd3_1
X_21210_ net4965 net6357 vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22190_ net322 net2050 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5726 _02950_ vssd1 vssd1 vccd1 vccd1 net6250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5737 _00424_ vssd1 vssd1 vccd1 vccd1 net6261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5748 _00814_ vssd1 vssd1 vccd1 vccd1 net6272 sky130_fd_sc_hd__dlygate4sd3_1
X_20906__320 clknet_1_0__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__inv_2
Xhold5759 _00423_ vssd1 vssd1 vccd1 vccd1 net6283 sky130_fd_sc_hd__dlygate4sd3_1
X_21141_ _04124_ _04125_ net4705 net65 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_111_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21072_ _04063_ _04064_ _04065_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20023_ _03581_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21974_ net199 net2333 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer30 net553 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer41 _06942_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer52 _06901_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer63 net586 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952__362 clknet_1_1__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__inv_2
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22457_ clknet_leaf_38_i_clk _01626_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ _05346_ _05376_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nor2_2
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21408_ clknet_leaf_79_i_clk net4481 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13190_ net2677 _06219_ _06216_ _04860_ _06345_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__a221o_1
X_22388_ net520 net1893 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
Xhold6983 net4203 vssd1 vssd1 vccd1 vccd1 net7507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ net4059 _04776_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__xnor2_1
X_21339_ clknet_leaf_42_i_clk net4132 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ rbzero.tex_r1\[39\] rbzero.tex_r1\[38\] _05071_ vssd1 vssd1 vccd1 vccd1 _05241_
+ sky130_fd_sc_hd__mux2_1
Xhold590 net5514 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net7260 net7012 _04310_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
X_15900_ _08952_ _08954_ _08953_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16880_ net4317 _09934_ _09936_ _08086_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
X_15831_ _08860_ _08897_ _08896_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__a21o_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _02561_ _02564_ _08246_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a21oi_1
X_15762_ _08827_ _08828_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__xnor2_2
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _06125_ _06127_ _06128_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__o211ai_4
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _10498_ _10499_ vssd1 vssd1 vccd1 vccd1 _10500_ sky130_fd_sc_hd__nor2_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 _01369_ vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _07862_ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__xnor2_1
X_11925_ net3218 vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__inv_2
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ net7360 rbzero.spi_registers.spi_cmd\[2\] _02501_ vssd1 vssd1 vccd1 vccd1
+ _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15693_ _08751_ _08767_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__xor2_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _10430_ _10431_ vssd1 vssd1 vccd1 vccd1 _10432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11856_ _04960_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__xnor2_1
X_14644_ _07743_ _07789_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__xor2_4
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10807_ net7165 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__clkbuf_1
X_17363_ _10258_ _10262_ _10362_ vssd1 vssd1 vccd1 vccd1 _10363_ sky130_fd_sc_hd__a21oi_1
X_14575_ _07697_ _07698_ _07699_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__a21o_1
X_11787_ _04944_ _04953_ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19102_ net5908 _03037_ _03041_ _03022_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__o211a_1
X_16314_ _09386_ _09387_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__and2b_1
Xclkbuf_0__05840_ _05840_ vssd1 vssd1 vccd1 vccd1 clknet_0__05840_ sky130_fd_sc_hd__clkbuf_16
X_10738_ net7249 net5886 _04236_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__mux2_1
X_13526_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17294_ _10172_ _10173_ _08584_ vssd1 vssd1 vccd1 vccd1 _10295_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19033_ net3958 _02988_ _02997_ _02993_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__o211a_1
X_16245_ _09317_ _09318_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__xnor2_1
X_13457_ _06503_ _06607_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__xor2_2
X_10669_ net2519 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ _04984_ _05574_ _05000_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16176_ _09250_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13388_ _06517_ _06528_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12339_ _05499_ _05506_ _05022_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15127_ net4599 net4513 _08219_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__mux2_1
Xhold3609 net7573 vssd1 vssd1 vccd1 vccd1 net4133 sky130_fd_sc_hd__dlygate4sd3_1
X_19935_ net1018 _03470_ _03480_ _03551_ _03529_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__o221a_1
X_15058_ _06625_ _08150_ _08154_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2908 net4500 vssd1 vssd1 vccd1 vccd1 net3432 sky130_fd_sc_hd__buf_1
X_14009_ _06970_ _07159_ _06869_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__mux2_1
Xhold2919 _01218_ vssd1 vssd1 vccd1 vccd1 net3443 sky130_fd_sc_hd__dlygate4sd3_1
X_19866_ net2999 _08467_ _03484_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18817_ _05396_ net4438 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__nand2_1
X_19797_ net6058 _03442_ net1567 _03441_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__o211a_1
X_18748_ net3281 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18679_ _02579_ net4697 net7572 net3689 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21690_ clknet_leaf_26_i_clk net5199 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20641_ net3930 _03972_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20572_ net2927 net3752 _03911_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22311_ net443 net2477 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6202 net1754 vssd1 vssd1 vccd1 vccd1 net6726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6213 _04483_ vssd1 vssd1 vccd1 vccd1 net6737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6224 net2074 vssd1 vssd1 vccd1 vccd1 net6748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6235 rbzero.tex_r1\[32\] vssd1 vssd1 vccd1 vccd1 net6759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22242_ net374 net1773 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold6246 net2048 vssd1 vssd1 vccd1 vccd1 net6770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5501 net3908 vssd1 vssd1 vccd1 vccd1 net6025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6257 rbzero.tex_r1\[44\] vssd1 vssd1 vccd1 vccd1 net6781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5512 rbzero.spi_registers.buf_texadd3\[21\] vssd1 vssd1 vccd1 vccd1 net6036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6268 net1794 vssd1 vssd1 vccd1 vccd1 net6792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5523 net2948 vssd1 vssd1 vccd1 vccd1 net6047 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5534 net1591 vssd1 vssd1 vccd1 vccd1 net6058 sky130_fd_sc_hd__clkbuf_2
Xhold6279 rbzero.tex_b0\[27\] vssd1 vssd1 vccd1 vccd1 net6803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4800 net905 vssd1 vssd1 vccd1 vccd1 net5324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5545 net3164 vssd1 vssd1 vccd1 vccd1 net6069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22173_ net305 net1075 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold4811 _01592_ vssd1 vssd1 vccd1 vccd1 net5335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5556 net3204 vssd1 vssd1 vccd1 vccd1 net6080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5567 _08204_ vssd1 vssd1 vccd1 vccd1 net6091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4822 net975 vssd1 vssd1 vccd1 vccd1 net5346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4833 _00693_ vssd1 vssd1 vccd1 vccd1 net5357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5578 net3409 vssd1 vssd1 vccd1 vccd1 net6102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5589 rbzero.spi_registers.buf_texadd3\[16\] vssd1 vssd1 vccd1 vccd1 net6113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4844 _00821_ vssd1 vssd1 vccd1 vccd1 net5368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21124_ _04108_ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__xnor2_1
Xhold4855 net945 vssd1 vssd1 vccd1 vccd1 net5379 sky130_fd_sc_hd__buf_1
Xhold4866 rbzero.spi_registers.buf_texadd0\[9\] vssd1 vssd1 vccd1 vccd1 net5390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4877 rbzero.spi_registers.buf_otherx\[4\] vssd1 vssd1 vccd1 vccd1 net5401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4888 rbzero.spi_registers.texadd3\[18\] vssd1 vssd1 vccd1 vccd1 net5412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4899 rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 net5423 sky130_fd_sc_hd__dlygate4sd3_1
X_21055_ _04048_ _04049_ _04050_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__o21a_1
X_20006_ rbzero.debug_overlay.facingY\[-7\] net3728 _03594_ vssd1 vssd1 vccd1 vccd1
+ _03603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21957_ net182 net2270 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
X_20876__293 clknet_1_0__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__inv_2
XFILLER_0_154_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _04862_ _04871_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__or3_1
XFILLER_0_178_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12690_ net15 _05850_ net11 net12 vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__and4b_1
X_21888_ clknet_leaf_97_i_clk net1273 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11641_ net3988 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__clkbuf_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14360_ _07473_ _07489_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__xnor2_1
X_11572_ _04714_ _04689_ _04741_ _04743_ _04160_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a311o_1
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__inv_2
Xinput19 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14291_ _07440_ _07441_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ _09086_ _08517_ _09085_ vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__or3_1
X_13242_ net2388 _06396_ _06202_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_165_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7492 _06158_ vssd1 vssd1 vccd1 vccd1 net8016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6780 net2861 vssd1 vssd1 vccd1 vccd1 net7304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ _06282_ _06284_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__04007_ clknet_0__04007_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04007_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6791 _02496_ vssd1 vssd1 vccd1 vccd1 net7315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _05028_ _05266_ _05274_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ _02027_ _02028_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19720_ net6172 _03393_ net2534 _03400_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__o211a_1
X_12055_ rbzero.tex_r1\[57\] rbzero.tex_r1\[56\] _05077_ vssd1 vssd1 vccd1 vccd1 _05224_
+ sky130_fd_sc_hd__mux2_1
X_16932_ _06221_ _08381_ vssd1 vssd1 vccd1 vccd1 _09950_ sky130_fd_sc_hd__xnor2_1
X_11006_ net7131 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__clkbuf_1
X_19651_ net6608 _03362_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__or2_1
X_16863_ _04165_ _04637_ _04603_ _04760_ vssd1 vssd1 vccd1 vccd1 _09924_ sky130_fd_sc_hd__and4_1
XFILLER_0_205_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20959__368 clknet_1_1__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__inv_2
X_18602_ _02611_ _02612_ _04624_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a21o_1
X_15814_ _08887_ _08888_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__nor2_1
X_19582_ _02501_ net797 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nor2_1
X_16794_ net3717 _09304_ vssd1 vssd1 vccd1 vccd1 _09864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18533_ net6237 net2919 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__nor2_1
X_15745_ _08819_ _08395_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _05077_ vssd1 vssd1 vccd1 vccd1 _05078_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _02487_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__clkbuf_1
X_15676_ _08750_ _08677_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__xor2_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _06045_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _09863_ _09864_ vssd1 vssd1 vccd1 vccd1 _10415_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _07772_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__xnor2_4
X_11839_ net80 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__buf_6
X_18395_ _02421_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _09538_ _09328_ _09447_ _09662_ vssd1 vssd1 vccd1 vccd1 _10346_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14558_ _07471_ _07524_ _07706_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03984_ clknet_0__03984_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03984_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _06659_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__clkbuf_2
X_17277_ _10276_ _10277_ vssd1 vssd1 vccd1 vccd1 _10278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14489_ _07562_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19016_ net3376 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
X_16228_ _09205_ _09185_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4107 _03583_ vssd1 vssd1 vccd1 vccd1 net4631 sky130_fd_sc_hd__dlygate4sd3_1
X_16159_ _09221_ _09233_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__xnor2_2
Xhold4118 _01020_ vssd1 vssd1 vccd1 vccd1 net4642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4129 net1504 vssd1 vssd1 vccd1 vccd1 net4653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3406 _05827_ vssd1 vssd1 vccd1 vccd1 net3930 sky130_fd_sc_hd__buf_4
Xhold3417 _03000_ vssd1 vssd1 vccd1 vccd1 net3941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_107_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3428 rbzero.debug_overlay.playerY\[5\] vssd1 vssd1 vccd1 vccd1 net3952 sky130_fd_sc_hd__buf_2
Xhold3439 _00951_ vssd1 vssd1 vccd1 vccd1 net3963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2705 rbzero.pov.ready_buffer\[18\] vssd1 vssd1 vccd1 vccd1 net3229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2716 net4466 vssd1 vssd1 vccd1 vccd1 net3240 sky130_fd_sc_hd__buf_1
X_19918_ _08377_ _03480_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_1
Xhold2727 _03943_ vssd1 vssd1 vccd1 vccd1 net3251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 rbzero.wall_tracer.visualWallDist\[-5\] vssd1 vssd1 vccd1 vccd1 net3262
+ sky130_fd_sc_hd__buf_2
Xhold2749 _08266_ vssd1 vssd1 vccd1 vccd1 net3273 sky130_fd_sc_hd__buf_1
XFILLER_0_177_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19849_ net4306 _03475_ net1157 _03454_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__o211a_1
X_21811_ clknet_leaf_10_i_clk net4677 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21742_ clknet_leaf_21_i_clk net4260 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21673_ clknet_leaf_14_i_clk net818 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdx\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20624_ _05825_ net3965 net4021 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20555_ net3490 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
Xhold6010 rbzero.tex_b0\[35\] vssd1 vssd1 vccd1 vccd1 net6534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6021 net1527 vssd1 vssd1 vccd1 vccd1 net6545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6032 rbzero.spi_registers.sclk_buffer\[1\] vssd1 vssd1 vccd1 vccd1 net6556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6043 rbzero.spi_registers.buf_texadd2\[1\] vssd1 vssd1 vccd1 vccd1 net6567 sky130_fd_sc_hd__dlygate4sd3_1
X_20486_ net3775 net1475 _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__mux2_1
Xhold6054 net1551 vssd1 vssd1 vccd1 vccd1 net6578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5320 rbzero.tex_g1\[46\] vssd1 vssd1 vccd1 vccd1 net5844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6065 rbzero.spi_registers.buf_texadd3\[3\] vssd1 vssd1 vccd1 vccd1 net6589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5331 _04351_ vssd1 vssd1 vccd1 vccd1 net5855 sky130_fd_sc_hd__dlygate4sd3_1
X_22225_ net357 net2773 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
Xhold6076 net1621 vssd1 vssd1 vccd1 vccd1 net6600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5342 _04497_ vssd1 vssd1 vccd1 vccd1 net5866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6087 _04417_ vssd1 vssd1 vccd1 vccd1 net6611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5353 _00663_ vssd1 vssd1 vccd1 vccd1 net5877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6098 net1729 vssd1 vssd1 vccd1 vccd1 net6622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5364 net2394 vssd1 vssd1 vccd1 vccd1 net5888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5375 net1781 vssd1 vssd1 vccd1 vccd1 net5899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4630 rbzero.spi_registers.buf_mapdx\[2\] vssd1 vssd1 vccd1 vccd1 net5154 sky130_fd_sc_hd__dlygate4sd3_1
X_22156_ net288 net2214 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
Xhold5386 rbzero.tex_r0\[2\] vssd1 vssd1 vccd1 vccd1 net5910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4641 net917 vssd1 vssd1 vccd1 vccd1 net5165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5397 _04455_ vssd1 vssd1 vccd1 vccd1 net5921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4652 _01066_ vssd1 vssd1 vccd1 vccd1 net5176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4663 _00847_ vssd1 vssd1 vccd1 vccd1 net5187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4674 _00859_ vssd1 vssd1 vccd1 vccd1 net5198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21107_ _04018_ _04096_ _04097_ _03083_ net4469 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a32o_1
Xhold3940 _03630_ vssd1 vssd1 vccd1 vccd1 net4464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4685 net1245 vssd1 vssd1 vccd1 vccd1 net5209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3951 net3327 vssd1 vssd1 vccd1 vccd1 net4475 sky130_fd_sc_hd__buf_1
Xhold4696 _01083_ vssd1 vssd1 vccd1 vccd1 net5220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22087_ clknet_leaf_74_i_clk net4024 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold3962 net7531 vssd1 vssd1 vccd1 vccd1 net4486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3973 net3381 vssd1 vssd1 vccd1 vccd1 net4497 sky130_fd_sc_hd__buf_1
Xhold3984 net7887 vssd1 vssd1 vccd1 vccd1 net4508 sky130_fd_sc_hd__dlygate4sd3_1
X_21038_ net985 net5424 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__nor2_1
Xhold3995 net1495 vssd1 vssd1 vccd1 vccd1 net4519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13860_ _06874_ _06878_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__or2b_1
XFILLER_0_57_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12811_ net4021 _05946_ _05956_ _05299_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13791_ _06939_ _06940_ _06941_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15530_ _08150_ _08104_ _08159_ _08047_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__a211oi_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ net21 _05901_ net17 net18 vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__and4b_1
XFILLER_0_85_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _05833_ _05834_ net7 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__mux2_1
X_15461_ _08534_ _08535_ _08295_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__a21o_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17200_ _09904_ _10201_ vssd1 vssd1 vccd1 vccd1 _10202_ sky130_fd_sc_hd__xnor2_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _07471_ _07509_ _07489_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__o21bai_2
X_11624_ _04727_ _04721_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__o21ai_1
X_18180_ _02225_ _02226_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__and2_1
X_20345__77 clknet_1_1__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
X_15392_ net3028 _08439_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17131_ _10131_ _10132_ vssd1 vssd1 vccd1 vccd1 _10133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14343_ _07492_ _07493_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__nand2_1
X_11555_ _04726_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17062_ _10066_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__clkbuf_1
X_14274_ _07416_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ rbzero.texu_hot\[1\] _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16013_ _09085_ _09087_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ _06185_ _06368_ _06380_ _06263_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ net3184 vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__inv_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ rbzero.tex_r1\[17\] rbzero.tex_r1\[16\] _05071_ vssd1 vssd1 vccd1 vccd1 _05276_
+ sky130_fd_sc_hd__mux2_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _02010_ _02011_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__and2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _06239_ _06240_ _06241_ _06242_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19703_ net1572 _03393_ net5729 _03384_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__o211a_1
X_12038_ net42 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__buf_6
X_16915_ net1144 _09941_ _09942_ net6123 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a22o_1
X_17895_ _01833_ _01837_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19634_ net5034 net798 _03353_ _03354_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__o211a_1
X_16846_ _04165_ net3976 vssd1 vssd1 vccd1 vccd1 _09915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19565_ net3112 _03305_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__or2_1
X_16777_ _09831_ _09832_ _09846_ vssd1 vssd1 vccd1 vccd1 _09847_ sky130_fd_sc_hd__a21o_1
X_13989_ _07099_ _07100_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ net4656 net715 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__or2_1
X_15728_ _08791_ _08792_ _08801_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19496_ net5783 _03266_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18447_ _09987_ _02472_ _02171_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a21o_1
X_15659_ _08433_ _08497_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18378_ _02412_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17329_ _06204_ _10329_ vssd1 vssd1 vccd1 vccd1 _10330_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03998_ _03998_ vssd1 vssd1 vccd1 vccd1 clknet_0__03998_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20271_ net3752 _03756_ net4840 _03761_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22010_ clknet_leaf_100_i_clk net3740 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3203 _00604_ vssd1 vssd1 vccd1 vccd1 net3727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3214 _03792_ vssd1 vssd1 vccd1 vccd1 net3738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3225 _02969_ vssd1 vssd1 vccd1 vccd1 net3749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3236 net7352 vssd1 vssd1 vccd1 vccd1 net3760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3247 _01003_ vssd1 vssd1 vccd1 vccd1 net3771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2502 net4682 vssd1 vssd1 vccd1 vccd1 net3026 sky130_fd_sc_hd__clkbuf_4
Xhold3258 net1381 vssd1 vssd1 vccd1 vccd1 net3782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2513 rbzero.spi_registers.spi_buffer\[12\] vssd1 vssd1 vccd1 vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 _08220_ vssd1 vssd1 vccd1 vccd1 net3048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3269 net4638 vssd1 vssd1 vccd1 vccd1 net3793 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2535 _02475_ vssd1 vssd1 vccd1 vccd1 net3059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1801 net7144 vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2546 net910 vssd1 vssd1 vccd1 vccd1 net3070 sky130_fd_sc_hd__buf_2
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1812 _01448_ vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2557 rbzero.pov.ready_buffer\[57\] vssd1 vssd1 vccd1 vccd1 net3081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _04544_ vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 net4819 vssd1 vssd1 vccd1 vccd1 net3092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _04365_ vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2579 net7916 vssd1 vssd1 vccd1 vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1845 _01522_ vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1856 _04190_ vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 _04552_ vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 net6913 vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1889 _04502_ vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_190_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21725_ clknet_leaf_2_i_clk net6031 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21656_ clknet_leaf_15_i_clk net5461 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_othery\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20607_ net4014 _05825_ net3965 net4021 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or4b_1
X_21587_ clknet_leaf_22_i_clk net5644 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ net2400 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_97 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_97/HI o_rgb[9] sky130_fd_sc_hd__conb_1
X_20538_ _03902_ net3287 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ net6812 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20469_ net3695 net1433 _03845_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13010_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xor2_1
Xhold5150 net1404 vssd1 vssd1 vccd1 vccd1 net5674 sky130_fd_sc_hd__dlygate4sd3_1
X_22208_ net340 net1643 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
Xhold5161 _08162_ vssd1 vssd1 vccd1 vccd1 net5685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5172 net1440 vssd1 vssd1 vccd1 vccd1 net5696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5183 _00387_ vssd1 vssd1 vccd1 vccd1 net5707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5194 net1214 vssd1 vssd1 vccd1 vccd1 net5718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4460 _00739_ vssd1 vssd1 vccd1 vccd1 net4984 sky130_fd_sc_hd__dlygate4sd3_1
X_22139_ net271 net1858 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
Xhold4471 net753 vssd1 vssd1 vccd1 vccd1 net4995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4482 rbzero.spi_registers.texadd1\[18\] vssd1 vssd1 vccd1 vccd1 net5006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4493 rbzero.spi_registers.texadd3\[16\] vssd1 vssd1 vccd1 vccd1 net5017 sky130_fd_sc_hd__dlygate4sd3_1
X_20653__92 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__inv_2
X_21003__5 clknet_1_0__leaf__03773_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
Xhold3770 net7379 vssd1 vssd1 vccd1 vccd1 net4294 sky130_fd_sc_hd__clkbuf_2
Xhold3781 net1305 vssd1 vssd1 vccd1 vccd1 net4305 sky130_fd_sc_hd__dlygate4sd3_1
X_14961_ _08100_ _08105_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__nand2_2
Xhold3792 rbzero.row_render.size\[1\] vssd1 vssd1 vccd1 vccd1 net4316 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03987_ clknet_0__03987_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03987_
+ sky130_fd_sc_hd__clkbuf_16
X_16700_ _09769_ net3029 vssd1 vssd1 vccd1 vccd1 _09771_ sky130_fd_sc_hd__nor2_1
X_13912_ _07031_ _07039_ _07040_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__or3_1
X_17680_ _10583_ _01731_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__xnor2_1
X_14892_ net7908 _08019_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16631_ _08471_ _08574_ _08588_ _08516_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__o22ai_2
X_13843_ _06922_ _06993_ _06921_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19350_ net4211 _03172_ net1218 _03181_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__o211a_1
X_16562_ _09631_ _09633_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__nor2_1
X_10986_ net2004 net6636 _04366_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__mux2_1
X_13774_ _06921_ _06924_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__nand2_1
X_18301_ _02344_ net4467 _02338_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15513_ _08550_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ net6555 _05843_ _05883_ net56 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_1
X_19281_ net5298 _03132_ _03145_ _03142_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__o211a_1
X_16493_ _09562_ _08962_ _08698_ _08701_ vssd1 vssd1 vccd1 vccd1 _09565_ sky130_fd_sc_hd__and4b_1
XFILLER_0_73_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18232_ _02204_ _02233_ _02234_ _02202_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__o31a_1
X_15444_ _08516_ _08517_ _08518_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ net4021 _05786_ _05796_ _05299_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18163_ _02208_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ rbzero.texu_hot\[0\] _04659_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__or2_1
X_12587_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _05541_ vssd1 vssd1 vccd1 vccd1 _05752_
+ sky130_fd_sc_hd__mux2_1
X_15375_ _08449_ _08411_ _08424_ _08433_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_136_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17114_ _10107_ _10115_ vssd1 vssd1 vccd1 vccd1 _10116_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14326_ _07465_ _07469_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18094_ _02140_ _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__nor2_1
X_11538_ rbzero.spi_registers.texadd0\[23\] _04709_ _04159_ vssd1 vssd1 vccd1 vccd1
+ _04710_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold408 net2252 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17045_ net3462 net4716 vssd1 vssd1 vccd1 vccd1 _10051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold419 net5274 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ _07388_ _07389_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__or2_1
X_11469_ _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _06217_ net3984 _06185_ net3804 vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__or4_1
X_14188_ _07337_ _07338_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__nand2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _06282_ _06284_ _06291_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18996_ net3749 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20900__315 clknet_1_1__leaf__04003_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__inv_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _01993_ _01994_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__nand2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _03453_ vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 _01377_ vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17878_ _01925_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ _09691_ _09761_ _09759_ vssd1 vssd1 vccd1 vccd1 _09899_ sky130_fd_sc_hd__a21oi_1
X_19617_ net4115 net799 net698 _03343_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19548_ net614 _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _04597_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21510_ clknet_leaf_44_i_clk net1009 vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21441_ clknet_leaf_88_i_clk net4665 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_20324__58 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21372_ clknet_leaf_59_i_clk _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold920 _01135_ vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold931 _01523_ vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold942 _01582_ vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold953 net6499 vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
X_20254_ net5588 _03743_ _03754_ _03748_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__o211a_1
Xhold964 rbzero.tex_r0\[0\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 _01144_ vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3000 net725 vssd1 vssd1 vccd1 vccd1 net3524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 net5532 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3011 _04819_ vssd1 vssd1 vccd1 vccd1 net3535 sky130_fd_sc_hd__buf_2
Xhold3022 _01007_ vssd1 vssd1 vccd1 vccd1 net3546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 rbzero.tex_b0\[0\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3033 net1409 vssd1 vssd1 vccd1 vccd1 net3557 sky130_fd_sc_hd__dlygate4sd3_1
X_20185_ net3651 _03704_ _03715_ _03709_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__o211a_1
Xhold3044 net1316 vssd1 vssd1 vccd1 vccd1 net3568 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_90_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold2310 net4777 vssd1 vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3055 rbzero.pov.ready_buffer\[49\] vssd1 vssd1 vccd1 vccd1 net3579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2321 net7289 vssd1 vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3066 net1170 vssd1 vssd1 vccd1 vccd1 net3590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2332 _04212_ vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3077 _01230_ vssd1 vssd1 vccd1 vccd1 net3601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2343 _04511_ vssd1 vssd1 vccd1 vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3088 _03887_ vssd1 vssd1 vccd1 vccd1 net3612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2354 _01405_ vssd1 vssd1 vccd1 vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3099 _08285_ vssd1 vssd1 vccd1 vccd1 net3623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 _04303_ vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2365 net3579 vssd1 vssd1 vccd1 vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2376 net6019 vssd1 vssd1 vccd1 vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1631 net5860 vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1642 net6925 vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2387 net3364 vssd1 vssd1 vccd1 vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1653 net5905 vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2398 net3610 vssd1 vssd1 vccd1 vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1664 net6749 vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1675 _01293_ vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1686 _04339_ vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1697 net7072 vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ net6866 net6500 _04288_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10771_ net6652 net1976 _04255_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _05230_ vssd1 vssd1 vccd1 vccd1 _05676_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13490_ _06612_ _06552_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__or2_1
X_21708_ clknet_leaf_19_i_clk net1705 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12441_ _05207_ _05603_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21639_ clknet_leaf_34_i_clk net1536 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12372_ _05248_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15160_ net3419 _08125_ _08249_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11323_ net1962 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
X_14111_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15091_ net645 _08201_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11254_ net6377 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ _06819_ _06869_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18850_ _02837_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11185_ net6974 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17801_ _01849_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__xnor2_1
Xhold4290 net3045 vssd1 vssd1 vccd1 vccd1 net4814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18781_ net6222 _02775_ _02714_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
X_15993_ _09063_ _09066_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17732_ _01781_ _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__nand2_1
X_14944_ net7433 net7457 vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_203_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17663_ _10301_ _01710_ _01714_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a21oi_1
X_14875_ net4931 net4027 _04622_ _06207_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__and4b_2
X_19402_ net5338 _03211_ _03214_ _03207_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__o211a_1
X_16614_ _09543_ _09552_ _09684_ vssd1 vssd1 vccd1 vccd1 _09685_ sky130_fd_sc_hd__a21oi_1
X_13826_ _06971_ _06976_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__xnor2_2
X_17594_ _10590_ _10591_ vssd1 vssd1 vccd1 vccd1 _10592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19333_ net5714 _03172_ _03175_ _03168_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ _09600_ _09616_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13757_ _06903_ _06904_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__a21o_1
X_10969_ net6894 net7133 _04355_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19264_ net4991 _03133_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or2_1
X_12708_ net12 _05848_ _05868_ net14 vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a22o_1
X_16476_ _09425_ _09547_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13688_ _06808_ _06814_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18215_ _02254_ _02255_ _02260_ _02261_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a22o_1
X_15427_ _08497_ _08501_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12639_ net56 _05790_ net6 _05799_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a41o_2
X_19195_ _02992_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6609 net2765 vssd1 vssd1 vccd1 vccd1 net7133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _01812_ _10539_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _08432_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5908 rbzero.tex_g1\[28\] vssd1 vssd1 vccd1 vccd1 net6432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5919 net1268 vssd1 vssd1 vccd1 vccd1 net6443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 net6334 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ _07407_ _07395_ _07435_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18077_ _02122_ _02124_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__xor2_1
Xhold216 net3427 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ _08362_ _08363_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold227 net5921 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _01272_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 net7676 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _10032_ _10035_ vssd1 vssd1 vccd1 vccd1 _10036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _09955_ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__xnor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21990_ net215 net1104 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20718__151 clknet_1_1__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__inv_2
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22473_ clknet_leaf_80_i_clk net4907 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21424_ clknet_leaf_45_i_clk net3920 vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21355_ clknet_leaf_42_i_clk net5971 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold750 net5048 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
X_21286_ clknet_leaf_65_i_clk _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold761 net5384 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 net5618 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 net5637 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
X_20237_ net3342 _03743_ _03745_ _03735_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold794 net5386 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20168_ net5591 _03704_ _03706_ _03696_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__o211a_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 _01378_ vssd1 vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2151 _04343_ vssd1 vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2162 net2647 vssd1 vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2173 _01465_ vssd1 vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20099_ net4865 net4797 net3562 vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__a21boi_1
X_12990_ _06139_ _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nor2_1
Xhold2184 net2396 vssd1 vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1450 _04298_ vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2195 _01349_ vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1461 net6891 vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1472 _04401_ vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ _05008_ _04992_ _04977_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a31o_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1483 net6851 vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1494 net6753 vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14660_ _07809_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__nor2b_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _05014_ vssd1 vssd1 vccd1 vccd1 _05042_
+ sky130_fd_sc_hd__mux2_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _06657_ _06658_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ net6604 net2902 _04277_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
X_14591_ _07690_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__and2b_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ net7380 net2935 _08293_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _06665_ _06619_ _06666_ _06628_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a31oi_4
X_10754_ net7018 net7004 _04244_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ _08564_ _08471_ _08516_ _08529_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ net2556 net5914 _04203_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13473_ _06613_ _06596_ _06609_ _06623_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__or4_4
X_18000_ _02033_ _02034_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15212_ _06367_ _08283_ _06267_ net1312 vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__a2bb2o_1
X_12424_ _05019_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__or2_1
X_16192_ _09265_ _09266_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__xor2_2
XFILLER_0_164_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20303__39 clknet_1_1__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_0_152_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15143_ net4933 vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__buf_4
X_12355_ _05507_ _05522_ _05027_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11306_ net2614 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
X_12286_ _05248_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__or2_1
X_19951_ net3893 _03560_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__or2_1
X_15074_ _06203_ _06384_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ net5902 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
X_14025_ _07168_ _07172_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__a21o_1
X_18902_ _02871_ _02886_ _02884_ _04623_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a31o_1
X_19882_ net4090 net3995 _03503_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__or3_1
XFILLER_0_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11168_ net2579 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
X_18833_ net7612 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18764_ _02750_ _02758_ net4800 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__o21a_1
X_15976_ _08430_ _08431_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__nand2_4
X_11099_ net6668 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
X_17715_ _10257_ _09538_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ net4435 _08074_ _08027_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__mux2_1
X_18695_ _04633_ _02699_ _02700_ _09933_ net3043 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a32o_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__04003_ clknet_0__04003_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04003_
+ sky130_fd_sc_hd__clkbuf_16
X_17646_ _01672_ _01697_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _07968_ _07970_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__xnor2_1
X_13809_ _06954_ _06959_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17577_ net4403 net7373 vssd1 vssd1 vccd1 vccd1 _10575_ sky130_fd_sc_hd__or2_1
X_14789_ _07937_ _07939_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19316_ net5053 _03159_ _03165_ _03155_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__o211a_1
X_16528_ _09594_ _09599_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7107 _02626_ vssd1 vssd1 vccd1 vccd1 net7631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19247_ net5030 _03120_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__or2_1
X_16459_ _09439_ _09441_ _09438_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__a21o_2
XFILLER_0_147_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7118 rbzero.traced_texa\[7\] vssd1 vssd1 vccd1 vccd1 net7642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7129 rbzero.wall_tracer.mapX\[6\] vssd1 vssd1 vccd1 vccd1 net7653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6406 net2209 vssd1 vssd1 vccd1 vccd1 net6930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6417 rbzero.tex_r1\[24\] vssd1 vssd1 vccd1 vccd1 net6941 sky130_fd_sc_hd__dlygate4sd3_1
X_19178_ net3254 net3144 _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6428 net2268 vssd1 vssd1 vccd1 vccd1 net6952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6439 _04414_ vssd1 vssd1 vccd1 vccd1 net6963 sky130_fd_sc_hd__dlygate4sd3_1
X_18129_ _01834_ _02084_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nor2_1
Xhold5705 net1531 vssd1 vssd1 vccd1 vccd1 net6229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5716 _02553_ vssd1 vssd1 vccd1 vccd1 net6240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5727 net6268 vssd1 vssd1 vccd1 vccd1 net6251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5738 rbzero.spi_registers.buf_texadd3\[9\] vssd1 vssd1 vccd1 vccd1 net6262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21140_ _04119_ _04121_ _04123_ _09919_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a31o_1
Xhold5749 net2543 vssd1 vssd1 vccd1 vccd1 net6273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21071_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20022_ _03577_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21973_ net198 net2029 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer20 net543 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer31 _07104_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer42 _07062_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ clknet_1_1__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__buf_1
Xrebuffer53 _06900_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer64 _06827_ vssd1 vssd1 vccd1 vccd1 net3132 sky130_fd_sc_hd__clkbuf_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22456_ clknet_leaf_40_i_clk _01625_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6940 net7923 vssd1 vssd1 vccd1 vccd1 net7464 sky130_fd_sc_hd__dlygate4sd3_1
X_21407_ clknet_leaf_24_i_clk net629 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi
+ sky130_fd_sc_hd__dfxtp_1
X_22387_ net519 net2570 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
Xhold6951 rbzero.wall_tracer.stepDistX\[-3\] vssd1 vssd1 vccd1 vccd1 net7475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6962 rbzero.traced_texVinit\[2\] vssd1 vssd1 vccd1 vccd1 net7486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6973 rbzero.traced_texVinit\[3\] vssd1 vssd1 vccd1 vccd1 net7497 sky130_fd_sc_hd__dlygate4sd3_1
X_12140_ _05298_ _05303_ _05308_ _04853_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or4b_2
X_21338_ clknet_leaf_46_i_clk net4148 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6995 _00501_ vssd1 vssd1 vccd1 vccd1 net7519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ rbzero.tex_r1\[37\] rbzero.tex_r1\[36\] _05072_ vssd1 vssd1 vccd1 vccd1 _05240_
+ sky130_fd_sc_hd__mux2_1
X_21269_ clknet_leaf_50_i_clk _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold580 _01159_ vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold591 net5761 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net6487 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15830_ _08900_ _08901_ _08904_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__a21bo_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _08528_ _08835_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__xnor2_4
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ net3857 net3135 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__or2_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _10496_ _10497_ vssd1 vssd1 vccd1 vccd1 _10499_ sky130_fd_sc_hd__and2_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1280 net6799 vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 net6741 vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _06918_ _07354_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__nor2_1
X_11924_ _05028_ _05063_ _05076_ _05093_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a31o_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ net3074 net3150 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15692_ _08760_ _08765_ _08766_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__a21oi_2
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17431_ _10428_ _10429_ vssd1 vssd1 vccd1 vccd1 _10431_ sky130_fd_sc_hd__and2_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14643_ _07742_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__xnor2_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _04961_ _04926_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__and2b_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ net7163 net2845 _04266_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
X_17362_ _10360_ _10361_ vssd1 vssd1 vccd1 vccd1 _10362_ sky130_fd_sc_hd__xnor2_1
X_14574_ _07723_ _07724_ _07675_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__o21ai_4
X_11786_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19101_ net5255 _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__or2_1
X_16313_ _09383_ _09385_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13525_ _06667_ _06675_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__nor2_4
X_10737_ net5888 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__clkbuf_1
X_17293_ _09863_ _09864_ _09086_ vssd1 vssd1 vccd1 vccd1 _10294_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19032_ net1608 _02990_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__or2_1
X_16244_ _09253_ _09256_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13456_ _06540_ net82 _06515_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__o21ai_4
X_10668_ net6626 net2518 _04192_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12407_ rbzero.tex_g1\[11\] rbzero.tex_g1\[10\] _05541_ vssd1 vssd1 vccd1 vccd1 _05574_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _08312_ _09249_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__or2_2
X_13387_ _06433_ _06535_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o21a_1
X_10599_ net4050 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ _08218_ _08235_ net3719 _08215_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__o211a_1
X_12338_ _05502_ _05505_ net80 vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19934_ _08475_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__inv_2
X_15057_ _08187_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
X_12269_ net3921 _05351_ _05384_ net2935 _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2909 net4512 vssd1 vssd1 vccd1 vccd1 net3433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14008_ _06781_ _06876_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19865_ net6130 _03475_ net2929 _03496_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18816_ net3807 _05393_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19796_ net6114 _03443_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__or2_1
X_15959_ _09010_ _09011_ _09032_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__and3_1
X_18747_ net3280 net4821 _06394_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
X_20936__347 clknet_1_1__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__inv_2
XFILLER_0_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18678_ rbzero.wall_tracer.rayAddendX\[6\] _09933_ _02684_ _04633_ vssd1 vssd1 vccd1
+ vccd1 _02685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17629_ _01678_ _01679_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20640_ net4002 _03970_ _03973_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20571_ net3814 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22310_ net442 net1843 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold6203 rbzero.tex_b0\[42\] vssd1 vssd1 vccd1 vccd1 net6727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6214 net1924 vssd1 vssd1 vccd1 vccd1 net6738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6225 rbzero.tex_b1\[44\] vssd1 vssd1 vccd1 vccd1 net6749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22241_ net373 net2136 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold6236 net1774 vssd1 vssd1 vccd1 vccd1 net6760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5502 _01253_ vssd1 vssd1 vccd1 vccd1 net6026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6247 rbzero.tex_r0\[43\] vssd1 vssd1 vccd1 vccd1 net6771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6258 net2224 vssd1 vssd1 vccd1 vccd1 net6782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5513 net2230 vssd1 vssd1 vccd1 vccd1 net6037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6269 _04450_ vssd1 vssd1 vccd1 vccd1 net6793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5524 gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 net6048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5535 rbzero.spi_registers.buf_texadd3\[17\] vssd1 vssd1 vccd1 vccd1 net6059 sky130_fd_sc_hd__dlygate4sd3_1
X_22172_ net304 net1752 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold4801 rbzero.color_floor\[2\] vssd1 vssd1 vccd1 vccd1 net5325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5546 rbzero.spi_registers.buf_texadd1\[22\] vssd1 vssd1 vccd1 vccd1 net6070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4812 net873 vssd1 vssd1 vccd1 vccd1 net5336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5557 rbzero.debug_overlay.playerY\[-8\] vssd1 vssd1 vccd1 vccd1 net6081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4823 _00783_ vssd1 vssd1 vccd1 vccd1 net5347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5568 net3334 vssd1 vssd1 vccd1 vccd1 net6092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21123_ _04109_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__and2b_1
Xhold4834 net948 vssd1 vssd1 vccd1 vccd1 net5358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5579 rbzero.spi_registers.spi_buffer\[19\] vssd1 vssd1 vccd1 vccd1 net6103 sky130_fd_sc_hd__dlygate4sd3_1
X_20681__117 clknet_1_0__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__inv_2
Xhold4845 net982 vssd1 vssd1 vccd1 vccd1 net5369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4856 _00503_ vssd1 vssd1 vccd1 vccd1 net5380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4867 net1045 vssd1 vssd1 vccd1 vccd1 net5391 sky130_fd_sc_hd__dlygate4sd3_1
X_20987__14 clknet_1_1__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_0_121_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4878 net1021 vssd1 vssd1 vccd1 vccd1 net5402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4889 net1029 vssd1 vssd1 vccd1 vccd1 net5413 sky130_fd_sc_hd__dlygate4sd3_1
X_21054_ net4763 _03519_ _04014_ _04052_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a22o_1
X_20005_ net3296 _03578_ net4515 _03602_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21956_ net181 net2818 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ clknet_leaf_97_i_clk net1281 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11640_ net3987 net2986 net3868 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11571_ _04648_ _04678_ _04682_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__o31a_1
XFILLER_0_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20769_ clknet_1_0__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__buf_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _06452_ _06460_ _06454_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ _07356_ _07400_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ _06179_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__clkbuf_4
X_22439_ clknet_leaf_39_i_clk net4742 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7493 net7440 vssd1 vssd1 vccd1 vccd1 net8017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6770 net2613 vssd1 vssd1 vccd1 vccd1 net7294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6781 _04323_ vssd1 vssd1 vccd1 vccd1 net7305 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__04006_ clknet_0__04006_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04006_
+ sky130_fd_sc_hd__clkbuf_16
X_13172_ _06280_ _06286_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6792 _00841_ vssd1 vssd1 vccd1 vccd1 net7316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12123_ _04978_ _05278_ _05283_ _05291_ _05050_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__o311a_1
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20293__30 clknet_1_1__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
X_17980_ _02027_ _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12054_ _05069_ _05220_ _05222_ _05034_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o211a_1
X_16931_ _06222_ _09294_ vssd1 vssd1 vccd1 vccd1 _09949_ sky130_fd_sc_hd__or2_1
X_11005_ net2325 net7129 _04377_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__mux2_1
X_16862_ net4075 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__clkbuf_1
X_19650_ _02996_ _03360_ net2077 _03354_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15813_ _08879_ _08882_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__and2b_1
X_18601_ _02611_ _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__nor2_1
X_19581_ net796 _02497_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nand2_1
X_16793_ _09740_ _09608_ _09304_ vssd1 vssd1 vccd1 vccd1 _09863_ sky130_fd_sc_hd__a21o_2
X_18532_ net4478 _02541_ _02542_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__o21a_1
X_15744_ _08396_ _08374_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__and2_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ _06109_ _06110_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__nand3_1
XFILLER_0_172_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ _04986_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__buf_4
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _02486_ net4342 net4920 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_4
X_15675_ _08678_ _08670_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__nand2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12887_ reg_gpout\[4\] clknet_1_1__leaf__06044_ net45 vssd1 vssd1 vccd1 vccd1 _06045_
+ sky130_fd_sc_hd__mux2_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _10403_ _10413_ vssd1 vssd1 vccd1 vccd1 _10414_ sky130_fd_sc_hd__xnor2_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14626_ _07773_ _07775_ _07776_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__a21bo_4
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _04957_ _04971_ _04997_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__nor3_2
X_18394_ net4487 net4423 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17345_ _09447_ _09662_ _10223_ vssd1 vssd1 vccd1 vccd1 _10345_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _07706_ _07707_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1__f__03983_ clknet_0__03983_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03983_
+ sky130_fd_sc_hd__clkbuf_16
X_11769_ _04934_ _04935_ net1583 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13508_ _06657_ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__nand2_2
X_17276_ _10255_ _10256_ _10275_ vssd1 vssd1 vccd1 vccd1 _10277_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _07520_ _07561_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19015_ _02982_ _02523_ net3375 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__and3b_1
X_16227_ _09268_ _09270_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__or2_4
X_13439_ _06540_ net82 _06516_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _09230_ _09232_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4108 _00985_ vssd1 vssd1 vccd1 vccd1 net4632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4119 net720 vssd1 vssd1 vccd1 vccd1 net4643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15109_ net3460 net3054 _08219_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3407 _01262_ vssd1 vssd1 vccd1 vccd1 net3931 sky130_fd_sc_hd__dlygate4sd3_1
X_16089_ _09149_ _09162_ _09163_ _09160_ _09161_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__o32a_1
Xhold3418 _03003_ vssd1 vssd1 vccd1 vccd1 net3942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3429 _03575_ vssd1 vssd1 vccd1 vccd1 net3953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2706 _03824_ vssd1 vssd1 vccd1 vccd1 net3230 sky130_fd_sc_hd__dlygate4sd3_1
X_19917_ net4893 _03530_ _03539_ _03496_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__o211a_1
Xhold2717 rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 net3241 sky130_fd_sc_hd__clkbuf_2
Xhold2728 _03944_ vssd1 vssd1 vccd1 vccd1 net3252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2739 net6125 vssd1 vssd1 vccd1 vccd1 net3263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19848_ net1156 _03477_ _03479_ _03486_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19779_ _08274_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__buf_4
X_21810_ clknet_leaf_10_i_clk net2894 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21741_ clknet_leaf_23_i_clk net1808 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire88 net3970 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_2
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21672_ clknet_leaf_13_i_clk net931 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20623_ net4021 _09929_ _03961_ net4018 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20554_ _03902_ net3489 vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__and2_1
Xhold6000 net1540 vssd1 vssd1 vccd1 vccd1 net6524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6011 net1497 vssd1 vssd1 vccd1 vccd1 net6535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6022 rbzero.tex_b1\[62\] vssd1 vssd1 vccd1 vccd1 net6546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ net3250 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__clkbuf_4
Xhold6033 net1577 vssd1 vssd1 vccd1 vccd1 net6557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6044 net1909 vssd1 vssd1 vccd1 vccd1 net6568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6055 _04272_ vssd1 vssd1 vccd1 vccd1 net6579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5310 rbzero.tex_g0\[34\] vssd1 vssd1 vccd1 vccd1 net5834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5321 _04336_ vssd1 vssd1 vccd1 vccd1 net5845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22224_ net356 net1984 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
Xhold6066 net1686 vssd1 vssd1 vccd1 vccd1 net6590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5332 net2002 vssd1 vssd1 vccd1 vccd1 net5856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6077 rbzero.spi_registers.buf_texadd1\[1\] vssd1 vssd1 vccd1 vccd1 net6601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5343 net2120 vssd1 vssd1 vccd1 vccd1 net5867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6088 net1878 vssd1 vssd1 vccd1 vccd1 net6612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5354 rbzero.tex_g1\[3\] vssd1 vssd1 vccd1 vccd1 net5878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6099 rbzero.spi_registers.buf_texadd3\[1\] vssd1 vssd1 vccd1 vccd1 net6623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5365 rbzero.tex_b1\[3\] vssd1 vssd1 vccd1 vccd1 net5889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4620 _00793_ vssd1 vssd1 vccd1 vccd1 net5144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5376 rbzero.tex_b1\[24\] vssd1 vssd1 vccd1 vccd1 net5900 sky130_fd_sc_hd__dlygate4sd3_1
X_22155_ net287 net2567 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold4631 net853 vssd1 vssd1 vccd1 vccd1 net5155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4642 _00723_ vssd1 vssd1 vccd1 vccd1 net5166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5387 net2562 vssd1 vssd1 vccd1 vccd1 net5911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5398 net751 vssd1 vssd1 vccd1 vccd1 net5922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4653 rbzero.spi_registers.buf_vshift\[3\] vssd1 vssd1 vccd1 vccd1 net5177 sky130_fd_sc_hd__dlygate4sd3_1
X_21106_ _04093_ _04094_ _04095_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4664 net883 vssd1 vssd1 vccd1 vccd1 net5188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3930 net7838 vssd1 vssd1 vccd1 vccd1 net4454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4675 net810 vssd1 vssd1 vccd1 vccd1 net5199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4686 _01045_ vssd1 vssd1 vccd1 vccd1 net5210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3941 _01013_ vssd1 vssd1 vccd1 vccd1 net4465 sky130_fd_sc_hd__dlygate4sd3_1
X_22086_ clknet_leaf_73_i_clk net3967 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3952 net4492 vssd1 vssd1 vccd1 vccd1 net4476 sky130_fd_sc_hd__buf_2
Xhold4697 rbzero.spi_registers.buf_texadd0\[8\] vssd1 vssd1 vccd1 vccd1 net5221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3963 net3314 vssd1 vssd1 vccd1 vccd1 net4487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3974 net7545 vssd1 vssd1 vccd1 vccd1 net4498 sky130_fd_sc_hd__dlygate4sd3_1
X_21037_ _04033_ _04034_ _04035_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o21a_1
Xhold3985 net2869 vssd1 vssd1 vccd1 vccd1 net4509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_156_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12810_ net26 _05965_ _05968_ net27 vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and4bb_1
X_13790_ _06736_ _06860_ net79 _06914_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__or4_4
XFILLER_0_9_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12741_ net20 _05898_ _05899_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ clknet_leaf_9_i_clk net4870 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _08130_ _08137_ _08144_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__or3_1
X_12672_ _04159_ _04718_ _04726_ _04777_ net4 net5 vssd1 vssd1 vccd1 vccd1 _05834_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14411_ _07520_ _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__nor2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11623_ _04714_ _04160_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__nand2_1
X_15391_ net695 _08465_ _08305_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17130_ _08317_ _08331_ _08548_ _08556_ vssd1 vssd1 vccd1 vccd1 _10132_ sky130_fd_sc_hd__or4_1
X_14342_ _07474_ _07471_ net558 vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__or3_4
XFILLER_0_53_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11554_ net6049 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17061_ _10065_ net3795 net4903 vssd1 vssd1 vccd1 vccd1 _10066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ _07417_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ rbzero.spi_registers.texadd3\[7\] rbzero.spi_registers.texadd1\[7\] rbzero.spi_registers.texadd0\[7\]
+ rbzero.spi_registers.texadd2\[7\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16012_ _09086_ _08517_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__nor2_1
Xhold7290 rbzero.wall_tracer.stepDistX\[7\] vssd1 vssd1 vccd1 vccd1 net7814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ _06217_ _06216_ _06369_ _06378_ _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__a311o_1
XFILLER_0_150_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__inv_2
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ rbzero.tex_r1\[19\] rbzero.tex_r1\[18\] _05219_ vssd1 vssd1 vccd1 vccd1 _05275_
+ sky130_fd_sc_hd__mux2_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _02010_ _02011_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__nor2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13086_ net2787 net1249 net977 net2768 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__or4_1
X_19702_ net5728 _03395_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__or2_1
X_12037_ net826 net7325 _05120_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__mux2_1
X_16914_ net1100 _09941_ _09942_ net7476 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17894_ _01836_ _01943_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19633_ _03294_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__clkbuf_4
X_16845_ _04164_ _04161_ net3975 vssd1 vssd1 vccd1 vccd1 _09914_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16776_ _09838_ _09845_ vssd1 vssd1 vccd1 vccd1 _09846_ sky130_fd_sc_hd__xnor2_1
X_19564_ net5371 _03303_ _03313_ _03314_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__o211a_1
X_13988_ _07135_ _07137_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_137_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15727_ _08791_ _08792_ _08801_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__a21oi_2
X_18515_ net4424 net701 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12939_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _03000_ _03265_ net2591 _03260_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__o211a_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15658_ _08731_ _08732_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18446_ _02470_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ _07753_ _07759_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__or2_1
X_18377_ _02410_ net4538 _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
X_15589_ _08663_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17328_ _10326_ _10328_ vssd1 vssd1 vccd1 vccd1 _10329_ sky130_fd_sc_hd__xor2_4
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20712__146 clknet_1_1__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__inv_2
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ _10259_ _08641_ _08754_ _08701_ vssd1 vssd1 vccd1 vccd1 _10260_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_0__03997_ _03997_ vssd1 vssd1 vccd1 vccd1 clknet_0__03997_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20270_ net3812 net4839 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3204 rbzero.pov.ready_buffer\[24\] vssd1 vssd1 vccd1 vccd1 net3728 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3215 _03793_ vssd1 vssd1 vccd1 vccd1 net3739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3226 _00621_ vssd1 vssd1 vccd1 vccd1 net3750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3237 _04813_ vssd1 vssd1 vccd1 vccd1 net3761 sky130_fd_sc_hd__buf_1
Xhold3248 net678 vssd1 vssd1 vccd1 vccd1 net3772 sky130_fd_sc_hd__clkbuf_2
Xhold2503 net4684 vssd1 vssd1 vccd1 vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3259 _03850_ vssd1 vssd1 vccd1 vccd1 net3783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 net616 vssd1 vssd1 vccd1 vccd1 net3038 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2525 net6283 vssd1 vssd1 vccd1 vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2536 _02482_ vssd1 vssd1 vccd1 vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1802 _04381_ vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2547 _00642_ vssd1 vssd1 vccd1 vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1813 net2366 vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 _03570_ vssd1 vssd1 vccd1 vccd1 net3082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1824 _01158_ vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2569 net6171 vssd1 vssd1 vccd1 vccd1 net3093 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1835 _01413_ vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1846 net6919 vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1857 _01568_ vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1868 _01151_ vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
X_20793__218 clknet_1_0__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__inv_2
Xhold1879 _04424_ vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ clknet_leaf_4_i_clk net4226 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21655_ clknet_leaf_15_i_clk net5404 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_otherx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20606_ _03947_ net4021 _05825_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21586_ clknet_leaf_22_i_clk net5596 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20687__123 clknet_1_1__leaf__03982_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__inv_2
Xtop_ew_algofoogle_98 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_98/HI o_rgb[10] sky130_fd_sc_hd__conb_1
X_20537_ net3286 net1400 _03889_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ net2653 net6810 _04514_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20468_ net3711 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5140 rbzero.pov.spi_buffer\[54\] vssd1 vssd1 vccd1 vccd1 net5664 sky130_fd_sc_hd__dlygate4sd3_1
X_22207_ net339 net2552 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
Xhold5151 _00759_ vssd1 vssd1 vccd1 vccd1 net5675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5162 _08169_ vssd1 vssd1 vccd1 vccd1 net5686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5173 _01017_ vssd1 vssd1 vccd1 vccd1 net5697 sky130_fd_sc_hd__dlygate4sd3_1
X_20399_ net3606 net1286 _03801_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__mux2_1
Xhold5184 net2769 vssd1 vssd1 vccd1 vccd1 net5708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4450 rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 net4974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5195 _03415_ vssd1 vssd1 vccd1 vccd1 net5719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4461 net780 vssd1 vssd1 vccd1 vccd1 net4985 sky130_fd_sc_hd__dlygate4sd3_1
X_22138_ net270 net1925 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4472 _00738_ vssd1 vssd1 vccd1 vccd1 net4996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4483 net763 vssd1 vssd1 vccd1 vccd1 net5007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4494 net855 vssd1 vssd1 vccd1 vccd1 net5018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3760 net1793 vssd1 vssd1 vccd1 vccd1 net4284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3771 _00974_ vssd1 vssd1 vccd1 vccd1 net4295 sky130_fd_sc_hd__dlygate4sd3_1
X_14960_ _08068_ _08104_ net6162 vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__a21oi_1
X_22069_ clknet_leaf_8_i_clk net3735 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3782 net7752 vssd1 vssd1 vccd1 vccd1 net4306 sky130_fd_sc_hd__clkbuf_2
Xhold3793 net3016 vssd1 vssd1 vccd1 vccd1 net4317 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03986_ clknet_0__03986_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03986_
+ sky130_fd_sc_hd__clkbuf_16
X_13911_ _07060_ _07061_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__xnor2_2
X_14891_ _07991_ _08017_ _08040_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16630_ _08470_ _08484_ _08574_ _08550_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__or4_1
X_13842_ _06960_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16561_ _09442_ _09508_ _09632_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__a21oi_1
X_13773_ _06736_ _06922_ _06923_ _06611_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10985_ net2135 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__clkbuf_1
X_15512_ _08387_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__clkbuf_4
X_18300_ _06206_ net7793 _10002_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__o21ai_1
X_12724_ net50 _05843_ _05852_ _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a31o_2
X_19280_ net1703 _03133_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__or2_1
X_16492_ _08701_ _08962_ _09563_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18231_ _02207_ _02231_ _02233_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a21oi_1
X_15443_ _08470_ _08492_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ net4020 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18162_ _08634_ _09538_ _02117_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ _04660_ _04662_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nand2_1
X_15374_ _08405_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__clkbuf_4
X_12586_ _05035_ _05746_ _05748_ _05750_ _04979_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17113_ _10108_ _10114_ vssd1 vssd1 vccd1 vccd1 _10115_ sky130_fd_sc_hd__xnor2_2
X_14325_ _07473_ _07475_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__xor2_1
X_18093_ _02001_ _02009_ _02007_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _04692_ _04693_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 _04334_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ _10041_ _10042_ _10043_ vssd1 vssd1 vccd1 vccd1 _10050_ sky130_fd_sc_hd__o21a_1
X_14256_ _07343_ _07393_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__nand2_2
X_11468_ _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__nor2_4
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ _06221_ net4897 _06244_ _06354_ _06362_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a221o_1
X_14187_ _07274_ _07309_ _07336_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__nand3_1
X_11399_ net2693 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ net3327 _06283_ _06292_ _06293_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a211o_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _02966_ _02967_ net3748 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__and3b_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17946_ _01993_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__or2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _04894_ _06216_ _06218_ _06220_ _06224_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o221a_1
Xhold1109 _00944_ vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
X_17877_ _01812_ _09484_ _01811_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__o31a_1
X_19616_ net3088 _03340_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or2_1
X_16828_ _09829_ _09897_ vssd1 vssd1 vccd1 vccd1 _09898_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19547_ net7312 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__buf_2
X_16759_ _09793_ _09828_ vssd1 vssd1 vccd1 vccd1 _09829_ sky130_fd_sc_hd__xnor2_1
X_19478_ _03000_ net3077 net1541 _03260_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309__45 clknet_1_0__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_0_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18429_ _02454_ _02455_ _01870_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21440_ clknet_leaf_87_i_clk net4761 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21371_ clknet_leaf_59_i_clk _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20322_ clknet_1_1__leaf__03773_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__buf_1
XFILLER_0_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold910 net5234 vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 net6484 vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 net4541 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20253_ net3568 _03744_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold943 net6306 vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 net6501 vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 net5776 vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3001 _03939_ vssd1 vssd1 vccd1 vccd1 net3525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 net7722 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__buf_1
Xhold987 net5534 vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3012 _01612_ vssd1 vssd1 vccd1 vccd1 net3536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 net5768 vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
X_20184_ net3557 _03705_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__or2_1
Xhold3023 rbzero.pov.ready_buffer\[26\] vssd1 vssd1 vccd1 vccd1 net3547 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3034 _03843_ vssd1 vssd1 vccd1 vccd1 net3558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3045 _03909_ vssd1 vssd1 vccd1 vccd1 net3569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2300 net5994 vssd1 vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3056 net2889 vssd1 vssd1 vccd1 vccd1 net3580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2311 net3572 vssd1 vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2322 _04276_ vssd1 vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3067 _03787_ vssd1 vssd1 vccd1 vccd1 net3591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2333 _01548_ vssd1 vssd1 vccd1 vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2344 _01281_ vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3089 _03888_ vssd1 vssd1 vccd1 vccd1 net3613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 net6875 vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2355 net6001 vssd1 vssd1 vccd1 vccd1 net2879 sky130_fd_sc_hd__clkbuf_2
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1621 _01469_ vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2366 _03545_ vssd1 vssd1 vccd1 vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1632 _03448_ vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2377 net6021 vssd1 vssd1 vccd1 vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 _04506_ vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2388 _03534_ vssd1 vssd1 vccd1 vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1654 _01309_ vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2399 _03541_ vssd1 vssd1 vccd1 vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1665 _04479_ vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1676 net6841 vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1687 _01437_ vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1698 _04232_ vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ net6397 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21707_ clknet_leaf_20_i_clk net5040 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ net42 _05604_ _05606_ net4077 vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a31o_1
XFILLER_0_212_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21638_ clknet_leaf_28_i_clk net6227 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12371_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _05230_ vssd1 vssd1 vccd1 vccd1 _05538_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21569_ clknet_leaf_16_i_clk net4997 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14110_ _07010_ _07021_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11322_ net6976 net6469 _04540_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
X_15090_ net3462 net3284 _08191_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ _06862_ net542 vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__nor2_1
X_11253_ net2866 net6375 _04503_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11184_ net2544 net6972 _04470_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__mux2_1
Xhold4280 net942 vssd1 vssd1 vccd1 vccd1 net4804 sky130_fd_sc_hd__dlygate4sd3_1
X_17800_ _01671_ _01726_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a21o_1
X_15992_ _09063_ _09066_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__or2_1
X_18780_ _04632_ _02767_ _02768_ _02773_ _02774_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a32o_1
Xhold3590 net602 vssd1 vssd1 vccd1 vccd1 net4114 sky130_fd_sc_hd__dlygate4sd3_1
X_17731_ _10379_ _09249_ _01780_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__o21ai_1
X_20741__172 clknet_1_0__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__inv_2
X_14943_ _06678_ _08035_ _08038_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17662_ _10302_ _01713_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14874_ _06625_ _08024_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__nand2_2
X_19401_ net1871 _03212_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__or2_1
X_16613_ _09551_ _09544_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__and2b_1
X_13825_ _06974_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xor2_2
X_17593_ _10477_ _10478_ _10476_ vssd1 vssd1 vccd1 vccd1 _10591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16544_ _09613_ _09615_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19332_ net1670 _03173_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or2_1
X_13756_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__nor2_1
X_10968_ net6514 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ net11 net12 net13 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a21oi_1
X_16475_ _09091_ _09251_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19263_ net5417 _03132_ _03135_ _03128_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__o211a_1
X_13687_ _06743_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__clkbuf_2
X_10899_ net7157 net2496 _04321_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
X_15426_ net3492 _06210_ _08309_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_66_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18214_ net3508 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__clkbuf_8
X_19194_ net1534 _03079_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12638_ clknet_leaf_69_i_clk _05785_ _05795_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__and3_2
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ net3102 _06210_ _08430_ _08431_ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__a2bb2o_2
X_18145_ _02190_ _02191_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__nor2_1
X_12569_ _04979_ _05721_ _05725_ _05028_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__o311a_1
XFILLER_0_171_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5909 net1206 vssd1 vssd1 vccd1 vccd1 net6433 sky130_fd_sc_hd__dlygate4sd3_1
X_14308_ _07432_ _07458_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18076_ _10257_ _09805_ _01991_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__o31a_1
Xhold206 _01119_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15288_ _08361_ _08342_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold217 net4461 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _01332_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ _10033_ _10034_ vssd1 vssd1 vccd1 vccd1 _10035_ sky130_fd_sc_hd__or2b_1
X_14239_ _07388_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__xnor2_2
Xhold239 net5006 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _09956_ _09949_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _01976_ net7798 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22472_ clknet_leaf_80_i_clk net4624 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21423_ clknet_leaf_85_i_clk net3199 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21354_ clknet_leaf_42_i_clk net4879 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold740 net5521 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
X_21285_ clknet_leaf_65_i_clk _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold751 net5050 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 net5553 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold773 net5620 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
X_20236_ net5432 _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or2_1
Xhold784 net5593 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 net5388 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799__224 clknet_1_0__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__inv_2
X_20167_ net5575 _03705_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or2_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2130 _04520_ vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2141 net7216 vssd1 vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2152 _01433_ vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2163 _04171_ vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20098_ net4797 net2630 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__nor2_1
Xhold2174 rbzero.tex_r1\[11\] vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2185 _04337_ vssd1 vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1440 net6659 vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 _01473_ vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2196 net2746 vssd1 vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ net4280 net4303 net4271 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor3_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1462 _04442_ vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1473 _01380_ vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1484 _04218_ vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _01436_ vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _05004_ _05038_ _05040_ _05010_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o211a_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13610_ _06759_ _06760_ _06676_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__o21a_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ net1760 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _07642_ _07689_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__nand2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ net5806 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16260_ _08564_ _08529_ _08471_ _08484_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__or4_1
X_20771__198 clknet_1_1__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__inv_2
X_13472_ _06614_ _06616_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__or3_1
X_10684_ net5983 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15211_ net3625 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__clkbuf_1
X_12423_ rbzero.tex_g1\[31\] rbzero.tex_g1\[30\] _05483_ vssd1 vssd1 vccd1 vccd1 _05590_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16191_ _08790_ _08804_ _08788_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15142_ _08246_ net4932 vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__nor2_1
X_12354_ _05514_ _05521_ _05022_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11305_ net7294 net6846 _04529_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15073_ net4689 net4687 _08191_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19950_ net4387 _03530_ net669 _03550_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__o211a_1
XFILLER_0_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12285_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _05071_ vssd1 vssd1 vccd1 vccd1 _05453_
+ sky130_fd_sc_hd__mux2_1
X_14024_ _07173_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__nor2_1
X_18901_ _02871_ _02884_ _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__a21oi_1
X_11236_ net2412 net5900 _04492_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__mux2_1
X_19881_ net2814 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__clkbuf_1
X_18832_ net4709 net7611 _02820_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__and3_1
X_11167_ net6441 net2578 _04459_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__mux2_1
X_18763_ net4799 net941 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15975_ net3539 _08313_ _08628_ _08430_ _09049_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__o41ai_2
X_11098_ net6666 net2128 _04426_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__mux2_1
X_17714_ _10257_ _09420_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14926_ net7433 _08062_ _08067_ _08073_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__a31o_2
XFILLER_0_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18694_ _02697_ _02698_ _02695_ _02696_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__04002_ clknet_0__04002_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04002_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17645_ _01695_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__nand2_1
X_14857_ net7908 _08007_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13808_ _06956_ _06958_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14788_ _07774_ _07590_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__nor2_1
X_17576_ net4403 net7373 vssd1 vssd1 vccd1 vccd1 _10574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19315_ net2487 _03160_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16527_ _09597_ _09598_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__nand2_1
X_13739_ _06844_ _06884_ _06886_ _06881_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246_ net5649 _03119_ _03125_ _03115_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__o211a_1
X_16458_ _09513_ _09514_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__or2_2
Xhold7108 rbzero.pov.ready_buffer\[2\] vssd1 vssd1 vccd1 vccd1 net7632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7119 rbzero.traced_texa\[6\] vssd1 vssd1 vccd1 vccd1 net7643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_144_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15409_ _08483_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__buf_2
X_16389_ _09445_ _09461_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__xnor2_1
Xhold6407 rbzero.tex_g0\[51\] vssd1 vssd1 vccd1 vccd1 net6931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19177_ _03038_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6418 net2373 vssd1 vssd1 vccd1 vccd1 net6942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6429 _04579_ vssd1 vssd1 vccd1 vccd1 net6953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5706 _03247_ vssd1 vssd1 vccd1 vccd1 net6230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18128_ _01984_ _02160_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5717 _02555_ vssd1 vssd1 vccd1 vccd1 net6241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5728 _01613_ vssd1 vssd1 vccd1 vccd1 net6252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5739 net1744 vssd1 vssd1 vccd1 vccd1 net6263 sky130_fd_sc_hd__dlygate4sd3_1
X_18059_ _02098_ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__xnor2_1
X_20748__178 clknet_1_0__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__inv_2
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21070_ _04063_ _04064_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ net3770 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21972_ net197 net2621 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer10 net533 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 net542 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xrebuffer32 _06827_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer43 _06857_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_1
Xrebuffer54 _06882_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer65 _07145_ vssd1 vssd1 vccd1 vccd1 net3163 sky130_fd_sc_hd__clkbuf_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22455_ clknet_leaf_40_i_clk _01624_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21406_ clknet_leaf_70_i_clk _00575_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22386_ net518 net2345 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6952 net4581 vssd1 vssd1 vccd1 vccd1 net7476 sky130_fd_sc_hd__clkbuf_4
Xhold6963 net4158 vssd1 vssd1 vccd1 vccd1 net7487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6974 net4182 vssd1 vssd1 vccd1 vccd1 net7498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21337_ clknet_leaf_46_i_clk net4154 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6996 net4298 vssd1 vssd1 vccd1 vccd1 net7520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20807__231 clknet_1_0__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__inv_2
XFILLER_0_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12070_ _05235_ _05236_ _05238_ _05034_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__o211a_1
Xhold570 net6380 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
X_21268_ clknet_leaf_50_i_clk _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold581 net5499 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _03206_ vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net6485 net2671 _04310_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__mux2_1
X_20219_ net5383 _03730_ _03734_ _03735_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__o211a_1
X_21199_ net4905 _02528_ _02579_ _04152_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a22o_1
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _08805_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__xnor2_4
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ net3876 net3085 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__or2_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 net6791 vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _05051_ _05092_ _04975_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a21bo_1
Xhold1281 _01113_ vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
X_14711_ _07232_ _07399_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1292 _04542_ vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _08752_ _08759_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__and2b_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _10428_ _10429_ vssd1 vssd1 vccd1 vccd1 _10430_ sky130_fd_sc_hd__nor2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14642_ _07740_ _07792_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__nor2_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11854_ _05013_ _05016_ _05020_ _05010_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a221o_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853__273 clknet_1_0__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__inv_2
X_10805_ net6830 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _09562_ _09312_ vssd1 vssd1 vccd1 vccd1 _10361_ sky130_fd_sc_hd__nor2_1
X_14573_ _07618_ _07438_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__or2_2
XFILLER_0_71_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ _04938_ _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19100_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__buf_2
X_16312_ _09383_ _09385_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__nor2_1
X_13524_ _06668_ _06630_ _06655_ _06674_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__or4_2
X_10736_ net5886 net5857 _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
X_17292_ _09593_ _10152_ vssd1 vssd1 vccd1 vccd1 _10293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16243_ _09315_ _09316_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__or2b_1
X_19031_ net3957 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__buf_4
X_13455_ _06604_ _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__xnor2_4
X_10667_ net2153 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12406_ _05177_ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16174_ net6148 _08299_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__nand2_4
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13386_ _06431_ _06135_ _06137_ _06536_ net4947 vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__a311o_1
X_10598_ net4049 vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__buf_4
X_15125_ net6150 _08223_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__or2_1
X_12337_ _05503_ _05504_ _04981_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19933_ net4358 _03530_ net2915 _03550_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__o211a_1
X_15056_ net4586 _08186_ _08138_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__mux2_1
X_12268_ net7427 _05383_ _05425_ rbzero.debug_overlay.playerX\[5\] _04807_ vssd1 vssd1
+ vccd1 vccd1 _05437_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14007_ _06865_ _06990_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nor2_1
X_11219_ _04332_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19864_ _03478_ net2928 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__or2_1
X_12199_ _05341_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__nor2_1
X_18815_ _02579_ _02801_ net4627 net3133 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19795_ net3100 _03442_ net1544 _03441_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ net3279 _02743_ _02261_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
X_15958_ _09010_ _09011_ _09032_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ net7568 _08057_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__nand2_1
X_18677_ _02682_ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__xnor2_1
X_15889_ _08958_ _08960_ _08963_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17628_ _01678_ _01679_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17559_ _10505_ _10557_ vssd1 vssd1 vccd1 vccd1 _10558_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20570_ _03924_ net3813 vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19229_ net5226 _03107_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__or2_1
Xhold6204 net2390 vssd1 vssd1 vccd1 vccd1 net6728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6215 rbzero.spi_registers.buf_texadd2\[3\] vssd1 vssd1 vccd1 vccd1 net6739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6226 net2188 vssd1 vssd1 vccd1 vccd1 net6750 sky130_fd_sc_hd__dlygate4sd3_1
X_22240_ net372 net1708 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold6237 _04206_ vssd1 vssd1 vccd1 vccd1 net6761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6248 net2304 vssd1 vssd1 vccd1 vccd1 net6772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5503 net2989 vssd1 vssd1 vccd1 vccd1 net6027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6259 rbzero.spi_registers.buf_texadd2\[18\] vssd1 vssd1 vccd1 vccd1 net6783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5514 _03456_ vssd1 vssd1 vccd1 vccd1 net6038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5525 net3987 vssd1 vssd1 vccd1 vccd1 net6049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22171_ net303 net2118 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold5536 net1844 vssd1 vssd1 vccd1 vccd1 net6060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4802 net1027 vssd1 vssd1 vccd1 vccd1 net5326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5547 net1670 vssd1 vssd1 vccd1 vccd1 net6071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5558 net3024 vssd1 vssd1 vccd1 vccd1 net6082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4813 rbzero.spi_registers.texadd3\[4\] vssd1 vssd1 vccd1 vccd1 net5337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4824 net976 vssd1 vssd1 vccd1 vccd1 net5348 sky130_fd_sc_hd__dlygate4sd3_1
X_21122_ net4176 net4744 vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__nand2_1
Xhold4835 rbzero.spi_registers.buf_vshift\[5\] vssd1 vssd1 vccd1 vccd1 net5359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4846 rbzero.spi_registers.buf_mapdy\[1\] vssd1 vssd1 vccd1 vccd1 net5370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4857 net946 vssd1 vssd1 vccd1 vccd1 net5381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4868 _00862_ vssd1 vssd1 vccd1 vccd1 net5392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4879 _00824_ vssd1 vssd1 vccd1 vccd1 net5403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21053_ _04048_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__xnor2_1
X_20004_ _03440_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ net180 net2610 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ clknet_leaf_98_i_clk net1390 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20357__87 clknet_1_0__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__inv_2
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _04714_ _04683_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13240_ net5706 _06179_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__xor2_1
X_22438_ clknet_leaf_39_i_clk net4746 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6760 net2668 vssd1 vssd1 vccd1 vccd1 net7284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _06318_ _06323_ _06325_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__and4bb_1
Xhold6771 rbzero.tex_g0\[54\] vssd1 vssd1 vccd1 vccd1 net7295 sky130_fd_sc_hd__dlygate4sd3_1
X_22369_ net501 net1450 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__04005_ clknet_0__04005_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04005_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6782 net2862 vssd1 vssd1 vccd1 vccd1 net7306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6793 rbzero.wall_hot\[1\] vssd1 vssd1 vccd1 vccd1 net7317 sky130_fd_sc_hd__dlygate4sd3_1
X_12122_ _05244_ _05286_ _05290_ _05023_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a211o_1
X_20883__299 clknet_1_1__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__inv_2
XFILLER_0_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12053_ _05002_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__or2_1
X_16930_ _06229_ _09294_ vssd1 vssd1 vccd1 vccd1 _09948_ sky130_fd_sc_hd__xnor2_2
X_11004_ net6960 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__clkbuf_1
X_16861_ net4074 _09920_ vssd1 vssd1 vccd1 vccd1 _09923_ sky130_fd_sc_hd__and2_1
X_18600_ _02590_ _02591_ net3838 _02569_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__o2bb2a_1
X_15812_ _08881_ _08880_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19580_ net5279 _03302_ _03322_ _03314_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__o211a_1
X_16792_ _09139_ _09861_ vssd1 vssd1 vccd1 vccd1 _09862_ sky130_fd_sc_hd__nor2_1
X_18531_ _05403_ net4424 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__or2_1
X_15743_ _08758_ _08809_ _08816_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__a21o_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__xor2_2
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ _05062_ _05066_ _05075_ _04979_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a211o_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18462_ net3062 _02485_ _02331_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__o21ai_1
X_15674_ _08747_ _08748_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__or2_4
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ net4083 _06000_ _06006_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__o22a_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17413_ _10405_ _10412_ vssd1 vssd1 vccd1 vccd1 _10413_ sky130_fd_sc_hd__xnor2_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _04983_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14625_ _07232_ _06918_ _07464_ _07438_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__or4_4
X_18393_ net4487 net4423 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _10278_ _10254_ vssd1 vssd1 vccd1 vccd1 _10344_ sky130_fd_sc_hd__or2b_1
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14556_ _07366_ _07523_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nor2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _04934_ _04936_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03982_ clknet_0__03982_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03982_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ net2699 net5976 _04225_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux2_1
X_13507_ _06626_ _06649_ _06656_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__o21ai_2
X_17275_ _10255_ _10256_ _10275_ vssd1 vssd1 vccd1 vccd1 _10276_ sky130_fd_sc_hd__a21o_1
X_14487_ _07585_ _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__nor2_1
X_11699_ net2043 _04600_ _04602_ _04868_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19014_ net3374 _02979_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__or2_1
X_16226_ _09184_ _09275_ _09273_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_181_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13438_ _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer1 net526 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16157_ _08612_ net7444 _09231_ _08620_ _08603_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__o32a_1
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13369_ net4406 net4787 vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4109 net858 vssd1 vssd1 vccd1 vccd1 net4633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _08218_ net3187 net6260 _08215_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__o211a_1
X_16088_ _09137_ _09142_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__nor2_1
Xhold3408 rbzero.spi_registers.spi_buffer\[3\] vssd1 vssd1 vccd1 vccd1 net3932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3419 _00633_ vssd1 vssd1 vccd1 vccd1 net3943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ net4368 _08173_ _08138_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__mux2_1
X_19916_ _03531_ _03538_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2707 _03825_ vssd1 vssd1 vccd1 vccd1 net3231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2718 _02572_ vssd1 vssd1 vccd1 vccd1 net3242 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2729 _01248_ vssd1 vssd1 vccd1 vccd1 net3253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19847_ _08342_ _08343_ _03485_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o21a_1
XFILLER_0_208_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19778_ net6263 _03429_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ net3919 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21740_ clknet_leaf_24_i_clk net2535 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21671_ clknet_leaf_13_i_clk net825 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20622_ net3898 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20553_ net733 net3488 _03911_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6001 _03259_ vssd1 vssd1 vccd1 vccd1 net6525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6012 _04559_ vssd1 vssd1 vccd1 vccd1 net6536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6023 net1518 vssd1 vssd1 vccd1 vccd1 net6547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6034 rbzero.spi_registers.buf_floor\[2\] vssd1 vssd1 vccd1 vccd1 net6558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20484_ net3521 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
Xhold6045 rbzero.tex_g0\[3\] vssd1 vssd1 vccd1 vccd1 net6569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5300 rbzero.tex_r1\[58\] vssd1 vssd1 vccd1 vccd1 net5824 sky130_fd_sc_hd__dlygate4sd3_1
X_22223_ net355 net1447 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
Xhold6056 net1552 vssd1 vssd1 vccd1 vccd1 net6580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5311 _04420_ vssd1 vssd1 vccd1 vccd1 net5835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5322 net2397 vssd1 vssd1 vccd1 vccd1 net5846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6067 rbzero.tex_b0\[41\] vssd1 vssd1 vccd1 vccd1 net6591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5333 rbzero.tex_r1\[4\] vssd1 vssd1 vccd1 vccd1 net5857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6078 net1652 vssd1 vssd1 vccd1 vccd1 net6602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5344 rbzero.tex_b1\[42\] vssd1 vssd1 vccd1 vccd1 net5868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6089 rbzero.tex_b0\[53\] vssd1 vssd1 vccd1 vccd1 net6613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4610 net802 vssd1 vssd1 vccd1 vccd1 net5134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5355 net2097 vssd1 vssd1 vccd1 vccd1 net5879 sky130_fd_sc_hd__dlygate4sd3_1
X_22154_ net286 net2580 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
Xhold5366 net1874 vssd1 vssd1 vccd1 vccd1 net5890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4621 net903 vssd1 vssd1 vccd1 vccd1 net5145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5377 _04501_ vssd1 vssd1 vccd1 vccd1 net5901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4632 _00839_ vssd1 vssd1 vccd1 vccd1 net5156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5388 _04313_ vssd1 vssd1 vccd1 vccd1 net5912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4643 rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 net5167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5399 rbzero.tex_b0\[2\] vssd1 vssd1 vccd1 vccd1 net5923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4654 net870 vssd1 vssd1 vccd1 vccd1 net5178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ _04093_ _04094_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a21o_1
Xhold3920 _00987_ vssd1 vssd1 vccd1 vccd1 net4444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4665 rbzero.spi_registers.buf_mapdx\[1\] vssd1 vssd1 vccd1 vccd1 net5189 sky130_fd_sc_hd__dlygate4sd3_1
X_22085_ clknet_leaf_74_i_clk net4019 vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold3931 net3217 vssd1 vssd1 vccd1 vccd1 net4455 sky130_fd_sc_hd__buf_1
Xhold4676 rbzero.spi_registers.buf_texadd0\[7\] vssd1 vssd1 vccd1 vccd1 net5200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3942 net7523 vssd1 vssd1 vccd1 vccd1 net4466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4687 rbzero.pov.spi_buffer\[43\] vssd1 vssd1 vccd1 vccd1 net5211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3953 _02539_ vssd1 vssd1 vccd1 vccd1 net4477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4698 net849 vssd1 vssd1 vccd1 vccd1 net5222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3964 net7529 vssd1 vssd1 vccd1 vccd1 net4488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3975 net3369 vssd1 vssd1 vccd1 vccd1 net4499 sky130_fd_sc_hd__buf_1
X_21036_ net5168 _03519_ _04014_ _04037_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a22o_1
Xhold3986 net7539 vssd1 vssd1 vccd1 vccd1 net4510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3997 _03586_ vssd1 vssd1 vccd1 vccd1 net4521 sky130_fd_sc_hd__dlygate4sd3_1
X_20919__332 clknet_1_0__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__inv_2
XFILLER_0_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ net4095 _05446_ net16 vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__mux2_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21938_ clknet_leaf_9_i_clk net1303 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _04162_ net3993 net4 vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ clknet_leaf_100_i_clk net1171 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14410_ _07546_ _07560_ _07558_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _04614_ _04790_ _04160_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21oi_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15390_ _08464_ net4358 _06178_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14341_ _07473_ _07489_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__a21bo_1
X_11553_ _04714_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17060_ _10062_ _10063_ _10064_ vssd1 vssd1 vccd1 vccd1 _10065_ sky130_fd_sc_hd__o21ai_1
X_14272_ _07418_ _07421_ _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11484_ rbzero.texu_hot\[2\] _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nand2_1
X_16011_ _08560_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7280 rbzero.wall_tracer.stepDistY\[-10\] vssd1 vssd1 vccd1 vccd1 net7804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ _06364_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__inv_2
X_20965__374 clknet_1_0__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__inv_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7291 _02077_ vssd1 vssd1 vccd1 vccd1 net7815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20664__102 clknet_1_1__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__inv_2
Xhold6590 rbzero.tex_r0\[8\] vssd1 vssd1 vccd1 vccd1 net7114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13154_ _06308_ net3233 _06309_ net3221 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12105_ _05268_ _05270_ _05273_ _05010_ _04978_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a221o_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17962_ _01890_ _01899_ _01897_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a21oi_1
X_13085_ net2388 net2907 net1130 net1064 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__or4_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19701_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__buf_2
X_16913_ _09935_ vssd1 vssd1 vccd1 vccd1 _09942_ sky130_fd_sc_hd__clkbuf_4
X_12036_ _05205_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17893_ _01936_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19632_ net4401 _03326_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or2_1
X_16844_ net7368 _08296_ _09912_ _09913_ _08195_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19563_ _03294_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__clkbuf_4
X_16775_ _09843_ _09844_ vssd1 vssd1 vccd1 vccd1 _09845_ sky130_fd_sc_hd__xor2_1
X_13987_ _07120_ _07134_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__and2b_1
X_18514_ _05403_ net715 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__nand2_1
X_15726_ _08799_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ net6294 _03266_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ net3876 net3018 vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__or2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18445_ _02460_ _02463_ _02461_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__o21ai_1
X_15657_ _08394_ _08471_ _08484_ _08411_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__o22ai_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ net4972 _05998_ _06007_ net4002 vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ _07471_ _07590_ _07754_ _07758_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__o31a_1
XFILLER_0_84_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18376_ net4920 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__buf_4
X_15588_ _06209_ _08613_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__nand2_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17327_ _10202_ _10204_ _10327_ vssd1 vssd1 vccd1 vccd1 _10328_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14539_ _07642_ _07689_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17258_ _08315_ vssd1 vssd1 vccd1 vccd1 _10259_ sky130_fd_sc_hd__buf_2
Xclkbuf_0__03996_ _03996_ vssd1 vssd1 vccd1 vccd1 clknet_0__03996_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16209_ _09178_ _09180_ vssd1 vssd1 vccd1 vccd1 _09284_ sky130_fd_sc_hd__xor2_4
XFILLER_0_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17189_ _10189_ _10190_ vssd1 vssd1 vccd1 vccd1 _10191_ sky130_fd_sc_hd__xor2_2
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3205 _03837_ vssd1 vssd1 vccd1 vccd1 net3729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3216 _01179_ vssd1 vssd1 vccd1 vccd1 net3740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3227 rbzero.pov.spi_buffer\[65\] vssd1 vssd1 vccd1 vccd1 net3751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3238 _05355_ vssd1 vssd1 vccd1 vccd1 net3762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2504 net6198 vssd1 vssd1 vccd1 vccd1 net3028 sky130_fd_sc_hd__clkbuf_4
Xhold3249 net6147 vssd1 vssd1 vccd1 vccd1 net3773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _00640_ vssd1 vssd1 vccd1 vccd1 net3039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2526 net6163 vssd1 vssd1 vccd1 vccd1 net3050 sky130_fd_sc_hd__clkbuf_2
Xhold2537 _02483_ vssd1 vssd1 vccd1 vccd1 net3061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1803 _01399_ vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 net6028 vssd1 vssd1 vccd1 vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1814 _04246_ vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2559 _03572_ vssd1 vssd1 vccd1 vccd1 net3083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1825 net6755 vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1836 net6843 vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1847 _04594_ vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 rbzero.tex_r1\[6\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 net5885 vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21723_ clknet_leaf_4_i_clk net2489 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21654_ clknet_leaf_16_i_clk net5112 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_otherx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20605_ net4014 net3965 vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21585_ clknet_leaf_21_i_clk net4193 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20536_ _08274_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_99 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_99/HI o_rgb[11] sky130_fd_sc_hd__conb_1
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20350__82 clknet_1_0__leaf__03779_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__inv_2
X_20467_ _03836_ net3710 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2_1
Xhold5130 net1331 vssd1 vssd1 vccd1 vccd1 net5654 sky130_fd_sc_hd__dlygate4sd3_1
X_22206_ net338 net2540 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
Xhold5141 net1400 vssd1 vssd1 vccd1 vccd1 net5665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5152 net1405 vssd1 vssd1 vccd1 vccd1 net5676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5163 rbzero.pov.spi_buffer\[35\] vssd1 vssd1 vccd1 vccd1 net5687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20398_ net3686 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5174 rbzero.map_overlay.i_mapdx\[4\] vssd1 vssd1 vccd1 vccd1 net5698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5185 rbzero.floor_leak\[2\] vssd1 vssd1 vccd1 vccd1 net5709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4440 gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4964 sky130_fd_sc_hd__dlygate4sd3_1
X_22137_ net269 net2175 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
Xhold4451 net707 vssd1 vssd1 vccd1 vccd1 net4975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5196 rbzero.spi_registers.vshift\[1\] vssd1 vssd1 vccd1 vccd1 net5720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4462 rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 net4986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4473 net754 vssd1 vssd1 vccd1 vccd1 net4997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4484 _00748_ vssd1 vssd1 vccd1 vccd1 net5008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3750 net7846 vssd1 vssd1 vccd1 vccd1 net4274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4495 _00794_ vssd1 vssd1 vccd1 vccd1 net5019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3761 rbzero.wall_tracer.visualWallDist\[2\] vssd1 vssd1 vccd1 vccd1 net4285 sky130_fd_sc_hd__clkbuf_1
X_22068_ clknet_leaf_8_i_clk net3708 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3772 net2992 vssd1 vssd1 vccd1 vccd1 net4296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3783 _00956_ vssd1 vssd1 vccd1 vccd1 net4307 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03985_ clknet_0__03985_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03985_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3794 net4321 vssd1 vssd1 vccd1 vccd1 net4318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21019_ _04020_ _04021_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__and2_1
X_13910_ _06948_ _06949_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__xnor2_2
X_14890_ net7434 _08011_ vssd1 vssd1 vccd1 vccd1 _08040_ sky130_fd_sc_hd__nor2_1
X_13841_ _06989_ _06991_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16560_ _09506_ _09507_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13772_ _06860_ _06864_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__xnor2_4
X_10984_ net6636 net6876 _04366_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15511_ _08583_ _08585_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12723_ clknet_1_1__leaf__04800_ _05843_ _05854_ vssd1 vssd1 vccd1 vccd1 _05884_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16491_ _08316_ _09562_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18230_ _02190_ _02193_ _02191_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__o21bai_1
X_15442_ _08501_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ net4034 vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__buf_4
XFILLER_0_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18161_ _08634_ _09420_ _09538_ _08643_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__o22a_1
X_12585_ _05004_ _05749_ _05461_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__o21a_1
X_15373_ _08405_ _08411_ _08422_ _08432_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17112_ _10112_ _10113_ vssd1 vssd1 vccd1 vccd1 _10114_ sky130_fd_sc_hd__nand2_1
X_14324_ _07474_ _07439_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11536_ rbzero.spi_registers.texadd2\[23\] _04642_ _04644_ rbzero.spi_registers.texadd1\[23\]
+ _04707_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a221o_1
X_18092_ _02129_ _02139_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03781_ _03781_ vssd1 vssd1 vccd1 vccd1 clknet_0__03781_ sky130_fd_sc_hd__clkbuf_16
X_17043_ _10049_ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__clkbuf_1
X_14255_ _07362_ _07397_ _07395_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11467_ net6496 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _06222_ _06186_ net3804 _06217_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__a22o_1
X_14186_ _07274_ _07309_ _07336_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__a21o_1
X_11398_ net7219 net6333 _04584_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ net3462 _06276_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__and2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18994_ net3213 net2978 net3747 vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _10130_ _09805_ _01881_ _01880_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__o31a_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ net2895 _06221_ _06213_ net2825 _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12019_ _04858_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__inv_2
X_17876_ _01809_ _01810_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19615_ net969 net799 _03344_ _03343_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__o211a_1
X_16827_ _09895_ _09896_ vssd1 vssd1 vccd1 vccd1 _09897_ sky130_fd_sc_hd__xor2_2
X_19546_ _02491_ _02497_ _02500_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nand3_2
X_16758_ _09826_ _09827_ vssd1 vssd1 vccd1 vccd1 _09828_ sky130_fd_sc_hd__nand2_1
X_15709_ _08781_ _08783_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_193_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19477_ _03141_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__clkbuf_4
X_16689_ _09757_ _09758_ vssd1 vssd1 vccd1 vccd1 _09760_ sky130_fd_sc_hd__and2_1
X_18428_ _02454_ _02455_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18359_ _02394_ _02395_ _10064_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21370_ clknet_leaf_59_i_clk _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold900 net6488 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 net6538 vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 net6486 vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold933 net4543 vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_20252_ net3568 _03743_ _03753_ _03748_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__o211a_1
Xhold944 _02991_ vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 _01477_ vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 _01459_ vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 net6480 vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3002 _03940_ vssd1 vssd1 vccd1 vccd1 net3526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3013 net4592 vssd1 vssd1 vccd1 vccd1 net3537 sky130_fd_sc_hd__buf_1
Xhold988 net6550 vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20183_ net3557 _03704_ net5482 _03709_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__o211a_1
Xhold3024 _03841_ vssd1 vssd1 vccd1 vccd1 net3548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 _01110_ vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3035 _03844_ vssd1 vssd1 vccd1 vccd1 net3559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3046 _03910_ vssd1 vssd1 vccd1 vccd1 net3570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2301 net5949 vssd1 vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__clkbuf_2
Xhold3057 _03892_ vssd1 vssd1 vccd1 vccd1 net3581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2312 _03535_ vssd1 vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2323 _01493_ vssd1 vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3068 _03788_ vssd1 vssd1 vccd1 vccd1 net3592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2334 net7267 vssd1 vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3079 _02615_ vssd1 vssd1 vccd1 vccd1 net3603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1600 _00654_ vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
X_20801__226 clknet_1_0__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__inv_2
Xhold2345 net7888 vssd1 vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__buf_2
Xhold1611 _04369_ vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2356 net6003 vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 net6845 vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2367 net6128 vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 net7308 vssd1 vssd1 vccd1 vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _00939_ vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1644 _01286_ vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2389 net4356 vssd1 vssd1 vccd1 vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1655 net2411 vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1666 _01310_ vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1677 _04476_ vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1688 net7118 vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1699 _01530_ vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21706_ clknet_leaf_20_i_clk net5097 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21637_ clknet_leaf_32_i_clk net3107 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _05457_ vssd1 vssd1 vccd1 vccd1 _05537_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21568_ clknet_leaf_16_i_clk net5024 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ net2503 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20519_ _03880_ net3276 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21499_ clknet_leaf_13_i_clk net2826 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _07185_ _07190_ _07156_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__or3b_4
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ net1801 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ net2323 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4270 net4836 vssd1 vssd1 vccd1 vccd1 net4794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4281 rbzero.wall_tracer.rayAddendX\[-7\] vssd1 vssd1 vccd1 vccd1 net4805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4292 _02906_ vssd1 vssd1 vccd1 vccd1 net4816 sky130_fd_sc_hd__dlygate4sd3_1
X_15991_ _09005_ _09065_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__or2_1
X_17730_ _10379_ _09249_ _01780_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__or3_1
Xhold3580 _04620_ vssd1 vssd1 vccd1 vccd1 net4104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3591 net7620 vssd1 vssd1 vccd1 vccd1 net4115 sky130_fd_sc_hd__dlygate4sd3_1
X_14942_ _08030_ _08032_ net7843 vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__a21o_1
X_20776__203 clknet_1_0__leaf__03991_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__inv_2
X_17661_ _09593_ _01712_ _10543_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
Xhold2890 _03862_ vssd1 vssd1 vccd1 vccd1 net3414 sky130_fd_sc_hd__dlygate4sd3_1
X_14873_ net7566 _08005_ _08023_ _06589_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__a211o_1
X_19400_ net5435 _03211_ _03213_ _03207_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16612_ _09672_ _09682_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__xnor2_1
X_13824_ _06889_ _06837_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__nor2_1
X_17592_ _10588_ _10589_ vssd1 vssd1 vccd1 vccd1 _10590_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ net5660 _03172_ _03174_ _03168_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__o211a_1
X_16543_ _09485_ _09491_ _09614_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__a21o_1
X_10967_ net2765 net6512 _04355_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__mux2_1
X_13755_ _06903_ _06904_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19262_ net5061 _03133_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or2_1
X_12706_ net4060 _05853_ _05854_ _05816_ _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a221o_1
X_16474_ _08724_ _09251_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__nor2_1
X_10898_ net7306 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13686_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18213_ _02258_ _02259_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__xnor2_1
X_15425_ _08486_ _08499_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19193_ net5356 _03078_ _03094_ _03074_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__o211a_1
X_12637_ net5 net4 vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__and2_2
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18144_ _01684_ _10520_ _01711_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__nor3_1
X_12568_ _05000_ _05728_ _05730_ _05732_ _05023_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a221o_1
X_15356_ net4382 _08379_ _08311_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ _07446_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__xnor2_1
X_11519_ _04689_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_145_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18075_ _01989_ _01990_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__nand2_1
X_12499_ _05663_ _05664_ _05235_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15287_ _08361_ _08342_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__nand2_1
Xhold207 net3316 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 net5010 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ net4556 net4719 vssd1 vssd1 vccd1 vccd1 _10034_ sky130_fd_sc_hd__nand2_1
Xhold229 net4994 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _07325_ _07334_ _07332_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ net568 _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ net3985 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _01865_ _01868_ _01866_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__o21a_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17859_ _01877_ _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19529_ _02996_ _03289_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22471_ clknet_leaf_81_i_clk net4441 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21422_ clknet_leaf_85_i_clk net4789 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21353_ clknet_leaf_35_i_clk net3220 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold730 net4852 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
X_21284_ clknet_leaf_64_i_clk _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold741 net5587 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 net5581 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 net5555 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
X_20235_ _03678_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold774 net7652 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold785 net5595 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 net5648 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20725__157 clknet_1_1__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__inv_2
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ _03678_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__buf_2
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2120 net7162 vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2131 _01273_ vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2142 _04438_ vssd1 vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2153 net5907 vssd1 vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__clkbuf_2
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2164 _01586_ vssd1 vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
X_20097_ net2629 net4796 _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__a21bo_1
Xhold2175 net2259 vssd1 vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1430 _04248_ vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2186 _01439_ vssd1 vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1441 _03436_ vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2197 _04316_ vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1452 net7078 vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1463 _01344_ vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1474 _06626_ vssd1 vssd1 vccd1 vccd1 net3457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_212_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 _01543_ vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _04983_ _05039_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__or2_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1496 net6783 vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10821_ net6744 net6604 _04277_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10752_ net5804 net1932 _04244_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__mux2_1
X_13540_ _06667_ _06675_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13471_ _06619_ _06621_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10683_ net5914 net5981 _04203_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12422_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _05541_ vssd1 vssd1 vccd1 vccd1 _05589_
+ sky130_fd_sc_hd__mux2_1
X_15210_ _08195_ net3624 vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _09247_ _09264_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _05517_ _05520_ net80 vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15141_ net4909 net2982 net4027 net4931 vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__or4b_1
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ net7040 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15072_ _08190_ _08196_ net3540 _01622_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__o211a_1
X_12284_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _05219_ vssd1 vssd1 vccd1 vccd1 _05452_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18900_ _02867_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__xnor2_1
X_14023_ _07168_ _07172_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__xnor2_1
X_11235_ net5964 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
X_19880_ _04597_ net2813 _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__or3_1
X_18831_ net4709 _02819_ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a21o_1
X_11166_ net2566 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18762_ _02751_ _02756_ _02757_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__o21a_1
X_15974_ _08409_ _08664_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__or2_1
X_11097_ net2528 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17713_ _01697_ _01672_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__or2b_1
X_14925_ _08068_ _08072_ net6162 vssd1 vssd1 vccd1 vccd1 _08073_ sky130_fd_sc_hd__a21o_1
X_18693_ _02695_ _02696_ _02697_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a211o_1
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 net5837 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_2
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__04001_ clknet_0__04001_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04001_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _01673_ _01674_ _01694_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nand3_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _07695_ _07971_ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__xor2_2
XFILLER_0_202_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ _06737_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_212_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17575_ _10573_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14787_ _07618_ _07805_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__nor2_1
X_11999_ net2955 _04598_ _04602_ _05160_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a221o_1
X_19314_ net5083 _03159_ _03164_ _03155_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__o211a_1
X_16526_ _09139_ _09595_ _09596_ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _06826_ _06888_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19245_ net5391 _03120_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or2_1
X_16457_ _09518_ _09520_ _09516_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__o21a_1
X_13669_ _06707_ _06696_ _06700_ _06662_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7109 rbzero.traced_texa\[-2\] vssd1 vssd1 vccd1 vccd1 net7633 sky130_fd_sc_hd__dlygate4sd3_1
X_20830__252 clknet_1_0__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__inv_2
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ _08477_ _08478_ _08482_ _08327_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__a22o_2
X_19176_ _04597_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__clkbuf_8
X_16388_ _09451_ _09460_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__xor2_2
XFILLER_0_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6408 net1950 vssd1 vssd1 vccd1 vccd1 net6932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6419 rbzero.tex_r0\[33\] vssd1 vssd1 vccd1 vccd1 net6943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18127_ _02157_ _02159_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__or2_1
X_15339_ _08412_ _08413_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__and2_1
Xhold5707 _00805_ vssd1 vssd1 vccd1 vccd1 net6231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5718 _02558_ vssd1 vssd1 vccd1 vccd1 net6242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5729 net692 vssd1 vssd1 vccd1 vccd1 net6253 sky130_fd_sc_hd__buf_2
X_18058_ _02103_ _02105_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17009_ _06204_ vssd1 vssd1 vccd1 vccd1 _10019_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20020_ _03261_ net3769 vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21971_ net196 net1896 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer11 _07103_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 _06896_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer33 net556 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_1
Xrebuffer44 net567 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__dlygate4sd2_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer55 _06882_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer66 _07114_ vssd1 vssd1 vccd1 vccd1 net3203 sky130_fd_sc_hd__clkbuf_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22454_ clknet_leaf_40_i_clk _01623_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21405_ clknet_leaf_29_i_clk net3215 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6920 net7945 vssd1 vssd1 vccd1 vccd1 net7444 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22385_ net517 net1776 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold6953 _08329_ vssd1 vssd1 vccd1 vccd1 net7477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6964 rbzero.wall_tracer.stepDistY\[1\] vssd1 vssd1 vccd1 vccd1 net7488 sky130_fd_sc_hd__dlygate4sd3_1
X_21336_ clknet_leaf_50_i_clk net5312 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6975 rbzero.traced_texVinit\[5\] vssd1 vssd1 vccd1 vccd1 net7499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6986 _08348_ vssd1 vssd1 vccd1 vccd1 net7510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6997 rbzero.wall_tracer.trackDistY\[8\] vssd1 vssd1 vccd1 vccd1 net7521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21267_ clknet_leaf_58_i_clk _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold560 _03177_ vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold571 _01352_ vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net1983 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold582 net5501 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
X_20218_ _08275_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold593 net4195 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21198_ _02756_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__xor2_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ _03440_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__clkbuf_4
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _06122_ _06126_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__nand2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1260 net1406 vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1271 net6793 vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _07618_ _07359_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__nor2_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _05084_ _05091_ _05023_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__mux2_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 net6255 vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 _01160_ vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ _08763_ _08764_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__xnor2_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _07790_ _07791_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__and2_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__clkbuf_8
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ net6828 net2644 _04266_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__mux2_1
X_17360_ _10236_ _10357_ _10359_ vssd1 vssd1 vccd1 vccd1 _10360_ sky130_fd_sc_hd__a21oi_1
X_11784_ _04937_ _04934_ _04936_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__and3_1
X_14572_ _06865_ _07467_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__nand2_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _09215_ _09237_ _09384_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__a21oi_2
X_20888__304 clknet_1_0__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__inv_2
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13523_ _06567_ _06565_ _06587_ _06671_ _06673_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__a41o_1
X_10735_ _04169_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__clkbuf_4
X_17291_ _10290_ _10291_ vssd1 vssd1 vccd1 vccd1 _10292_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19030_ net1608 _02988_ _02995_ _02993_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__o211a_1
X_16242_ _09188_ _09303_ _09314_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ net2518 net5811 _04192_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13454_ _06560_ _06593_ _06429_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12405_ rbzero.tex_g1\[9\] rbzero.tex_g1\[8\] _05476_ vssd1 vssd1 vccd1 vccd1 _05572_
+ sky130_fd_sc_hd__mux2_1
X_16173_ _08744_ _08722_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13385_ net7476 _06431_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ net4558 net4573 _08219_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__mux2_1
X_12336_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _05493_ vssd1 vssd1 vccd1 vccd1 _05504_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19932_ _03440_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__clkbuf_4
X_12267_ net3853 _05368_ _05347_ net3995 _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a221o_1
X_15055_ _08150_ _08149_ _08047_ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11218_ net1810 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
X_14006_ _07115_ _07116_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19863_ net2927 _08441_ _03484_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
X_12198_ _05348_ _05361_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ net5922 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
X_18814_ _04633_ _02804_ _02805_ _09933_ rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a32o_1
XFILLER_0_207_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19794_ net6549 _03443_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18745_ _06197_ _06195_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__xnor2_1
X_15957_ _09012_ _09030_ _09031_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ _06838_ _08054_ _08056_ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__a21o_1
X_18676_ _02650_ _02668_ _02670_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a21o_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _08962_ _08665_ _08917_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17627_ _08643_ _08708_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nor2_1
X_14839_ _06690_ _07989_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17558_ _10555_ _10556_ vssd1 vssd1 vccd1 vccd1 _10557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16509_ _09560_ _09580_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__xnor2_2
X_17489_ _10358_ _10487_ vssd1 vssd1 vccd1 vccd1 _10488_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19228_ net5788 _03106_ _03114_ _03115_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6205 rbzero.spi_registers.buf_texadd1\[6\] vssd1 vssd1 vccd1 vccd1 net6729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6216 net1868 vssd1 vssd1 vccd1 vccd1 net6740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6227 rbzero.tex_g1\[42\] vssd1 vssd1 vccd1 vccd1 net6751 sky130_fd_sc_hd__dlygate4sd3_1
X_19159_ net5279 _03066_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__or2_1
Xhold6238 net1775 vssd1 vssd1 vccd1 vccd1 net6762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6249 _04268_ vssd1 vssd1 vccd1 vccd1 net6773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5504 rbzero.spi_registers.spi_buffer\[17\] vssd1 vssd1 vccd1 vccd1 net6028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5515 _00946_ vssd1 vssd1 vccd1 vccd1 net6039 sky130_fd_sc_hd__dlygate4sd3_1
X_22170_ net302 net1717 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold5526 rbzero.spi_registers.buf_texadd3\[22\] vssd1 vssd1 vccd1 vccd1 net6050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5537 rbzero.spi_registers.buf_texadd1\[21\] vssd1 vssd1 vccd1 vccd1 net6061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4803 _00696_ vssd1 vssd1 vccd1 vccd1 net5327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5548 _03389_ vssd1 vssd1 vccd1 vccd1 net6072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4814 net1025 vssd1 vssd1 vccd1 vccd1 net5338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21121_ net4176 net4744 vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__nor2_1
Xhold5559 _00971_ vssd1 vssd1 vccd1 vccd1 net6083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4825 rbzero.spi_registers.buf_texadd0\[14\] vssd1 vssd1 vccd1 vccd1 net5349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4836 net962 vssd1 vssd1 vccd1 vccd1 net5360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4847 net993 vssd1 vssd1 vccd1 vccd1 net5371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4858 rbzero.pov.spi_buffer\[42\] vssd1 vssd1 vccd1 vccd1 net5382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21052_ _04049_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__and2b_1
Xhold4869 net1046 vssd1 vssd1 vccd1 vccd1 net5393 sky130_fd_sc_hd__dlygate4sd3_1
X_20003_ rbzero.debug_overlay.facingY\[-8\] _03582_ vssd1 vssd1 vccd1 vccd1 _03601_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ net179 net1949 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837__258 clknet_1_1__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__inv_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ clknet_leaf_98_i_clk net5542 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22437_ clknet_leaf_38_i_clk net4655 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6750 net2740 vssd1 vssd1 vccd1 vccd1 net7274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13170_ _06324_ net3314 _06316_ net3460 vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__o2bb2a_1
Xhold6761 rbzero.tex_g1\[11\] vssd1 vssd1 vccd1 vccd1 net7285 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__04004_ clknet_0__04004_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04004_
+ sky130_fd_sc_hd__clkbuf_16
X_22368_ net500 net2730 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6772 net2897 vssd1 vssd1 vccd1 vccd1 net7296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ _05019_ _05287_ _05289_ _05009_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6783 gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 net7307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6794 _04638_ vssd1 vssd1 vccd1 vccd1 net7318 sky130_fd_sc_hd__dlygate4sd3_1
X_21319_ clknet_leaf_72_i_clk _00488_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22299_ net431 net1432 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
X_12052_ rbzero.tex_r1\[49\] rbzero.tex_r1\[48\] _05071_ vssd1 vssd1 vccd1 vccd1 _05221_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold390 net4807 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net2599 net6958 _04377_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
X_16860_ net4039 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__clkbuf_1
X_15811_ _08837_ _08885_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__xnor2_2
X_20993__19 clknet_1_0__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
X_16791_ _09603_ vssd1 vssd1 vccd1 vccd1 _09861_ sky130_fd_sc_hd__clkbuf_4
X_18530_ _05403_ net4424 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__nand2_1
X_15742_ _08758_ _08809_ _08816_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__nand3_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__or2_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 net5764 vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _05004_ _05067_ _05074_ _05035_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__o211a_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18461_ net4332 net3061 _01870_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a21o_1
X_15673_ _08695_ _08680_ _08694_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__a21oi_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _06019_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__or2_2
XFILLER_0_201_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ _10410_ _10411_ vssd1 vssd1 vccd1 vccd1 _10412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _07439_ _07774_ _07090_ _07466_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11836_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _04988_ vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__mux2_1
X_18392_ _02424_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17343_ _10234_ _10248_ _10246_ vssd1 vssd1 vccd1 vccd1 _10343_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14555_ _07367_ _07358_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__or2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03981_ clknet_0__03981_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03981_
+ sky130_fd_sc_hd__clkbuf_16
X_11767_ net2776 _04931_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13506_ _06626_ _06649_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__or3_4
X_17274_ _10264_ _10274_ vssd1 vssd1 vccd1 vccd1 _10275_ sky130_fd_sc_hd__xnor2_1
X_10718_ net5929 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__clkbuf_1
X_14486_ _07586_ _07633_ _07636_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ net2917 vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__inv_2
X_19013_ net3969 _02979_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__and2_1
X_16225_ net4376 _08296_ _09298_ _09299_ _08239_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__o221a_1
X_13437_ _06557_ _06565_ _06567_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__and4b_2
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ net2224 net6564 _04181_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__mux2_1
Xrebuffer2 _07110_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ _06211_ _08618_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__nand2_4
Xclkbuf_leaf_41_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13368_ _06471_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__xor2_2
X_15107_ net6259 _08223_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__or2_1
X_12319_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _05262_ vssd1 vssd1 vccd1 vccd1 _05487_
+ sky130_fd_sc_hd__mux2_1
X_16087_ _09156_ _09159_ _09160_ _09161_ vssd1 vssd1 vccd1 vccd1 _09162_ sky130_fd_sc_hd__o211a_1
X_13299_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__or2_1
X_20942__353 clknet_1_0__leaf__04007_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__inv_2
Xhold3409 net3123 vssd1 vssd1 vccd1 vccd1 net3933 sky130_fd_sc_hd__dlygate4sd3_1
X_19915_ net3713 _08356_ _03484_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_1
X_15038_ _06589_ _08172_ _08047_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__a21o_2
Xhold2708 _01193_ vssd1 vssd1 vccd1 vccd1 net3232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2719 _03631_ vssd1 vssd1 vccd1 vccd1 net3243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19846_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__clkbuf_4
X_16989_ _09171_ _09173_ vssd1 vssd1 vccd1 vccd1 _10001_ sky130_fd_sc_hd__and2_1
X_19777_ net6172 _03427_ net1690 _03424_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18728_ net3918 _06185_ _06394_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18659_ _02634_ _02652_ _02627_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire79 _06856_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_4
X_21670_ clknet_leaf_13_i_clk net854 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_mapdx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20621_ _03959_ net3966 _03960_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20552_ net3485 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6002 rbzero.tex_g1\[12\] vssd1 vssd1 vccd1 vccd1 net6526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6013 net1498 vssd1 vssd1 vccd1 vccd1 net6537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20483_ _03858_ net3520 vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__and2_1
Xhold6024 rbzero.spi_registers.buf_texadd3\[15\] vssd1 vssd1 vccd1 vccd1 net6548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6035 net1615 vssd1 vssd1 vccd1 vccd1 net6559 sky130_fd_sc_hd__dlygate4sd3_1
X_22222_ net354 net2673 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
Xhold6046 net1610 vssd1 vssd1 vccd1 vccd1 net6570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5301 _04176_ vssd1 vssd1 vccd1 vccd1 net5825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5312 net1957 vssd1 vssd1 vccd1 vccd1 net5836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6057 rbzero.tex_g1\[30\] vssd1 vssd1 vccd1 vccd1 net6581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6068 net1824 vssd1 vssd1 vccd1 vccd1 net6592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5323 rbzero.tex_b1\[61\] vssd1 vssd1 vccd1 vccd1 net5847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5334 _04235_ vssd1 vssd1 vccd1 vccd1 net5858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6079 rbzero.tex_r0\[28\] vssd1 vssd1 vccd1 vccd1 net6603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5345 _04482_ vssd1 vssd1 vccd1 vccd1 net5869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4600 net867 vssd1 vssd1 vccd1 vccd1 net5124 sky130_fd_sc_hd__dlygate4sd3_1
X_22153_ net285 net1269 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
Xhold5356 _04383_ vssd1 vssd1 vccd1 vccd1 net5880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4611 rbzero.spi_registers.texadd1\[5\] vssd1 vssd1 vccd1 vccd1 net5135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5367 _04524_ vssd1 vssd1 vccd1 vccd1 net5891 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_3_7_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_i_clk sky130_fd_sc_hd__clkbuf_8
Xhold4622 rbzero.spi_registers.texadd3\[1\] vssd1 vssd1 vccd1 vccd1 net5146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4633 rbzero.spi_registers.texadd1\[20\] vssd1 vssd1 vccd1 vccd1 net5157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5378 net2180 vssd1 vssd1 vccd1 vccd1 net5902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5389 net2563 vssd1 vssd1 vccd1 vccd1 net5913 sky130_fd_sc_hd__dlygate4sd3_1
X_21104_ _04088_ _04091_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__nand2_1
Xhold4644 net859 vssd1 vssd1 vccd1 vccd1 net5168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4655 _00833_ vssd1 vssd1 vccd1 vccd1 net5179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3910 net7825 vssd1 vssd1 vccd1 vccd1 net4434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3921 net952 vssd1 vssd1 vccd1 vccd1 net4445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4666 net898 vssd1 vssd1 vccd1 vccd1 net5190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22084_ clknet_leaf_47_i_clk net6027 vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_1
Xhold3932 _08060_ vssd1 vssd1 vccd1 vccd1 net4456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4677 net815 vssd1 vssd1 vccd1 vccd1 net5201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3943 net3240 vssd1 vssd1 vccd1 vccd1 net4467 sky130_fd_sc_hd__buf_1
Xhold4688 net1228 vssd1 vssd1 vccd1 vccd1 net5212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3954 _02540_ vssd1 vssd1 vccd1 vccd1 net4478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4699 _00861_ vssd1 vssd1 vccd1 vccd1 net5223 sky130_fd_sc_hd__dlygate4sd3_1
X_21035_ _04033_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3965 net3221 vssd1 vssd1 vccd1 vccd1 net4489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3976 net7525 vssd1 vssd1 vccd1 vccd1 net4500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3987 net3426 vssd1 vssd1 vccd1 vccd1 net4511 sky130_fd_sc_hd__buf_1
XFILLER_0_22_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3998 _00988_ vssd1 vssd1 vccd1 vccd1 net4522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21937_ clknet_leaf_7_i_clk net1221 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12670_ _05826_ _05831_ net7 vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__mux2_1
X_21868_ clknet_leaf_100_i_clk net1238 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _04637_ _04605_ _04606_ _04740_ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a41o_1
XFILLER_0_182_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21799_ clknet_leaf_12_i_clk net1037 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ _07479_ _07472_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ net3869 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14271_ net569 _07410_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nand2_1
X_11483_ rbzero.spi_registers.texadd3\[8\] rbzero.spi_registers.texadd1\[8\] rbzero.spi_registers.texadd0\[8\]
+ rbzero.spi_registers.texadd2\[8\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ _08559_ _08493_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__or2_1
Xhold7270 rbzero.wall_tracer.stepDistX\[-7\] vssd1 vssd1 vccd1 vccd1 net7794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7281 _02350_ vssd1 vssd1 vccd1 vccd1 net7805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13222_ net3984 net3804 _06371_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7292 rbzero.wall_tracer.stepDistY\[-6\] vssd1 vssd1 vccd1 vccd1 net7816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6580 rbzero.tex_g1\[9\] vssd1 vssd1 vccd1 vccd1 net7104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6591 net2292 vssd1 vssd1 vccd1 vccd1 net7115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13153_ net3417 vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12104_ _05271_ _05272_ _05235_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__mux2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5890 rbzero.tex_g1\[18\] vssd1 vssd1 vccd1 vccd1 net6414 sky130_fd_sc_hd__dlygate4sd3_1
X_17961_ _02001_ _02009_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__xnor2_1
X_13084_ net3921 rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__or2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16912_ _09933_ vssd1 vssd1 vccd1 vccd1 _09941_ sky130_fd_sc_hd__clkbuf_4
X_12035_ reg_rgb\[6\] _05203_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__mux2_4
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19700_ _02491_ _02514_ net3076 vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__and3_2
X_17892_ _01825_ _01941_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__xnor2_1
X_16843_ _09778_ _09911_ _08296_ vssd1 vssd1 vccd1 vccd1 _09913_ sky130_fd_sc_hd__o21ai_1
X_19631_ net4607 net798 _03352_ _03343_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ net1727 _03305_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__or2_1
X_16774_ _09702_ _09704_ _09701_ vssd1 vssd1 vccd1 vccd1 _09844_ sky130_fd_sc_hd__a21boi_2
X_13986_ net536 _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18513_ net4446 net4806 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15725_ _08796_ _08798_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__and2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _06093_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_1
X_19493_ _02998_ _03265_ net1736 _03260_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _02468_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__nand2_1
X_15656_ _08394_ _08411_ _08470_ _08484_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__or4_1
XFILLER_0_185_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12868_ net6265 _06012_ _06008_ net3964 vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _07755_ _07757_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nand2_1
X_11819_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__buf_4
X_18375_ _10010_ net3396 _02409_ _10080_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__o31ai_1
X_15587_ _08327_ net4954 _08540_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__or3b_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12799_ _05955_ net22 vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__nor2_2
X_20336__69 clknet_1_1__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
X_17326_ _09904_ _10201_ vssd1 vssd1 vccd1 vccd1 _10327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14538_ _07643_ _07684_ _07688_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _08315_ _08331_ _08641_ _08548_ vssd1 vssd1 vccd1 vccd1 _10258_ sky130_fd_sc_hd__or4_2
Xclkbuf_0__03995_ _03995_ vssd1 vssd1 vccd1 vccd1 clknet_0__03995_ sky130_fd_sc_hd__clkbuf_16
X_14469_ _07618_ _07509_ _07619_ _07536_ _06611_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__o221a_2
X_16208_ _09281_ _09282_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17188_ _09850_ _09892_ _09891_ vssd1 vssd1 vccd1 vccd1 _10190_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _09208_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3206 _03838_ vssd1 vssd1 vccd1 vccd1 net3730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3217 net7524 vssd1 vssd1 vccd1 vccd1 net3741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3228 net1355 vssd1 vssd1 vccd1 vccd1 net3752 sky130_fd_sc_hd__buf_1
XFILLER_0_110_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3239 _00476_ vssd1 vssd1 vccd1 vccd1 net3763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2505 net7447 vssd1 vssd1 vccd1 vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2516 net4343 vssd1 vssd1 vccd1 vccd1 net3040 sky130_fd_sc_hd__clkbuf_2
Xhold2527 _00635_ vssd1 vssd1 vccd1 vccd1 net3051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2538 _02484_ vssd1 vssd1 vccd1 vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1804 net6785 vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2549 _00645_ vssd1 vssd1 vccd1 vccd1 net3073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 _01521_ vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1826 _04453_ vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_19829_ net625 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
Xhold1837 _04431_ vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1848 _01112_ vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 net7090 vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21722_ clknet_leaf_8_i_clk net2595 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21653_ clknet_leaf_16_i_clk net5564 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_otherx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20604_ _04881_ _05816_ _03033_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or3b_1
XFILLER_0_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21584_ clknet_leaf_21_i_clk net5726 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20949__359 clknet_1_1__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__inv_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20535_ net3362 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20466_ net3709 net1274 _03845_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5120 net1346 vssd1 vssd1 vccd1 vccd1 net5644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5131 rbzero.floor_leak\[3\] vssd1 vssd1 vccd1 vccd1 net5655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22205_ net337 net2267 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
Xhold5142 _01090_ vssd1 vssd1 vccd1 vccd1 net5666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5153 rbzero.mapdyw\[1\] vssd1 vssd1 vccd1 vccd1 net5677 sky130_fd_sc_hd__dlygate4sd3_1
X_20397_ _03791_ net3685 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5164 _01071_ vssd1 vssd1 vccd1 vccd1 net5688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4430 _08661_ vssd1 vssd1 vccd1 vccd1 net4954 sky130_fd_sc_hd__clkbuf_4
Xhold5175 net3619 vssd1 vssd1 vccd1 vccd1 net5699 sky130_fd_sc_hd__dlygate4sd3_1
X_22136_ net268 net1758 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5186 net1524 vssd1 vssd1 vccd1 vccd1 net5710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4441 net664 vssd1 vssd1 vccd1 vccd1 net4965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4452 _01590_ vssd1 vssd1 vccd1 vccd1 net4976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5197 net1529 vssd1 vssd1 vccd1 vccd1 net5721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4463 net717 vssd1 vssd1 vccd1 vccd1 net4987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4474 rbzero.spi_registers.texadd3\[10\] vssd1 vssd1 vccd1 vccd1 net4998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4485 net764 vssd1 vssd1 vccd1 vccd1 net5009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3740 net7845 vssd1 vssd1 vccd1 vccd1 net4264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4496 net856 vssd1 vssd1 vccd1 vccd1 net5020 sky130_fd_sc_hd__dlygate4sd3_1
X_22067_ clknet_leaf_8_i_clk net3261 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3751 net1603 vssd1 vssd1 vccd1 vccd1 net4275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3762 _00512_ vssd1 vssd1 vccd1 vccd1 net4286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03984_ clknet_0__03984_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03984_
+ sky130_fd_sc_hd__clkbuf_16
X_21018_ _04018_ _04021_ _04022_ _04017_ net4975 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a32o_1
Xhold3784 net1158 vssd1 vssd1 vccd1 vccd1 net4308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3795 _00648_ vssd1 vssd1 vccd1 vccd1 net4319 sky130_fd_sc_hd__dlygate4sd3_1
X_13840_ _06931_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20694__129 clknet_1_0__leaf__03983_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__inv_2
XFILLER_0_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _06916_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__buf_6
X_10983_ net6648 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15510_ _08560_ _08574_ _08582_ _08584_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_168_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ net13 net12 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__and2b_1
X_16490_ _08372_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__clkbuf_4
X_15441_ _08484_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__clkbuf_4
X_12653_ _05806_ _05814_ net8 vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__o21ba_1
X_18160_ _02093_ _02107_ _02206_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a21bo_1
X_11604_ net6025 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__clkbuf_4
X_15372_ _08397_ _08446_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12584_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _04989_ vssd1 vssd1 vccd1 vccd1 _05749_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17111_ _10110_ _10111_ vssd1 vssd1 vccd1 vccd1 _10113_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14323_ net534 vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18091_ _02137_ _02138_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__nor2_1
X_11535_ _04692_ rbzero.spi_registers.texadd3\[23\] vssd1 vssd1 vccd1 vccd1 _04707_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17042_ _10048_ net4560 net4903 vssd1 vssd1 vccd1 vccd1 _10049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03780_ _03780_ vssd1 vssd1 vccd1 vccd1 clknet_0__03780_ sky130_fd_sc_hd__clkbuf_16
X_14254_ _07351_ _07398_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__nor2_8
X_11466_ net7317 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13205_ net3984 _06183_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11397_ net2810 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
X_14185_ _07324_ _07335_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _06287_ net3426 net3542 _06285_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__a22o_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _02523_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__clkbuf_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17944_ _01991_ _01992_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__xnor2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ net4345 _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__xnor2_1
X_12018_ _05119_ _05121_ net4077 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__mux2_1
X_17875_ _01923_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19614_ net3038 _03340_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or2_1
X_16826_ _09716_ _09755_ _09754_ vssd1 vssd1 vccd1 vccd1 _09896_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757_ _09711_ _09714_ _09825_ vssd1 vssd1 vccd1 vccd1 _09827_ sky130_fd_sc_hd__nand3_1
XFILLER_0_159_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19545_ _03302_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__clkbuf_4
X_13969_ _07096_ _07097_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15708_ _08710_ _08782_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__xnor2_2
X_16688_ _09757_ _09758_ vssd1 vssd1 vccd1 vccd1 _09759_ sky130_fd_sc_hd__nor2_1
X_19476_ _02492_ _03238_ net3076 net6524 vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ _08712_ _08713_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__and2_1
X_18427_ _02445_ _02448_ _02446_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _02390_ _02393_ _01870_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ _10279_ _10309_ vssd1 vssd1 vccd1 vccd1 _10310_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18289_ net4475 net4315 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold901 net6490 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 net6540 vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _01392_ vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
X_20251_ net3646 _03744_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold934 net7088 vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold945 _00628_ vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 net6472 vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 net5438 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__buf_1
Xhold978 net6482 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20182_ net5481 _03705_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__or2_1
Xhold3003 _01246_ vssd1 vssd1 vccd1 vccd1 net3527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 net6552 vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3025 _03842_ vssd1 vssd1 vccd1 vccd1 net3549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3036 _01202_ vssd1 vssd1 vccd1 vccd1 net3560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3047 _01232_ vssd1 vssd1 vccd1 vccd1 net3571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2302 net5951 vssd1 vssd1 vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3058 _03893_ vssd1 vssd1 vccd1 vccd1 net3582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2313 _03536_ vssd1 vssd1 vccd1 vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 net7291 vssd1 vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3069 _01177_ vssd1 vssd1 vccd1 vccd1 net3593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2335 _04517_ vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1601 net6889 vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2346 net7301 vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1612 _01410_ vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2357 net7297 vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1623 _04538_ vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2368 net3359 vssd1 vssd1 vccd1 vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2379 _04285_ vssd1 vssd1 vccd1 vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 net4678 vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__buf_1
XFILLER_0_208_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1645 net7202 vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1656 net5901 vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1667 net5934 vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1678 _01313_ vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1689 net6885 vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21705_ clknet_leaf_20_i_clk net5036 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21636_ clknet_leaf_28_i_clk net1533 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21567_ clknet_leaf_26_i_clk net5028 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11320_ net7123 net6976 _04540_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20518_ net2990 net3275 _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21498_ clknet_leaf_13_i_clk net2896 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11251_ net6375 net6696 _04503_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__mux2_1
X_20449_ net3549 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ net6972 net7042 _04470_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4260 _08226_ vssd1 vssd1 vccd1 vccd1 net4784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4271 _03653_ vssd1 vssd1 vccd1 vccd1 net4795 sky130_fd_sc_hd__dlygate4sd3_1
X_22119_ net251 net1437 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15990_ _08449_ _08501_ _08514_ _09064_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__o22a_1
Xhold4282 net913 vssd1 vssd1 vccd1 vccd1 net4806 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold4293 _02907_ vssd1 vssd1 vccd1 vccd1 net4817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3570 _04908_ vssd1 vssd1 vccd1 vccd1 net4094 sky130_fd_sc_hd__dlygate4sd3_1
X_14941_ _08087_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__clkbuf_1
Xhold3581 net4218 vssd1 vssd1 vccd1 vccd1 net4105 sky130_fd_sc_hd__clkbuf_2
Xhold3592 _00866_ vssd1 vssd1 vccd1 vccd1 net4116 sky130_fd_sc_hd__dlygate4sd3_1
X_17660_ _09593_ _01711_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__nor2_1
Xhold2880 net4948 vssd1 vssd1 vccd1 vccd1 net3404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2891 _01210_ vssd1 vssd1 vccd1 vccd1 net3415 sky130_fd_sc_hd__dlygate4sd3_1
X_14872_ net7891 _08016_ _08022_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__a21oi_1
X_16611_ _09680_ _09681_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13823_ _06895_ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__nor2_1
X_17591_ _09805_ _09447_ vssd1 vssd1 vccd1 vccd1 _10589_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16542_ _09371_ _09490_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__nor2_1
X_19330_ net1712 _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or2_1
X_13754_ _06869_ _06893_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__or2_4
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10966_ net1822 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19261_ net5395 _03132_ _03134_ _03128_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__o211a_1
X_12705_ net4021 _05844_ _05852_ _05299_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a22o_1
X_16473_ _09091_ _08795_ vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__nor2_1
X_13685_ _06830_ _06832_ _06835_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__and3_1
X_10897_ net2496 net7304 _04321_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18212_ _02073_ _02076_ _02074_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15424_ _08493_ _08498_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19192_ net1790 _03079_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__or2_1
X_12636_ net57 _05795_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ _01684_ _10520_ _01711_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ _08428_ _08429_ _08305_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__a21o_2
X_12567_ _05003_ _05731_ _05009_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14306_ _07454_ _07456_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18074_ _02120_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11518_ rbzero.spi_registers.texadd3\[16\] rbzero.spi_registers.texadd1\[16\] rbzero.spi_registers.texadd0\[16\]
+ rbzero.spi_registers.texadd2\[16\] _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04690_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15286_ net5463 vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__inv_2
X_12498_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _05219_ vssd1 vssd1 vccd1 vccd1 _05664_
+ sky130_fd_sc_hd__mux2_1
Xhold208 net4636 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ net4556 net4719 vssd1 vssd1 vccd1 vccd1 _10033_ sky130_fd_sc_hd__nor2_1
Xhold219 net5012 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ _07386_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__nand2_1
X_11449_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ _07313_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _06269_ net4577 net3780 _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__o22a_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _07189_ _07230_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__and2_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _02953_ net3984 _01749_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__mux2_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17858_ _01906_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16809_ _09875_ _09876_ _09878_ vssd1 vssd1 vccd1 vccd1 _09879_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17789_ _01709_ _01717_ _01715_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19528_ net5428 _03288_ _03291_ _03280_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19459_ net3104 net2995 _03241_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22470_ clknet_leaf_79_i_clk net4793 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21421_ clknet_leaf_85_i_clk net3196 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21352_ clknet_leaf_35_i_clk net3380 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21283_ clknet_leaf_63_i_clk _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold720 net5508 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold731 net5604 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 net5589 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold753 net5583 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
X_20234_ _03675_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__clkbuf_4
Xhold764 net5516 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 net4448 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 net5608 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 net5650 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
X_20165_ _03675_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__clkbuf_4
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2110 _01446_ vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2121 net7164 vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2132 net7210 vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2143 _01348_ vssd1 vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_20096_ net3562 net2938 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__and2_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2154 net5909 vssd1 vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 net7192 vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 net6665 vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2176 _04229_ vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1431 _01519_ vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1442 _00931_ vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2187 net7124 vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2198 _01457_ vssd1 vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 net7080 vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1464 rbzero.spi_registers.buf_texadd3\[12\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1475 net7631 vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 net7057 vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _03418_ vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10820_ net2061 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10751_ net2338 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13470_ _06428_ _06620_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ net1180 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _05177_ _05585_ _05587_ _05244_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__o211a_1
X_21619_ clknet_leaf_18_i_clk net5001 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15140_ _04621_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__buf_4
X_12352_ _05518_ _05519_ _04991_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ net7038 net2613 _04529_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15071_ net3539 _06386_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__nand2_1
X_12283_ net3378 _05448_ _05450_ _05115_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_121_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ _07158_ _07160_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__xnor2_1
X_11234_ net5900 net5962 _04492_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__mux2_1
X_18830_ _02811_ _02812_ _02813_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a21bo_1
X_11165_ net2578 net7119 _04459_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4090 rbzero.pov.ready_buffer\[0\] vssd1 vssd1 vccd1 vccd1 net4614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15973_ _08456_ _08626_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__nor2_1
X_11096_ net7032 net6666 _04426_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
X_18761_ net4640 net4905 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17712_ _10596_ _01666_ _01664_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a21o_1
X_14924_ net7458 _08071_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__nor2_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ _02680_ _02681_ _02683_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__and3_1
Xhold80 _03127_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__04000_ clknet_0__04000_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04000_
+ sky130_fd_sc_hd__clkbuf_16
Xhold91 net4259 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _01673_ _01674_ _01694_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a21o_1
X_14855_ _07995_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__buf_2
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ _06933_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__clkbuf_4
X_17574_ _10572_ net4501 net4903 vssd1 vssd1 vccd1 vccd1 _10573_ sky130_fd_sc_hd__mux2_1
X_14786_ _07232_ _07524_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__or2_1
XFILLER_0_203_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ _05160_ net4009 _04604_ _05161_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__o221a_1
X_16525_ _09086_ _09595_ _09596_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__or3_1
X_19313_ net2593 _03160_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__or2_1
X_13737_ _06781_ _06796_ _06806_ net563 vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__a211o_2
X_10949_ net5899 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16456_ net4313 _08296_ _09527_ _09528_ _08239_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19244_ net5353 _03119_ _03124_ _03115_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13668_ _06733_ _06812_ _06815_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _08481_ _04846_ _08381_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__mux2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19175_ net5996 _03078_ net1635 _03074_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__o211a_1
X_12619_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__inv_2
X_16387_ _09458_ _09459_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__nor2_1
X_13599_ _06743_ _06746_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__or3_1
Xhold6409 rbzero.tex_b0\[28\] vssd1 vssd1 vccd1 vccd1 net6933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_171_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _02173_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ net4294 _08375_ net3003 vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5708 rbzero.spi_registers.buf_texadd3\[5\] vssd1 vssd1 vccd1 vccd1 net6232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5719 net2920 vssd1 vssd1 vccd1 vccd1 net6243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18057_ _01812_ _10407_ _02043_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15269_ _08341_ _08342_ _08343_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__or3_1
X_17008_ _10014_ _10017_ vssd1 vssd1 vccd1 vccd1 _10018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20999__25 clknet_1_1__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_0_10_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18959_ _02864_ net3018 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__xor2_1
XFILLER_0_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21970_ net195 net1419 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer12 net3203 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_2
Xrebuffer23 net546 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_1
Xrebuffer34 _07058_ vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer45 net568 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer56 net581 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer67 _06624_ vssd1 vssd1 vccd1 vccd1 net3237 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22453_ clknet_leaf_51_i_clk _01622_ vssd1 vssd1 vccd1 vccd1 reg_vsync sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6910 net7912 vssd1 vssd1 vccd1 vccd1 net7434 sky130_fd_sc_hd__clkbuf_2
X_21404_ clknet_leaf_44_i_clk net1213 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6921 rbzero.debug_overlay.playerY\[-2\] vssd1 vssd1 vccd1 vccd1 net7445 sky130_fd_sc_hd__dlygate4sd3_1
X_22384_ net516 net2637 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6943 rbzero.wall_tracer.stepDistY\[-3\] vssd1 vssd1 vccd1 vccd1 net7467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6954 _06721_ vssd1 vssd1 vccd1 vccd1 net7478 sky130_fd_sc_hd__buf_1
Xhold6965 net4371 vssd1 vssd1 vccd1 vccd1 net7489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21335_ clknet_leaf_50_i_clk net5473 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6976 net4165 vssd1 vssd1 vccd1 vccd1 net7500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6987 _08349_ vssd1 vssd1 vccd1 vccd1 net7511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6998 rbzero.wall_tracer.trackDistX\[-10\] vssd1 vssd1 vccd1 vccd1 net7522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold550 net6392 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
X_21266_ clknet_leaf_58_i_clk _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold561 net4192 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 net5486 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 net6364 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
X_20217_ net1318 _03731_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21197_ _02751_ _02757_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__or2b_1
Xhold594 net5522 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20148_ net5554 _03692_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20079_ net3702 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__clkbuf_1
X_12970_ net3857 net3135 vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nand2_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 net6759 vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1261 _03416_ vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ _05087_ _05090_ _05009_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__mux2_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 _01337_ vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _03406_ vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1294 net6827 vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _07696_ _07739_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__xor2_2
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__buf_4
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ net2308 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__clkbuf_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _07083_ _07618_ _07464_ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _04945_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__nor2_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20814__237 clknet_1_1__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__inv_2
X_16310_ _09234_ _09236_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13522_ _06579_ _06581_ _06672_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and3b_1
X_10734_ net5859 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__clkbuf_1
X_17290_ _10281_ _10289_ vssd1 vssd1 vccd1 vccd1 _10291_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _09188_ _09303_ _09314_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ _06511_ _06513_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__nand2_2
X_10665_ net5813 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ _05569_ _05570_ _05235_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__mux2_1
X_16172_ _09245_ _09246_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _06532_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ _08218_ _08233_ net3628 _08215_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__o211a_1
X_12335_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _05493_ vssd1 vssd1 vccd1 vccd1 _05503_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19931_ net2914 _03477_ _03532_ _03548_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a211o_1
X_15054_ _08185_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
X_12266_ net3008 _05373_ _05381_ net4218 vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14005_ _07119_ _07147_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11217_ net6493 net6776 _04481_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__mux2_1
X_20708__142 clknet_1_0__leaf__03984_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__inv_2
XFILLER_0_43_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19862_ net4300 _03475_ net2946 _03496_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__o211a_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__clkbuf_4
X_12197_ _05343_ _05357_ _05364_ _05365_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20860__279 clknet_1_0__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__inv_2
X_18813_ _05396_ _02803_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__nand2_1
X_11148_ net750 net5920 _04448_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__mux2_1
X_19793_ net3070 _03442_ net2156 _03441_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18744_ net3895 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__clkbuf_1
X_15956_ _09013_ _09029_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__nor2_1
X_11079_ net5985 net5834 _04415_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14907_ _08006_ _08014_ _08055_ _06663_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__o211a_1
X_15887_ _08961_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__clkbuf_4
X_18675_ _02680_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nand2_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17626_ _01676_ _01677_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ _07986_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__xor2_2
XFILLER_0_188_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17557_ _10553_ _10554_ vssd1 vssd1 vccd1 vccd1 _10556_ sky130_fd_sc_hd__and2_1
X_14769_ _07532_ _07805_ _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16508_ _09561_ _09579_ vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__xnor2_2
X_20754__184 clknet_1_1__leaf__03988_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__inv_2
X_17488_ _10383_ _08795_ vssd1 vssd1 vccd1 vccd1 _10487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19227_ _02992_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__clkbuf_4
X_16439_ _09510_ _09511_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6206 net2274 vssd1 vssd1 vccd1 vccd1 net6730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6217 rbzero.tex_b0\[51\] vssd1 vssd1 vccd1 vccd1 net6741 sky130_fd_sc_hd__dlygate4sd3_1
X_19158_ net5442 _03065_ _03072_ _03061_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__o211a_1
Xhold6228 net2017 vssd1 vssd1 vccd1 vccd1 net6752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6239 rbzero.tex_b1\[54\] vssd1 vssd1 vccd1 vccd1 net6763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5505 net3072 vssd1 vssd1 vccd1 vccd1 net6029 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5516 gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 net6040 sky130_fd_sc_hd__dlygate4sd3_1
X_18109_ _02082_ _02156_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ net2123 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
Xhold5527 net2282 vssd1 vssd1 vccd1 vccd1 net6051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5538 net1712 vssd1 vssd1 vccd1 vccd1 net6062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4804 net1028 vssd1 vssd1 vccd1 vccd1 net5328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5549 _00899_ vssd1 vssd1 vccd1 vccd1 net6073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21120_ _04103_ _04104_ _04105_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o21ba_1
Xhold4815 _00782_ vssd1 vssd1 vccd1 vccd1 net5339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4826 net606 vssd1 vssd1 vccd1 vccd1 net5350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4837 _00835_ vssd1 vssd1 vccd1 vccd1 net5361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4848 _00844_ vssd1 vssd1 vccd1 vccd1 net5372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4859 net1284 vssd1 vssd1 vccd1 vccd1 net5383 sky130_fd_sc_hd__dlygate4sd3_1
X_21051_ net4152 net4763 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20002_ net3902 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21953_ net178 net2736 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21884_ clknet_leaf_98_i_clk net1277 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ clknet_1_1__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__buf_1
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22436_ clknet_leaf_38_i_clk net4651 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6740 net2793 vssd1 vssd1 vccd1 vccd1 net7264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7485 rbzero.debug_overlay.playerX\[-7\] vssd1 vssd1 vccd1 vccd1 net8009 sky130_fd_sc_hd__dlygate4sd3_1
X_22367_ net499 net2087 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold6751 rbzero.tex_b0\[12\] vssd1 vssd1 vccd1 vccd1 net7275 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__04003_ clknet_0__04003_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04003_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6762 net2876 vssd1 vssd1 vccd1 vccd1 net7286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6773 rbzero.tex_b1\[12\] vssd1 vssd1 vccd1 vccd1 net7297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6784 rbzero.tex_r0\[27\] vssd1 vssd1 vccd1 vccd1 net7308 sky130_fd_sc_hd__dlygate4sd3_1
X_12120_ _04992_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or2_1
Xhold6795 _09945_ vssd1 vssd1 vccd1 vccd1 net7319 sky130_fd_sc_hd__dlygate4sd3_1
X_21318_ clknet_leaf_72_i_clk net2994 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_22298_ net430 net2109 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12051_ rbzero.tex_r1\[51\] rbzero.tex_r1\[50\] _05219_ vssd1 vssd1 vccd1 vccd1 _05220_
+ sky130_fd_sc_hd__mux2_1
Xhold380 net5321 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21249_ clknet_leaf_50_i_clk net3358 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold391 net5329 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net6345 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__clkbuf_1
X_15810_ _08871_ _08883_ _08884_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__a21oi_2
X_16790_ _09852_ _09859_ vssd1 vssd1 vccd1 vccd1 _09860_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15741_ _08810_ _08811_ _08812_ _08815_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__a22o_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nand2_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 net6257 vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 net6558 vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _05069_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or2_1
X_15672_ _08695_ _08680_ _08694_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__and3_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ net4332 net3061 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__nor2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ net33 _06034_ _06041_ _05996_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__a22o_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _09582_ _09484_ vssd1 vssd1 vccd1 vccd1 _10411_ sky130_fd_sc_hd__nor2_1
X_14623_ _06918_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__buf_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _04989_ vssd1 vssd1 vccd1 vccd1 _05005_
+ sky130_fd_sc_hd__mux2_1
X_18391_ _02423_ net4536 _02411_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _10340_ _10341_ vssd1 vssd1 vccd1 vccd1 _10342_ sky130_fd_sc_hd__nor2_2
XFILLER_0_157_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _07474_ _07589_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nor2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__03980_ clknet_0__03980_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03980_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11766_ net1583 _04934_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13505_ _06628_ _06651_ _06655_ _06648_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__or4b_2
X_17273_ _10272_ _10273_ vssd1 vssd1 vccd1 vccd1 _10274_ sky130_fd_sc_hd__and2b_1
X_10717_ net5927 net1683 _04225_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14485_ _07634_ _07635_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11697_ net4971 net2536 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ _09292_ _09293_ net7407 _08633_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__a31o_1
X_19012_ net3887 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
X_13436_ _06579_ _06581_ _06584_ _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__and4b_2
X_10648_ net2380 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer3 _07963_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ _09223_ _09229_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__xnor2_2
X_13367_ _06478_ net82 _06485_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15106_ _08200_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__clkbuf_2
X_12318_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _05262_ vssd1 vssd1 vccd1 vccd1 _05486_
+ sky130_fd_sc_hd__mux2_1
X_16086_ _09138_ _08874_ _09158_ vssd1 vssd1 vccd1 vccd1 _09161_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19914_ net2837 _03537_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__nor2_1
X_15037_ net7431 _06714_ _08123_ _08171_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ rbzero.debug_overlay.facingX\[10\] _05371_ _05417_ vssd1 vssd1 vccd1 vccd1
+ _05418_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2709 net4537 vssd1 vssd1 vccd1 vccd1 net3233 sky130_fd_sc_hd__buf_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19845_ _03038_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__nor2_4
X_19776_ net1689 _03429_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__or2_1
X_16988_ _09171_ _09173_ vssd1 vssd1 vccd1 vccd1 _10000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18727_ net3917 _06227_ _02261_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
X_15939_ _09004_ _09005_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__xor2_1
XFILLER_0_211_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18658_ _02663_ net4767 _02662_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ _01659_ _01660_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18589_ net4666 rbzero.wall_tracer.rayAddendX\[1\] vssd1 vssd1 vccd1 vccd1 _02601_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20620_ _05825_ net3965 net3979 _04597_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a31o_1
XFILLER_0_188_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20551_ _03902_ net3484 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6003 net1515 vssd1 vssd1 vccd1 vccd1 net6527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6014 rbzero.tex_b1\[22\] vssd1 vssd1 vccd1 vccd1 net6538 sky130_fd_sc_hd__dlygate4sd3_1
X_20482_ net3519 net1341 _03845_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6025 net1543 vssd1 vssd1 vccd1 vccd1 net6549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22221_ net353 net2133 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold6036 _03256_ vssd1 vssd1 vccd1 vccd1 net6560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6047 _04454_ vssd1 vssd1 vccd1 vccd1 net6571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5302 net2428 vssd1 vssd1 vccd1 vccd1 net5826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6058 net1680 vssd1 vssd1 vccd1 vccd1 net6582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5313 rbzero.spi_registers.spi_buffer\[10\] vssd1 vssd1 vccd1 vccd1 net5837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6069 rbzero.tex_b1\[55\] vssd1 vssd1 vccd1 vccd1 net6593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5324 net1832 vssd1 vssd1 vccd1 vccd1 net5848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5335 net1459 vssd1 vssd1 vccd1 vccd1 net5859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4601 _00827_ vssd1 vssd1 vccd1 vccd1 net5125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5346 net1857 vssd1 vssd1 vccd1 vccd1 net5870 sky130_fd_sc_hd__dlygate4sd3_1
X_22152_ net284 net1487 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5357 net2098 vssd1 vssd1 vccd1 vccd1 net5881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4612 net925 vssd1 vssd1 vccd1 vccd1 net5136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5368 net1875 vssd1 vssd1 vccd1 vccd1 net5892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4623 net896 vssd1 vssd1 vccd1 vccd1 net5147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5379 rbzero.tex_b1\[43\] vssd1 vssd1 vccd1 vccd1 net5903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4634 net892 vssd1 vssd1 vccd1 vccd1 net5158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21103_ net4186 net4469 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nand2_1
Xhold3900 rbzero.debug_overlay.vplaneX\[-9\] vssd1 vssd1 vccd1 vccd1 net4424 sky130_fd_sc_hd__buf_2
Xhold4645 _01593_ vssd1 vssd1 vccd1 vccd1 net5169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4656 net871 vssd1 vssd1 vccd1 vccd1 net5180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3911 net3193 vssd1 vssd1 vccd1 vccd1 net4435 sky130_fd_sc_hd__buf_1
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22083_ clknet_leaf_49_i_clk net1452 vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync
+ sky130_fd_sc_hd__dfxtp_1
Xhold3922 rbzero.debug_overlay.vplaneX\[-7\] vssd1 vssd1 vccd1 vccd1 net4446 sky130_fd_sc_hd__buf_2
Xhold4667 _00838_ vssd1 vssd1 vccd1 vccd1 net5191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3933 net7542 vssd1 vssd1 vccd1 vccd1 net4457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4678 _00860_ vssd1 vssd1 vccd1 vccd1 net5202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3944 rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 net4468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4689 _01079_ vssd1 vssd1 vccd1 vccd1 net5213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3955 _02544_ vssd1 vssd1 vccd1 vccd1 net4479 sky130_fd_sc_hd__dlygate4sd3_1
X_21034_ _04034_ _04035_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3966 net7543 vssd1 vssd1 vccd1 vccd1 net4490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3977 net3432 vssd1 vssd1 vccd1 vccd1 net4501 sky130_fd_sc_hd__buf_1
Xhold3988 net7527 vssd1 vssd1 vccd1 vccd1 net4512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3999 net722 vssd1 vssd1 vccd1 vccd1 net4523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21936_ clknet_leaf_9_i_clk net1412 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21867_ clknet_leaf_100_i_clk net955 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _04761_ _04789_ _04791_ _04613_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a31o_1
XFILLER_0_182_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21798_ clknet_leaf_11_i_clk net727 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _04699_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14270_ _07419_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__xnor2_1
X_11482_ rbzero.texu_hot\[3\] _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13221_ _06372_ _06376_ _06222_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__a21oi_1
Xhold7271 net4369 vssd1 vssd1 vccd1 vccd1 net7795 sky130_fd_sc_hd__dlygate4sd3_1
X_22419_ clknet_leaf_66_i_clk net1082 vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold7282 rbzero.wall_tracer.stepDistY\[0\] vssd1 vssd1 vccd1 vccd1 net7806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7293 net4373 vssd1 vssd1 vccd1 vccd1 net7817 sky130_fd_sc_hd__dlygate4sd3_1
X_20926__338 clknet_1_0__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__inv_2
XFILLER_0_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6570 rbzero.tex_g0\[44\] vssd1 vssd1 vccd1 vccd1 net7094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ net3047 vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__inv_2
Xhold6581 net2478 vssd1 vssd1 vccd1 vccd1 net7105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6592 _04306_ vssd1 vssd1 vccd1 vccd1 net7116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ rbzero.tex_r1\[7\] rbzero.tex_r1\[6\] _05072_ vssd1 vssd1 vccd1 vccd1 _05272_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5880 _04289_ vssd1 vssd1 vccd1 vccd1 net6404 sky130_fd_sc_hd__dlygate4sd3_1
X_17960_ _02007_ _02008_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__nor2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ net3921 net6216 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__nand2_1
Xhold5891 net1201 vssd1 vssd1 vccd1 vccd1 net6415 sky130_fd_sc_hd__dlygate4sd3_1
X_16911_ net4179 _09939_ _09940_ net7552 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
X_12034_ net45 vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__clkbuf_8
X_17891_ _01937_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19630_ net4322 _03326_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__or2_1
XFILLER_0_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16842_ _09778_ _09911_ vssd1 vssd1 vccd1 vccd1 _09912_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19561_ net5065 _03303_ _03312_ _03295_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__o211a_1
X_16773_ _09839_ _09842_ vssd1 vssd1 vccd1 vccd1 _09843_ sky130_fd_sc_hd__xor2_1
X_13985_ _07115_ _07116_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ net4493 net4791 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15724_ _08796_ _08798_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__nor2_1
X_12936_ reg_gpout\[5\] clknet_1_1__leaf__06092_ net45 vssd1 vssd1 vccd1 vccd1 _06093_
+ sky130_fd_sc_hd__mux2_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ net6290 _03266_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__or2_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18443_ net4437 net4380 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__nand2_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _08728_ _08729_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ net31 net32 _06021_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a32o_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20671__108 clknet_1_1__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__inv_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11818_ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__buf_4
X_14606_ _07754_ _07756_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__xnor2_1
X_15586_ rbzero.wall_tracer.visualWallDist\[-10\] _08298_ vssd1 vssd1 vccd1 vccd1
+ _08661_ sky130_fd_sc_hd__nand2_1
X_18374_ _02407_ net3234 net3395 _02399_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__and2_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _10324_ _10325_ vssd1 vssd1 vccd1 vccd1 _10326_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14537_ _07685_ _07687_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__or2b_1
X_11749_ net785 net2467 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03994_ _03994_ vssd1 vssd1 vccd1 vccd1 clknet_0__03994_ sky130_fd_sc_hd__clkbuf_16
X_17256_ _08556_ vssd1 vssd1 vccd1 vccd1 _10257_ sky130_fd_sc_hd__buf_2
X_14468_ _07533_ _07535_ _07465_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13419_ _06472_ _06477_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__nand2_1
X_16207_ net4893 net5463 net4088 vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__mux2_2
X_17187_ _10149_ _10188_ vssd1 vssd1 vccd1 vccd1 _10189_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14399_ _07549_ _07545_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _09211_ _09212_ vssd1 vssd1 vccd1 vccd1 _09213_ sky130_fd_sc_hd__xnor2_2
X_20866__285 clknet_1_1__leaf__03999_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__inv_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _09137_ _09142_ _09143_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__a21oi_1
Xhold3207 _01199_ vssd1 vssd1 vccd1 vccd1 net3731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3218 net3058 vssd1 vssd1 vccd1 vccd1 net3742 sky130_fd_sc_hd__buf_1
Xhold3229 _03927_ vssd1 vssd1 vccd1 vccd1 net3753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2506 rbzero.pov.ready_buffer\[62\] vssd1 vssd1 vccd1 vccd1 net3030 sky130_fd_sc_hd__buf_1
Xhold2517 net7823 vssd1 vssd1 vccd1 vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2528 net6197 vssd1 vssd1 vccd1 vccd1 net3052 sky130_fd_sc_hd__buf_1
XFILLER_0_209_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2539 net5683 vssd1 vssd1 vccd1 vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 net6787 vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1816 net6861 vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
X_19828_ net6322 _03026_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__and2_1
Xhold1827 _01334_ vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1838 _01354_ vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 net6941 vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
X_19759_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__buf_2
XFILLER_0_155_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21721_ clknet_leaf_8_i_clk net1694 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21652_ clknet_leaf_16_i_clk net5369 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_otherx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20603_ net1108 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21583_ clknet_leaf_21_i_clk net5716 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20534_ _03880_ net3361 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20465_ net3766 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5110 _00758_ vssd1 vssd1 vccd1 vccd1 net5634 sky130_fd_sc_hd__dlygate4sd3_1
X_22204_ net336 net2220 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
Xhold5121 rbzero.pov.spi_buffer\[38\] vssd1 vssd1 vccd1 vccd1 net5645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5132 net1326 vssd1 vssd1 vccd1 vccd1 net5656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5143 rbzero.pov.spi_buffer\[39\] vssd1 vssd1 vccd1 vccd1 net5667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5154 net1312 vssd1 vssd1 vccd1 vccd1 net5678 sky130_fd_sc_hd__dlygate4sd3_1
X_20396_ net2900 net3684 _03801_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__mux2_1
Xhold4420 gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5165 rbzero.spi_registers.texadd3\[8\] vssd1 vssd1 vccd1 vccd1 net5689 sky130_fd_sc_hd__dlygate4sd3_1
X_22135_ net267 net2598 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4431 gpout1.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5176 _00670_ vssd1 vssd1 vccd1 vccd1 net5700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5187 _00684_ vssd1 vssd1 vccd1 vccd1 net5711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4442 _01648_ vssd1 vssd1 vccd1 vccd1 net4966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4453 net708 vssd1 vssd1 vccd1 vccd1 net4977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5198 _00701_ vssd1 vssd1 vccd1 vccd1 net5722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4464 _01589_ vssd1 vssd1 vccd1 vccd1 net4988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3730 net7662 vssd1 vssd1 vccd1 vccd1 net4254 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold4475 net803 vssd1 vssd1 vccd1 vccd1 net4999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3741 net1600 vssd1 vssd1 vccd1 vccd1 net4265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4486 rbzero.spi_registers.buf_texadd0\[15\] vssd1 vssd1 vccd1 vccd1 net5010 sky130_fd_sc_hd__dlygate4sd3_1
X_22066_ clknet_leaf_7_i_clk net3479 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3752 _00483_ vssd1 vssd1 vccd1 vccd1 net4276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4497 rbzero.spi_registers.texadd1\[7\] vssd1 vssd1 vccd1 vccd1 net5021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3763 net1101 vssd1 vssd1 vccd1 vccd1 net4287 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03983_ clknet_0__03983_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03983_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3774 net7519 vssd1 vssd1 vccd1 vccd1 net4298 sky130_fd_sc_hd__dlygate4sd3_1
X_21017_ _04019_ _04020_ _04016_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a21bo_1
Xhold3785 net7804 vssd1 vssd1 vccd1 vccd1 net4309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3796 net644 vssd1 vssd1 vccd1 vccd1 net4320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13770_ _06668_ _06736_ _06918_ _06916_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__or4_2
X_10982_ net2134 net6646 _04366_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_40_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12721_ net57 _05854_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__a21o_1
X_21919_ clknet_leaf_93_i_clk net1307 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15440_ _08497_ _08514_ vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__or2_1
X_12652_ _05790_ net6 _05807_ _05810_ _05813_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a311o_1
XFILLER_0_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _04714_ _04771_ _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__or3_1
X_15371_ _08426_ _08445_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12583_ _04984_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17110_ _10110_ _10111_ vssd1 vssd1 vccd1 vccd1 _10112_ sky130_fd_sc_hd__nand2_1
X_14322_ _07470_ _07472_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18090_ _02130_ _02038_ _02136_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__and3_1
X_11534_ _04701_ _04704_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _10045_ _10046_ _10047_ vssd1 vssd1 vccd1 vccd1 _10048_ sky130_fd_sc_hd__o21ai_1
X_14253_ _07356_ _07354_ _07401_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11465_ _04599_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__buf_4
Xhold7090 rbzero.wall_tracer.rayAddendX\[-8\] vssd1 vssd1 vccd1 vccd1 net7614 sky130_fd_sc_hd__dlygate4sd3_1
X_13204_ _06216_ _06185_ _06190_ _06219_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ _07325_ _07334_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11396_ net7276 net7219 _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__mux2_1
X_13135_ _06286_ _06288_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18992_ net3747 net3213 net2978 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__and3_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _10257_ _09805_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__or2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ net6216 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__clkbuf_4
X_12017_ net4076 _04975_ _05180_ _05181_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17874_ _01812_ _09861_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19613_ net5121 net799 _03342_ _03343_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__o211a_1
X_16825_ _09893_ _09894_ vssd1 vssd1 vccd1 vccd1 _09895_ sky130_fd_sc_hd__or2_4
XFILLER_0_75_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19544_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__clkbuf_2
X_16756_ _09711_ _09714_ _09825_ vssd1 vssd1 vccd1 vccd1 _09826_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13968_ _07113_ _07117_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__o21a_1
X_15707_ _08721_ _08720_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19475_ net3125 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__clkbuf_1
X_12919_ _06070_ _06074_ _06075_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and3_1
X_16687_ _09581_ _09625_ _09624_ vssd1 vssd1 vccd1 vccd1 _09758_ sky130_fd_sc_hd__a21oi_1
X_13899_ _07047_ _07048_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18426_ _02452_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__or2b_1
X_15638_ _08433_ _08516_ _08711_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18357_ net7801 _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__nor2_1
X_15569_ _08643_ _08632_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17308_ _10307_ _10308_ vssd1 vssd1 vccd1 vccd1 _10309_ sky130_fd_sc_hd__xor2_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18288_ _02333_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17239_ _10238_ _10239_ vssd1 vssd1 vccd1 vccd1 _10240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold902 _01507_ vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _01288_ vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20250_ net3646 _03743_ _03752_ _03748_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__o211a_1
Xhold924 net6519 vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 net5858 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 net5174 vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 net6474 vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
X_20181_ net5481 _03704_ _03713_ _03709_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__o211a_1
Xhold968 net5440 vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3004 net4585 vssd1 vssd1 vccd1 vccd1 net3528 sky130_fd_sc_hd__buf_1
XFILLER_0_110_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold979 _01395_ vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3015 net6122 vssd1 vssd1 vccd1 vccd1 net3539 sky130_fd_sc_hd__buf_2
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3026 _01201_ vssd1 vssd1 vccd1 vccd1 net3550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3037 net4843 vssd1 vssd1 vccd1 vccd1 net3561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2303 net7279 vssd1 vssd1 vccd1 vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3048 rbzero.pov.ready_buffer\[45\] vssd1 vssd1 vccd1 vccd1 net3572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3059 _01224_ vssd1 vssd1 vccd1 vccd1 net3583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2314 net6083 vssd1 vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2325 _04259_ vssd1 vssd1 vccd1 vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2336 _01276_ vssd1 vssd1 vccd1 vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 _04349_ vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2347 _04416_ vssd1 vssd1 vccd1 vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 _04515_ vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 net6909 vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _01163_ vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 _03556_ vssd1 vssd1 vccd1 vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1635 net4680 vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 _04263_ vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1657 _01290_ vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 net5936 vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 net7047 vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21704_ clknet_leaf_1_i_clk net4609 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21635_ clknet_leaf_32_i_clk net3183 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21566_ clknet_leaf_17_i_clk net5138 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20517_ net3249 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21497_ clknet_leaf_14_i_clk net2775 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11250_ net1881 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20448_ _03836_ net3548 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ net2250 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20379_ net3189 net1204 _03782_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__mux2_1
Xhold4250 _01015_ vssd1 vssd1 vccd1 vccd1 net4774 sky130_fd_sc_hd__dlygate4sd3_1
X_22118_ net250 net2798 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4261 _00425_ vssd1 vssd1 vccd1 vccd1 net4785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4272 _03655_ vssd1 vssd1 vccd1 vccd1 net4796 sky130_fd_sc_hd__buf_1
Xhold4283 _01638_ vssd1 vssd1 vccd1 vccd1 net4807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4294 _02908_ vssd1 vssd1 vccd1 vccd1 net4818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3560 _08281_ vssd1 vssd1 vccd1 vccd1 net4084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14940_ net4382 _08086_ _08027_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__mux2_1
X_22049_ clknet_leaf_91_i_clk net3443 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3571 _05203_ vssd1 vssd1 vccd1 vccd1 net4095 sky130_fd_sc_hd__buf_4
Xhold3582 _09909_ vssd1 vssd1 vccd1 vccd1 net4106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3593 net699 vssd1 vssd1 vccd1 vccd1 net4117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2870 _02400_ vssd1 vssd1 vccd1 vccd1 net3394 sky130_fd_sc_hd__clkdlybuf4s25_1
X_14871_ _06664_ _06678_ _08021_ net7566 vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__a31o_1
Xhold2892 net4927 vssd1 vssd1 vccd1 vccd1 net3416 sky130_fd_sc_hd__dlygate4sd3_1
X_16610_ _09673_ _09679_ vssd1 vssd1 vccd1 vccd1 _09681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13822_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__buf_6
X_17590_ _10474_ _10586_ _10587_ vssd1 vssd1 vccd1 vccd1 _10588_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _09604_ _09612_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__xnor2_1
X_13753_ _06846_ _06898_ net554 vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a21oi_2
X_10965_ net6512 net6836 _04355_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ net14 net15 _05861_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and4b_1
X_19260_ net5011 _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__or2_1
X_16472_ _09448_ _09450_ _09446_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_183_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13684_ _06743_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__or2_1
X_10896_ net6413 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__clkbuf_1
X_18211_ _02256_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nand2_1
X_15423_ _08497_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__buf_2
X_12635_ net54 _05786_ _05796_ net55 vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19191_ net2997 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18142_ _01812_ _10416_ _02101_ _02099_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15354_ _08080_ _08085_ _08295_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__a21o_1
X_12566_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _05014_ vssd1 vssd1 vccd1 vccd1 _05731_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14305_ _07417_ _07455_ _07422_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__o21a_1
X_11517_ _04643_ _04687_ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18073_ _10383_ _09805_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nor2_1
X_15285_ net3206 _08297_ _08307_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__a21oi_1
X_12497_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _05263_ vssd1 vssd1 vccd1 vccd1 _05663_
+ sky130_fd_sc_hd__mux2_1
X_20783__209 clknet_1_0__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__inv_2
X_17024_ _10026_ _10024_ _10025_ vssd1 vssd1 vccd1 vccd1 _10032_ sky130_fd_sc_hd__a21boi_2
X_14236_ _07322_ _07364_ _07385_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__or3_1
Xhold209 rbzero.pov.ready_buffer\[59\] vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__buf_4
XFILLER_0_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ _07314_ _07317_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11379_ net6351 net2656 _04573_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ net3742 vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__inv_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _07191_ _07245_ _07247_ _07248_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__or4_4
X_18975_ _02261_ _09954_ _02951_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a31o_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13049_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__clkbuf_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ net4599 net4530 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20978__386 clknet_1_0__leaf__04010_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__inv_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ _01820_ _01878_ _01905_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20677__114 clknet_1_0__leaf__03981_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__inv_2
X_16808_ _08613_ _09877_ _09741_ _09742_ _09734_ vssd1 vssd1 vccd1 vccd1 _09878_ sky130_fd_sc_hd__a32o_1
X_17788_ _01837_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19527_ net1608 _03289_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
X_16739_ _09677_ _09808_ vssd1 vssd1 vccd1 vccd1 _09809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19458_ _02998_ _03241_ net1532 _03233_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18409_ net4458 net5684 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _03141_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21420_ clknet_leaf_85_i_clk net4814 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21351_ clknet_leaf_39_i_clk net4157 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 net6420 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
X_21282_ clknet_leaf_62_i_clk _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold721 net5208 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold732 net5606 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 net6440 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_20233_ net5432 _03730_ _03742_ _03735_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 net5113 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 net5518 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 net5628 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 net5610 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
X_20164_ net5575 _03691_ _03703_ _03696_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__o211a_1
Xhold798 net3645 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2100 _01504_ vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2111 net7174 vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2122 _01494_ vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 _04577_ vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2144 net7283 vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ net2937 net4796 _03659_ net4968 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__or4b_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _01520_ vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2155 net7120 vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2166 _04260_ vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 net6667 vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2177 _01533_ vssd1 vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1432 net2023 vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1443 net2288 vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2188 _04574_ vssd1 vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2199 net7248 vssd1 vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 _01510_ vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1465 net600 vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1476 net4755 vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _04297_ vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 _00919_ vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ net2367 net5942 _04244_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ net5981 net6419 _04203_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _05019_ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21618_ clknet_leaf_17_i_clk net5104 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12351_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _04986_ vssd1 vssd1 vccd1 vccd1 _05519_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21549_ clknet_leaf_3_i_clk net4151 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ net2290 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _08197_
+ sky130_fd_sc_hd__inv_2
X_12282_ _05106_ _05449_ _05104_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o21ai_1
X_14021_ _07169_ _07170_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__a21bo_1
X_11233_ net1384 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ net6886 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4080 net7902 vssd1 vssd1 vccd1 vccd1 net4604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4091 net1587 vssd1 vssd1 vccd1 vccd1 net4615 sky130_fd_sc_hd__dlygate4sd3_1
X_18760_ _02752_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15972_ _09044_ _09046_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__nand2_1
X_11095_ net6459 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17711_ _01760_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__nor2_1
Xhold3390 _02974_ vssd1 vssd1 vccd1 vccd1 net3914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14923_ _08069_ _08070_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__nand2_1
X_18691_ _02676_ net3242 _02677_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 net1562 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 net4122 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _01692_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__nand2_1
Xhold92 net3037 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _06664_ _08001_ _08004_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__a21o_1
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ _06931_ _06955_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17573_ _10010_ _10460_ _10461_ _10571_ vssd1 vssd1 vccd1 vccd1 _10572_ sky130_fd_sc_hd__o31ai_1
X_14785_ _07924_ _07927_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__xnor2_1
X_11997_ _05161_ _04604_ _04776_ _05162_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19312_ net5614 _03159_ _03163_ _03155_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__o211a_1
X_16524_ _09375_ _09482_ _08584_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__a21o_1
X_10948_ net5854 net5897 _04344_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
X_13736_ _06880_ _06881_ _06884_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__nand4_4
XFILLER_0_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19243_ net5222 _03120_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__or2_1
X_16455_ net7407 _09526_ _08633_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10879_ net5913 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__clkbuf_1
X_13667_ _06724_ _06765_ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__and3_1
XFILLER_0_171_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15406_ _08479_ _08480_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ _05781_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
X_19174_ net5783 _03079_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _09456_ _09457_ vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__and2_1
X_13598_ _06747_ _06748_ _06676_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18125_ _02172_ net4497 _01749_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
X_12549_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _04994_ vssd1 vssd1 vccd1 vccd1 _05714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15337_ net3003 net4294 _08375_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__or3_1
XFILLER_0_152_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5709 net1661 vssd1 vssd1 vccd1 vccd1 net6233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18056_ _02041_ _02042_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__nand2_1
XANTENNA_1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15268_ net4306 net4335 vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__and2_1
X_17007_ _10015_ _10016_ vssd1 vssd1 vccd1 vccd1 _10017_ sky130_fd_sc_hd__or2b_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ _07368_ _07369_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15199_ _08279_ net4066 vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18958_ _02934_ _02935_ _02933_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__o21a_1
XFILLER_0_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17909_ _01849_ _01851_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__and2b_1
X_18889_ rbzero.wall_tracer.rayAddendY\[4\] _02875_ _02714_ vssd1 vssd1 vccd1 vccd1
+ _02876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer13 _07141_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_1
Xrebuffer24 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 _07231_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_2
Xrebuffer46 _07035_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_1
Xrebuffer57 net584 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer68 _06886_ vssd1 vssd1 vccd1 vccd1 net3246 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22452_ clknet_leaf_46_i_clk net651 vssd1 vssd1 vccd1 vccd1 reg_hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20731__163 clknet_1_0__leaf__03986_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__inv_2
X_21403_ clknet_leaf_65_i_clk _00572_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_22383_ net515 net1181 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6922 net4358 vssd1 vssd1 vccd1 vccd1 net7446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6933 net7568 vssd1 vssd1 vccd1 vccd1 net7457 sky130_fd_sc_hd__clkbuf_2
Xhold6944 net3504 vssd1 vssd1 vccd1 vccd1 net7468 sky130_fd_sc_hd__dlygate4sd3_1
X_21334_ clknet_leaf_54_i_clk net5381 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6955 rbzero.wall_tracer.stepDistX\[2\] vssd1 vssd1 vccd1 vccd1 net7479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6966 rbzero.wall_tracer.trackDistY\[6\] vssd1 vssd1 vccd1 vccd1 net7490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6977 rbzero.traced_texVinit\[4\] vssd1 vssd1 vccd1 vccd1 net7501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6999 rbzero.wall_tracer.trackDistY\[-10\] vssd1 vssd1 vccd1 vccd1 net7523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 net5509 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21265_ clknet_leaf_71_i_clk net4831 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold551 _01342_ vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold562 net5451 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
X_20216_ net5387 _03730_ _03733_ _03722_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold573 net5488 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold584 _03946_ vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21196_ _02529_ _02755_ net4622 _02528_ net738 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a32o_1
Xhold595 net5524 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20147_ net5554 _03691_ _03694_ _03683_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__o211a_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _03616_ net3701 vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__or2_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1240 _01561_ vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 net6761 vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _05088_ _05089_ _04982_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__mux2_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1262 _00917_ vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 net6683 vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1284 _00910_ vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 net6829 vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _04959_ _04971_ _04976_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__or3_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ net7173 net6828 _04266_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14570_ _07674_ _07720_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _04947_ _04950_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__or3_2
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10733_ net5857 net1458 _04225_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_1
X_13521_ _06584_ _06586_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _09309_ _09313_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _06601_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__xnor2_2
X_10664_ net5811 net5798 _04192_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12403_ rbzero.tex_g1\[15\] rbzero.tex_g1\[14\] _05263_ vssd1 vssd1 vccd1 vccd1 _05570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16171_ _09242_ _09244_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13383_ _06533_ _06476_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__nor2_1
X_12334_ _05500_ _05501_ _04992_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15122_ net6148 _08223_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19930_ _08464_ _03476_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__nor2_1
X_15053_ net4380 _08184_ _08138_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12265_ net7369 _05382_ _05379_ net2933 vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__a22o_1
X_14004_ _07150_ _07154_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nand2_1
X_11216_ net2207 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
X_19861_ _03440_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__clkbuf_4
X_12196_ _05348_ _05345_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nor2_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__buf_1
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18812_ _05396_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ net6572 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
X_19792_ net5861 _03443_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ net3894 _06183_ _06394_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11078_ net2238 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
X_15955_ _09013_ _09029_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__xor2_1
XFILLER_0_208_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14906_ _08006_ _08021_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__nand2_1
X_18674_ _02646_ net4463 net3242 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__or3b_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _08391_ _08392_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__nand2_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _10259_ _08630_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__nor2_1
X_14837_ _07493_ _07982_ _07987_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__nand3_2
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ _10553_ _10554_ vssd1 vssd1 vccd1 vccd1 _10555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14768_ _07534_ _07590_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16507_ _09569_ _09578_ vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__xor2_2
X_13719_ _06869_ _06858_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__nor2_1
X_17487_ _10360_ _10361_ _10359_ vssd1 vssd1 vccd1 vccd1 _10486_ sky130_fd_sc_hd__a21o_1
X_14699_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20789__215 clknet_1_1__leaf__03992_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__inv_2
X_19226_ net5072 _03107_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__or2_1
X_16438_ _09415_ _09416_ _09509_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6207 rbzero.tex_b0\[14\] vssd1 vssd1 vccd1 vccd1 net6731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19157_ net5243 _03066_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__or2_1
Xhold6218 net1815 vssd1 vssd1 vccd1 vccd1 net6742 sky130_fd_sc_hd__dlygate4sd3_1
X_16369_ _09440_ _09441_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6229 _04340_ vssd1 vssd1 vccd1 vccd1 net6753 sky130_fd_sc_hd__dlygate4sd3_1
X_18108_ _02154_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__nor2_1
Xhold5506 _00894_ vssd1 vssd1 vccd1 vccd1 net6030 sky130_fd_sc_hd__dlygate4sd3_1
X_19088_ net4884 _03026_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__and2_1
Xhold5517 net3929 vssd1 vssd1 vccd1 vccd1 net6041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5528 _03457_ vssd1 vssd1 vccd1 vccd1 net6052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5539 _03388_ vssd1 vssd1 vccd1 vccd1 net6063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4805 rbzero.color_floor\[0\] vssd1 vssd1 vccd1 vccd1 net5329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18039_ _01833_ _02025_ _02085_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4816 net1026 vssd1 vssd1 vccd1 vccd1 net5340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4827 _00867_ vssd1 vssd1 vccd1 vccd1 net5351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4838 net963 vssd1 vssd1 vccd1 vccd1 net5362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4849 net994 vssd1 vssd1 vccd1 vccd1 net5373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21050_ net4152 net4763 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20001_ _03261_ net3901 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__or2_1
X_20761__189 clknet_1_0__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__inv_2
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21952_ net177 net2811 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21883_ clknet_leaf_99_i_clk net5502 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22435_ clknet_leaf_38_i_clk net4471 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6730 rbzero.tex_g0\[19\] vssd1 vssd1 vccd1 vccd1 net7254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7475 rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 net7999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22366_ net498 net1685 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold6741 rbzero.tex_r1\[17\] vssd1 vssd1 vccd1 vccd1 net7265 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__04002_ clknet_0__04002_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04002_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7486 _09282_ vssd1 vssd1 vccd1 vccd1 net8010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6752 net2809 vssd1 vssd1 vccd1 vccd1 net7276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6763 rbzero.tex_g1\[41\] vssd1 vssd1 vccd1 vccd1 net7287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6774 net2881 vssd1 vssd1 vccd1 vccd1 net7298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21317_ clknet_leaf_73_i_clk net4266 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6785 net2902 vssd1 vssd1 vccd1 vccd1 net7309 sky130_fd_sc_hd__dlygate4sd3_1
X_22297_ net429 net2294 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
X_12050_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__clkbuf_8
Xhold370 net5235 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
X_21248_ clknet_leaf_54_i_clk net3208 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold381 net5323 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net2514 net6343 _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
Xhold392 net5331 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
X_21179_ net4231 _04140_ _04141_ _10454_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15740_ _08754_ _08631_ _08811_ _08813_ _08814_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__a32oi_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__inv_2
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 net5744 vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _03368_ vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _05072_ vssd1 vssd1 vccd1 vccd1 _05073_
+ sky130_fd_sc_hd__mux2_1
Xhold1092 net6560 vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _08697_ _08745_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__xnor2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _06036_ _06037_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a21o_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _10408_ _10409_ vssd1 vssd1 vccd1 vccd1 _10410_ sky130_fd_sc_hd__nand2_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20738__169 clknet_1_1__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__inv_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _07618_ _07400_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__nor2_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__buf_4
X_18390_ _09987_ _02421_ net3236 _10330_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a31o_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _10250_ _10338_ _10339_ vssd1 vssd1 vccd1 vccd1 _10341_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ net869 net1529 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__or2_1
X_14553_ _07702_ _07703_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ net6882 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13504_ _06652_ _06640_ _06650_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__a22o_1
X_17272_ _10269_ _10271_ vssd1 vssd1 vccd1 vccd1 _10273_ sky130_fd_sc_hd__nand2_1
X_14484_ _07595_ _07614_ _07612_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__a21o_1
X_11696_ _04801_ net2536 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19011_ _02979_ _02967_ net3886 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and3b_1
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16223_ _09292_ _09293_ net7407 vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10647_ net6564 net7006 _04181_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _06576_ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer4 _07156_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_1
X_16154_ _09227_ _09228_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__xor2_2
X_13366_ _04635_ _06489_ _06491_ _06495_ _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15105_ net3186 net3174 _08219_ vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__mux2_1
X_12317_ _04993_ _05484_ _04999_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16085_ _09150_ _09155_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__nand2_1
X_13297_ _06446_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__nor2_2
X_12248_ net3786 _05381_ _05412_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a211o_1
X_19913_ net6082 _03530_ _08276_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o21ai_1
X_15036_ _08092_ _08148_ net7430 _06715_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__o211a_1
X_20903__317 clknet_1_0__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__inv_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19844_ net41 net40 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nor2_2
XFILLER_0_177_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12179_ net4010 _04616_ net3989 vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__mux2_2
X_19775_ net6164 _03427_ net2071 _03424_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16987_ net3508 vssd1 vssd1 vccd1 vccd1 _09999_ sky130_fd_sc_hd__buf_6
X_18726_ net3198 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_1
X_15938_ _08978_ _08979_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18657_ _02662_ _02663_ net4767 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__or3_1
X_15869_ _08940_ _08942_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__nand2_2
XFILLER_0_149_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ _01658_ _01657_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__and2b_1
X_18588_ net6117 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17539_ _10530_ _10537_ vssd1 vssd1 vccd1 vccd1 _10538_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20550_ net3483 net1265 _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19209_ net3130 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20481_ net3667 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
Xhold6004 _04373_ vssd1 vssd1 vccd1 vccd1 net6528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6015 net1435 vssd1 vssd1 vccd1 vccd1 net6539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6026 rbzero.tex_g1\[35\] vssd1 vssd1 vccd1 vccd1 net6550 sky130_fd_sc_hd__dlygate4sd3_1
X_22220_ net352 net2303 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6037 rbzero.spi_registers.buf_texadd1\[12\] vssd1 vssd1 vccd1 vccd1 net6561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5303 rbzero.tex_r1\[57\] vssd1 vssd1 vccd1 vccd1 net5827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6048 net1611 vssd1 vssd1 vccd1 vccd1 net6572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6059 _04353_ vssd1 vssd1 vccd1 vccd1 net6583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5314 net614 vssd1 vssd1 vccd1 vccd1 net5838 sky130_fd_sc_hd__clkbuf_2
Xhold5325 _04461_ vssd1 vssd1 vccd1 vccd1 net5849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22151_ net283 net2151 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5336 rbzero.spi_registers.buf_texadd3\[14\] vssd1 vssd1 vccd1 vccd1 net5860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5347 rbzero.tex_b1\[29\] vssd1 vssd1 vccd1 vccd1 net5871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4602 net868 vssd1 vssd1 vccd1 vccd1 net5126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5358 rbzero.spi_registers.vshift\[4\] vssd1 vssd1 vccd1 vccd1 net5882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4613 _00735_ vssd1 vssd1 vccd1 vccd1 net5137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4624 _00779_ vssd1 vssd1 vccd1 vccd1 net5148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5369 rbzero.tex_g1\[52\] vssd1 vssd1 vccd1 vccd1 net5893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21102_ net4186 net4469 vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4635 _00750_ vssd1 vssd1 vccd1 vccd1 net5159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22082_ clknet_leaf_79_i_clk net1109 vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
Xhold3901 _02533_ vssd1 vssd1 vccd1 vccd1 net4425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4646 net860 vssd1 vssd1 vccd1 vccd1 net5170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4657 rbzero.spi_registers.texadd1\[12\] vssd1 vssd1 vccd1 vccd1 net5181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3912 net7521 vssd1 vssd1 vccd1 vccd1 net4436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold3923 _03624_ vssd1 vssd1 vccd1 vccd1 net4447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4668 rbzero.pov.spi_buffer\[44\] vssd1 vssd1 vccd1 vccd1 net5192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20843__264 clknet_1_0__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__inv_2
Xhold3934 net3209 vssd1 vssd1 vccd1 vccd1 net4458 sky130_fd_sc_hd__buf_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4679 net816 vssd1 vssd1 vccd1 vccd1 net5203 sky130_fd_sc_hd__dlygate4sd3_1
X_21033_ net5379 net5168 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__nand2_1
Xhold3945 net1583 vssd1 vssd1 vccd1 vccd1 net4469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3956 _00577_ vssd1 vssd1 vccd1 vccd1 net4480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3967 net3373 vssd1 vssd1 vccd1 vccd1 net4491 sky130_fd_sc_hd__buf_1
Xhold3978 rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 net4502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3989 net3433 vssd1 vssd1 vccd1 vccd1 net4513 sky130_fd_sc_hd__buf_1
XFILLER_0_201_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20983__10 clknet_1_0__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
XFILLER_0_59_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21935_ clknet_leaf_9_i_clk net1361 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21866_ clknet_leaf_6_i_clk net4970 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21797_ clknet_leaf_11_i_clk net6184 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11550_ _04696_ _04697_ _04698_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11481_ rbzero.spi_registers.texadd3\[9\] rbzero.spi_registers.texadd1\[9\] rbzero.spi_registers.texadd0\[9\]
+ rbzero.spi_registers.texadd2\[9\] rbzero.wall_hot\[1\] rbzero.wall_hot\[0\] vssd1
+ vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__mux4_1
XFILLER_0_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _06221_ _06244_ _06373_ _06374_ _06375_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_162_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22418_ clknet_leaf_66_i_clk net667 vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold7272 _10027_ vssd1 vssd1 vccd1 vccd1 net7796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7283 rbzero.wall_tracer.stepDistX\[-10\] vssd1 vssd1 vccd1 vccd1 net7807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7294 _02379_ vssd1 vssd1 vccd1 vccd1 net7818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6560 rbzero.tex_r0\[12\] vssd1 vssd1 vccd1 vccd1 net7084 sky130_fd_sc_hd__dlygate4sd3_1
X_13151_ net4483 _06305_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__o21ba_1
Xhold6571 net2265 vssd1 vssd1 vccd1 vccd1 net7095 sky130_fd_sc_hd__dlygate4sd3_1
X_22349_ net481 net2103 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
Xhold6582 rbzero.tex_b1\[37\] vssd1 vssd1 vccd1 vccd1 net7106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ rbzero.tex_r1\[5\] rbzero.tex_r1\[4\] _05072_ vssd1 vssd1 vccd1 vccd1 _05271_
+ sky130_fd_sc_hd__mux2_1
Xhold6593 net2293 vssd1 vssd1 vccd1 vccd1 net7117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5870 rbzero.tex_r0\[54\] vssd1 vssd1 vccd1 vccd1 net6394 sky130_fd_sc_hd__dlygate4sd3_1
X_13082_ _06226_ net4874 _06228_ _06237_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a211o_1
Xhold5881 net1160 vssd1 vssd1 vccd1 vccd1 net6405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5892 _04367_ vssd1 vssd1 vccd1 vccd1 net6416 sky130_fd_sc_hd__dlygate4sd3_1
X_12033_ net83 _05191_ net4044 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__o21a_1
X_16910_ net4167 _09939_ _09940_ net6259 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__a22o_1
X_17890_ _01938_ _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _09908_ net4107 vssd1 vssd1 vccd1 vccd1 _09911_ sky130_fd_sc_hd__xnor2_1
X_19560_ _03000_ _03305_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__or2_1
X_16772_ _09840_ _09841_ vssd1 vssd1 vccd1 vccd1 _09842_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13984_ _07120_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18511_ _09935_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__clkbuf_4
X_15723_ _08797_ _08709_ _08703_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ _02996_ _03265_ net2554 _03260_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ _06053_ _06064_ _06090_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__o31a_2
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18442_ net4437 net4380 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__or2_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _08725_ _08726_ _08727_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _04760_ _04603_ _04637_ _04165_ net28 net29 vssd1 vssd1 vccd1 vccd1 _06024_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14605_ _07366_ _07589_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__nor2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11817_ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__buf_4
X_18373_ _02399_ net3395 net3234 _02407_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ net3722 _08327_ _08379_ _08579_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__or4b_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _05955_ net22 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__and2_2
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _10213_ _10214_ _10323_ vssd1 vssd1 vccd1 vccd1 _10325_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _07651_ _07666_ _07686_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__o21ai_2
X_11748_ net785 net2467 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17255_ _10151_ _10160_ vssd1 vssd1 vccd1 vccd1 _10256_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__03993_ _03993_ vssd1 vssd1 vccd1 vccd1 clknet_0__03993_ sky130_fd_sc_hd__clkbuf_16
X_14467_ _06922_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11679_ _04846_ _04726_ net2986 _04847_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16206_ _09181_ _09183_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__xor2_4
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ _06479_ _06568_ _06433_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__o21a_1
X_17186_ _10186_ _10187_ vssd1 vssd1 vccd1 vccd1 _10188_ sky130_fd_sc_hd__xor2_2
XFILLER_0_52_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14398_ _07525_ _07526_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16137_ _08564_ _08684_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13349_ _06445_ _06458_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16068_ _09129_ _09136_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__nor2_1
Xhold3208 net6007 vssd1 vssd1 vccd1 vccd1 net3732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3219 rbzero.pov.ready_buffer\[25\] vssd1 vssd1 vccd1 vccd1 net3743 sky130_fd_sc_hd__buf_1
X_15019_ _08156_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
Xhold2507 _03490_ vssd1 vssd1 vccd1 vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2518 net7907 vssd1 vssd1 vccd1 vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2529 _00637_ vssd1 vssd1 vccd1 vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1806 _01544_ vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
X_19827_ _03468_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
Xhold1817 net6863 vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 net7673 vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1839 net7152 vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19758_ _02491_ _02500_ _02514_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__and3_2
X_18709_ _02556_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__buf_4
XFILLER_0_190_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19689_ net4672 _03361_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21720_ clknet_leaf_8_i_clk net1627 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21651_ clknet_leaf_16_i_clk net5257 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_otherx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20602_ net6365 _03026_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21582_ clknet_leaf_21_i_clk net5662 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20533_ net3360 net1337 _03889_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20464_ _03836_ net3765 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5100 _01089_ vssd1 vssd1 vccd1 vccd1 net5624 sky130_fd_sc_hd__dlygate4sd3_1
X_22203_ net335 net1193 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5111 net1369 vssd1 vssd1 vccd1 vccd1 net5635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5122 net1475 vssd1 vssd1 vccd1 vccd1 net5646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5133 _00685_ vssd1 vssd1 vccd1 vccd1 net5657 sky130_fd_sc_hd__dlygate4sd3_1
X_20395_ net3319 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5144 rbzero.spi_registers.texadd0\[2\] vssd1 vssd1 vccd1 vccd1 net5668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5155 _00681_ vssd1 vssd1 vccd1 vccd1 net5679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4410 _08267_ vssd1 vssd1 vccd1 vccd1 net4934 sky130_fd_sc_hd__dlygate4sd3_1
X_22134_ net266 net2589 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
X_20767__195 clknet_1_1__leaf__03990_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__inv_2
Xhold5166 net1415 vssd1 vssd1 vccd1 vccd1 net5690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4421 net666 vssd1 vssd1 vccd1 vccd1 net4945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5177 rbzero.floor_leak\[4\] vssd1 vssd1 vccd1 vccd1 net5701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4432 net660 vssd1 vssd1 vccd1 vccd1 net4956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4443 rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 net4967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5188 net1525 vssd1 vssd1 vccd1 vccd1 net5712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4454 rbzero.spi_registers.texadd3\[21\] vssd1 vssd1 vccd1 vccd1 net4978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5199 rbzero.spi_registers.texadd1\[23\] vssd1 vssd1 vccd1 vccd1 net5723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4465 net718 vssd1 vssd1 vccd1 vccd1 net4989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3720 _03191_ vssd1 vssd1 vccd1 vccd1 net4244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3731 _00498_ vssd1 vssd1 vccd1 vccd1 net4255 sky130_fd_sc_hd__dlygate4sd3_1
X_22065_ clknet_leaf_7_i_clk net3491 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4476 _00788_ vssd1 vssd1 vccd1 vccd1 net5000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4487 net742 vssd1 vssd1 vccd1 vccd1 net5011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3742 _00486_ vssd1 vssd1 vccd1 vccd1 net4266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3753 net7942 vssd1 vssd1 vccd1 vccd1 net4277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4498 net813 vssd1 vssd1 vccd1 vccd1 net5022 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03982_ clknet_0__03982_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03982_
+ sky130_fd_sc_hd__clkbuf_16
X_21016_ _04016_ _04019_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__nand3b_1
Xhold3764 rbzero.debug_overlay.playerY\[-1\] vssd1 vssd1 vccd1 vccd1 net4288 sky130_fd_sc_hd__clkbuf_2
Xhold3775 net1012 vssd1 vssd1 vccd1 vccd1 net4299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3786 net3005 vssd1 vssd1 vccd1 vccd1 net4310 sky130_fd_sc_hd__buf_1
Xhold3797 rbzero.spi_registers.spi_buffer\[20\] vssd1 vssd1 vccd1 vccd1 net4321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10981_ net6417 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ net54 _05844_ _05852_ net55 vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21918_ clknet_leaf_93_i_clk net1396 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12651_ net6 _05812_ net7 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__and3b_1
X_21849_ clknet_leaf_81_i_clk net4617 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11602_ rbzero.spi_registers.texadd0\[1\] _04680_ _04772_ _04773_ _04724_ vssd1 vssd1
+ vccd1 vccd1 _04774_ sky130_fd_sc_hd__o221a_1
X_12582_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _05541_ vssd1 vssd1 vccd1 vccd1 _05747_
+ sky130_fd_sc_hd__mux2_1
X_15370_ _08433_ _08444_ vssd1 vssd1 vccd1 vccd1 _08445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20326__60 clknet_1_0__leaf__03777_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14321_ _07471_ _07464_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ _04160_ _04701_ _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ _10019_ _09403_ vssd1 vssd1 vccd1 vccd1 _10047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ _07401_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__xnor2_1
X_11464_ net4947 _04628_ _04630_ net3403 vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a31o_1
XFILLER_0_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20341__74 clknet_1_0__leaf__03778_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7091 rbzero.wall_tracer.rayAddendY\[-9\] vssd1 vssd1 vccd1 vccd1 net7615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _06346_ net4915 _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_208_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11395_ _04242_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__clkbuf_4
X_14183_ _07332_ _07333_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6390 net2402 vssd1 vssd1 vccd1 vccd1 net6914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ net3780 _06274_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and2_1
X_18991_ net3266 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__clkbuf_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _01989_ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__xnor2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ net6248 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12016_ net1402 _05027_ _04975_ net4076 _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17873_ _01921_ _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16824_ _09891_ _09892_ _09850_ vssd1 vssd1 vccd1 vccd1 _09894_ sky130_fd_sc_hd__a21oi_1
X_19612_ _03294_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19543_ _02491_ _02497_ _02500_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16755_ _09807_ _09824_ vssd1 vssd1 vccd1 vccd1 _09825_ sky130_fd_sc_hd__xnor2_1
X_13967_ _06862_ net573 vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15706_ _08779_ _08780_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__nand2_2
XFILLER_0_158_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19474_ _03088_ net3124 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or2_1
X_12918_ net53 _06065_ _06066_ net40 _06048_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__a221o_1
X_16686_ _09716_ _09756_ vssd1 vssd1 vccd1 vccd1 _09757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13898_ _06861_ net79 _06864_ _06844_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__or4b_1
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18425_ net4573 net4386 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15637_ _08433_ _08484_ _08711_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__or3_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12849_ net29 net28 vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_201_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18356_ _02391_ net3393 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _08320_ _08576_ _08578_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17307_ _10161_ _10183_ _10182_ vssd1 vssd1 vccd1 vccd1 _10308_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14519_ _07659_ _07665_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__xor2_4
X_18287_ _02332_ net4577 _01749_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_4
X_15499_ _08542_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17238_ _09311_ _09447_ vssd1 vssd1 vccd1 vccd1 _10239_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20909__323 clknet_1_1__leaf__04004_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__inv_2
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold903 net6511 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17169_ _09096_ _10168_ _10170_ vssd1 vssd1 vccd1 vccd1 _10171_ sky130_fd_sc_hd__or3b_1
Xhold914 net3650 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 net6521 vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _01527_ vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 net5495 vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _01267_ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
X_20180_ net3843 _03705_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__or2_1
Xhold969 net5431 vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3005 net5667 vssd1 vssd1 vccd1 vccd1 net3529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3016 _08198_ vssd1 vssd1 vccd1 vccd1 net3540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3038 _03652_ vssd1 vssd1 vccd1 vccd1 net3562 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2304 _04220_ vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3049 net2835 vssd1 vssd1 vccd1 vccd1 net3573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 net5972 vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__clkbuf_2
Xhold2326 _01509_ vssd1 vssd1 vccd1 vccd1 net2850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2337 net7303 vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1603 _01428_ vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 _01368_ vssd1 vssd1 vccd1 vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1614 _04185_ vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2359 _01278_ vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1625 net6763 vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1636 net7037 vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1647 _01505_ vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1658 net5961 vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1669 _01331_ vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
X_20955__365 clknet_1_0__leaf__04008_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__inv_2
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21703_ clknet_leaf_101_i_clk net5163 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21634_ clknet_leaf_34_i_clk net1597 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21565_ clknet_leaf_17_i_clk net5344 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20516_ net3613 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21496_ clknet_leaf_14_i_clk net4685 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20447_ net3547 net1335 _03823_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ net7042 net7046 _04470_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20378_ net3739 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4240 _01596_ vssd1 vssd1 vccd1 vccd1 net4764 sky130_fd_sc_hd__dlygate4sd3_1
X_22117_ net249 net2168 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold4251 rbzero.pov.ready_buffer\[12\] vssd1 vssd1 vccd1 vccd1 net4775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4262 net3056 vssd1 vssd1 vccd1 vccd1 net4786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4273 _03658_ vssd1 vssd1 vccd1 vccd1 net4797 sky130_fd_sc_hd__buf_1
Xhold4284 net914 vssd1 vssd1 vccd1 vccd1 net4808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4295 _00611_ vssd1 vssd1 vccd1 vccd1 net4819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3550 _05353_ vssd1 vssd1 vccd1 vccd1 net4074 sky130_fd_sc_hd__dlygate4sd3_1
X_22048_ clknet_leaf_91_i_clk net3304 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3561 _00461_ vssd1 vssd1 vccd1 vccd1 net4085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3572 _08277_ vssd1 vssd1 vccd1 vccd1 net4096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3583 _09910_ vssd1 vssd1 vccd1 vccd1 net4107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3594 net7622 vssd1 vssd1 vccd1 vccd1 net4118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2860 _03937_ vssd1 vssd1 vccd1 vccd1 net3384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2871 _02405_ vssd1 vssd1 vccd1 vccd1 net3395 sky130_fd_sc_hd__dlygate4sd3_1
X_14870_ _06690_ _08017_ _08020_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__a21o_1
Xhold2882 _02589_ vssd1 vssd1 vccd1 vccd1 net3406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2893 net3066 vssd1 vssd1 vccd1 vccd1 net3417 sky130_fd_sc_hd__clkbuf_2
X_13821_ _06846_ _06898_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__and2_4
XFILLER_0_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _09609_ _09611_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _06885_ net546 vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10964_ net1866 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12703_ net4043 _05853_ _05862_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a211o_1
X_16471_ _09429_ _09430_ _09428_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _06739_ _06833_ _06678_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__mux2_1
X_10895_ net2861 net6411 _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18210_ net3780 net4605 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__or2_1
X_15422_ _08328_ _08495_ _08496_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__o21a_2
X_19190_ _03088_ net2996 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12634_ net5 net4 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__and2b_2
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18141_ _02186_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15353_ _08295_ net7766 vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__nand2_1
X_12565_ _04983_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ _07423_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__inv_2
X_18072_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__nand2_1
X_11516_ rbzero.spi_registers.texadd3\[15\] rbzero.spi_registers.texadd1\[15\] rbzero.spi_registers.texadd0\[15\]
+ rbzero.spi_registers.texadd2\[15\] _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15284_ _08297_ _08358_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__or2_1
X_12496_ _05035_ _05657_ _05661_ _04979_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a211o_1
X_17023_ _10031_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ _07322_ _07364_ _07385_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11378_ net2204 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
X_14166_ _07315_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13117_ _06271_ net3369 _06272_ net3852 vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a22o_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _07227_ _07229_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__nor2_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _04823_ _02261_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__nor2_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ net4911 vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__buf_4
X_17925_ net4599 net4530 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ _01820_ _01878_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _09873_ _09738_ _09305_ vssd1 vssd1 vccd1 vccd1 _09877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17787_ _01832_ _01836_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__or2_1
X_14999_ _08139_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
X_16738_ _09674_ _09678_ vssd1 vssd1 vccd1 vccd1 _09808_ sky130_fd_sc_hd__or2b_1
X_19526_ net5247 _03288_ _03290_ _03280_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19457_ _02492_ _02498_ _03238_ net6229 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16669_ net3127 _09486_ vssd1 vssd1 vccd1 vccd1 _09740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18408_ net4458 net5684 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nand2_1
X_19388_ net1115 _03199_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18339_ _02376_ _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__or2b_1
XFILLER_0_189_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20305__41 clknet_1_0__leaf__03775_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
X_21350_ clknet_leaf_39_i_clk net4138 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold700 net3683 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
X_21281_ clknet_leaf_71_i_clk _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold711 net6422 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20320__55 clknet_1_1__leaf__03776_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
Xhold722 net5210 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 net7718 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_1
X_20232_ net3275 _03731_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_1
Xhold744 net6442 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 net5115 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold766 net5192 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold777 net5630 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 net5677 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
X_20163_ net5540 _03692_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold799 _01092_ vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2101 net7166 vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2112 _04207_ vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2123 net2685 vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
X_20094_ net3825 net1601 net2628 net3328 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or4b_1
Xhold2134 _01128_ vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 net6737 vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2145 _04281_ vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2156 _04251_ vssd1 vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 net6965 vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_54_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2167 _01508_ vssd1 vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _01356_ vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 net5835 vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2178 net7265 vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1444 net5818 vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2189 _01131_ vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 net6777 vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
X_20879__296 clknet_1_0__leaf__04001_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__inv_2
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1466 _03446_ vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1477 net2233 vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1488 _01474_ vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 rbzero.tex_g0\[33\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10680_ net2636 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21617_ clknet_leaf_25_i_clk net5692 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12350_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _05493_ vssd1 vssd1 vccd1 vccd1 _05518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21548_ clknet_leaf_3_i_clk net4123 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ net2289 net7038 _04529_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_1
X_12281_ net4239 _05102_ _05097_ _05004_ _05010_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21479_ clknet_leaf_1_i_clk net4320 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11232_ net5962 net6504 _04492_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__mux2_1
X_14020_ _06826_ _06861_ _06864_ _06885_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ net2212 net6884 _04459_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4070 net7546 vssd1 vssd1 vccd1 vccd1 net4594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4081 net3565 vssd1 vssd1 vccd1 vccd1 net4605 sky130_fd_sc_hd__dlygate4sd3_1
X_15971_ _08432_ _08626_ _09022_ _09045_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__a2bb2o_1
X_11094_ net6457 net2527 _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
Xhold4092 _01018_ vssd1 vssd1 vccd1 vccd1 net4616 sky130_fd_sc_hd__dlygate4sd3_1
X_17710_ _01668_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3380 net7356 vssd1 vssd1 vccd1 vccd1 net3904 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3391 _02975_ vssd1 vssd1 vccd1 vccd1 net3915 sky130_fd_sc_hd__dlygate4sd3_1
X_14922_ net7434 _08017_ _08042_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__a21bo_1
X_18690_ _02647_ net3242 _05401_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__or3b_4
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 _03195_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _01682_ _01691_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__or2_1
Xhold2690 _02525_ vssd1 vssd1 vccd1 vccd1 net3214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net5349 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _06664_ _08003_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__nor2_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 net5797 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _06882_ _06885_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__xor2_4
X_17572_ _10462_ _10464_ _10568_ _10570_ vssd1 vssd1 vccd1 vccd1 _10571_ sky130_fd_sc_hd__a31o_2
X_14784_ _07933_ _07934_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__and2_1
XFILLER_0_212_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11996_ _05122_ net3987 net3908 _05162_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__o221a_1
X_19311_ net1692 _03160_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or2_1
X_16523_ _09364_ vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13735_ net579 _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__xnor2_4
X_10947_ net2126 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19242_ net5230 _03119_ _03123_ _03115_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__o211a_1
X_16454_ net7407 _09526_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13666_ _06731_ _06816_ _06717_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__mux2_1
X_10878_ net5911 net5775 _04310_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15405_ net3028 _08439_ net4105 vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__o21ai_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19173_ net5702 _03078_ _03081_ _03074_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__o211a_1
X_12617_ reg_vsync _04620_ _05204_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__mux2_2
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _09456_ _09457_ vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _06595_ _06667_ _06686_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _09987_ net7815 _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a21o_1
X_15336_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__clkbuf_4
X_12548_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _04989_ vssd1 vssd1 vccd1 vccd1 _05713_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18055_ _02101_ _02102_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15267_ net4306 net4335 vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__nor2_1
X_12479_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _05262_ vssd1 vssd1 vccd1 vccd1 _05645_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17006_ net4528 net4727 vssd1 vssd1 vccd1 vccd1 _10016_ sky130_fd_sc_hd__nand2_1
X_14218_ _06737_ net543 _07366_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__or3_1
X_15198_ _08275_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _07296_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ net3085 _02557_ _09943_ _02936_ _02938_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__o221a_1
XFILLER_0_207_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17908_ _01876_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18888_ _02866_ _02874_ _04632_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__mux2_1
X_17839_ _01887_ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__xor2_2
Xrebuffer14 _06530_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_1
Xrebuffer25 _07112_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 _07249_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_2
Xrebuffer47 _07076_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_1
Xrebuffer58 _06780_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer69 net3246 vssd1 vssd1 vccd1 vccd1 net3333 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_7_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19509_ net5110 _03274_ _03279_ _03280_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7602 _06146_ vssd1 vssd1 vccd1 vccd1 net8126 sky130_fd_sc_hd__dlygate4sd3_1
X_22451_ clknet_leaf_65_i_clk _01620_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21402_ clknet_leaf_65_i_clk _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_22382_ net514 net2495 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6912 _06765_ vssd1 vssd1 vccd1 vccd1 net7436 sky130_fd_sc_hd__buf_1
Xhold6923 _09770_ vssd1 vssd1 vccd1 vccd1 net7447 sky130_fd_sc_hd__dlygate4sd3_1
X_21333_ clknet_leaf_54_i_clk net4204 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6934 _06800_ vssd1 vssd1 vccd1 vccd1 net7458 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6956 net4348 vssd1 vssd1 vccd1 vccd1 net7480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6967 rbzero.traced_texVinit\[6\] vssd1 vssd1 vccd1 vccd1 net7491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6978 net4163 vssd1 vssd1 vccd1 vccd1 net7502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6989 _00500_ vssd1 vssd1 vccd1 vccd1 net7513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21264_ clknet_leaf_71_i_clk net4782 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold530 net5441 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 net5511 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold552 net7639 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20215_ net1491 _03731_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__or2_1
Xhold563 net5453 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold574 net7645 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
X_21195_ _02752_ net4621 net4439 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__a21bo_1
Xhold585 _01251_ vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 net6410 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20146_ net3684 _03692_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__or2_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20077_ net3700 net3636 _03580_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__mux2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 net6725 vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 net6677 vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 _01554_ vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1263 net6681 vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 net6685 vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 net6775 vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 _01495_ vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _05017_ _05018_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ net6580 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ net924 net1364 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ clknet_1_0__leaf__04800_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__buf_1
XFILLER_0_71_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ _06669_ _06634_ _06639_ _06670_ _06552_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a311o_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ net7091 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13451_ _06560_ _06593_ _06514_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__a21o_1
X_10663_ net5800 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12402_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _05263_ vssd1 vssd1 vccd1 vccd1 _05569_
+ sky130_fd_sc_hd__mux2_1
X_16170_ _09242_ _09244_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__nor2_1
X_13382_ _06472_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15121_ net4433 net4483 _08219_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__mux2_1
X_12333_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _05493_ vssd1 vssd1 vccd1 vccd1 _05501_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15052_ _08150_ _08142_ _08183_ _08176_ _08047_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12264_ net4306 _05377_ _05378_ net4338 vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _07151_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11215_ net6776 net6790 _04481_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12195_ _05359_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__nor2_1
X_19860_ _03479_ net2945 vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__or2_1
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__buf_1
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__clkbuf_4
X_18811_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.debug_overlay.vplaneY\[-7\] _05393_
+ _02765_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__o31a_1
X_11146_ net6570 net750 _04448_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19791_ net3088 _03442_ net1719 _03441_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11077_ net7028 net5985 _04415_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
X_15954_ _09014_ _09027_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__a21oi_1
X_18742_ net3893 _02740_ _02261_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14905_ _07999_ _08053_ _07995_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__mux2_1
X_18673_ _02676_ _02677_ _02678_ _02679_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _08917_ _08959_ vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__xnor2_1
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _08329_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__or2_1
X_14836_ _07356_ _07509_ _07498_ net7757 vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__o211a_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__04012_ _04012_ vssd1 vssd1 vccd1 vccd1 clknet_0__04012_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17555_ _10402_ _10432_ _10430_ vssd1 vssd1 vccd1 vccd1 _10554_ sky130_fd_sc_hd__a21oi_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14767_ _07882_ _07917_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__xnor2_2
X_11979_ _04604_ _05138_ _05137_ _04602_ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16506_ _09576_ _09577_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13718_ _06796_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__clkbuf_4
X_17486_ _10483_ _10484_ vssd1 vssd1 vccd1 vccd1 _10485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14698_ _07847_ _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20715__148 clknet_1_1__leaf__03985_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__inv_2
X_16437_ _09415_ _09416_ _09509_ vssd1 vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19225_ net5740 _03106_ _03113_ _03096_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__o211a_1
X_13649_ _06742_ _06713_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19156_ net5447 _03065_ _03071_ _03061_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__o211a_1
X_16368_ _09315_ _09316_ _09256_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__and3b_1
Xhold6208 net1947 vssd1 vssd1 vccd1 vccd1 net6732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6219 rbzero.tex_r0\[29\] vssd1 vssd1 vccd1 vccd1 net6743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18107_ _02152_ _02153_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__and2_1
X_15319_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19087_ net622 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
Xhold5507 net1861 vssd1 vssd1 vccd1 vccd1 net6031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ _09365_ _09372_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5518 rbzero.spi_registers.buf_texadd1\[23\] vssd1 vssd1 vccd1 vccd1 net6042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5529 _00947_ vssd1 vssd1 vccd1 vccd1 net6053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _01833_ _02025_ _02085_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4806 net915 vssd1 vssd1 vccd1 vccd1 net5330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4817 rbzero.spi_registers.texadd1\[4\] vssd1 vssd1 vccd1 vccd1 net5341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4828 rbzero.spi_registers.texadd0\[8\] vssd1 vssd1 vccd1 vccd1 net5352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4839 rbzero.spi_registers.texadd0\[23\] vssd1 vssd1 vccd1 vccd1 net5363 sky130_fd_sc_hd__dlygate4sd3_1
X_20000_ rbzero.debug_overlay.facingY\[-9\] net3756 _03594_ vssd1 vssd1 vccd1 vccd1
+ _03599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19989_ net3141 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21951_ net176 net2694 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ clknet_1_1__leaf__04000_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__buf_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21882_ clknet_leaf_99_i_clk net1163 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7421 _08623_ vssd1 vssd1 vccd1 vccd1 net7945 sky130_fd_sc_hd__dlygate4sd3_1
X_22434_ clknet_leaf_40_i_clk net4940 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6720 rbzero.tex_g0\[48\] vssd1 vssd1 vccd1 vccd1 net7244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__04001_ clknet_0__04001_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04001_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6731 net2717 vssd1 vssd1 vccd1 vccd1 net7255 sky130_fd_sc_hd__dlygate4sd3_1
X_22365_ net497 net2261 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold6742 net2702 vssd1 vssd1 vccd1 vccd1 net7266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6753 rbzero.tex_r1\[1\] vssd1 vssd1 vccd1 vccd1 net7277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6764 net2830 vssd1 vssd1 vccd1 vccd1 net7288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6775 rbzero.tex_r0\[4\] vssd1 vssd1 vccd1 vccd1 net7299 sky130_fd_sc_hd__dlygate4sd3_1
X_21316_ clknet_leaf_73_i_clk net4279 vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_22296_ net428 net2697 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold6786 rbzero.pov.ready_buffer\[69\] vssd1 vssd1 vccd1 vccd1 net7310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6797 _02931_ vssd1 vssd1 vccd1 vccd1 net7321 sky130_fd_sc_hd__dlygate4sd3_1
X_21247_ clknet_leaf_53_i_clk net3335 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold360 net5309 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 net5237 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 net5246 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _04332_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__clkbuf_4
Xhold393 net5164 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
X_21178_ net4201 _04140_ _04141_ _10329_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__a22o_1
X_20129_ net3817 _03676_ _03684_ _03683_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__o211a_1
X_20820__243 clknet_1_0__leaf__03995_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__inv_2
XFILLER_0_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _06105_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__and2_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 net4470 vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1071 net6244 vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__clkbuf_8
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _08722_ _08744_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__xnor2_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _00882_ vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 _00810_ vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _05997_ _06038_ _06039_ _06012_ _05999_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__a221o_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _07723_ _07724_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__xnor2_2
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__buf_4
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _10250_ _10338_ _10339_ vssd1 vssd1 vccd1 vccd1 _10340_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _07697_ _07700_ _07701_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__nand3_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ net869 net1529 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nand2_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__inv_2
X_17271_ _10269_ _10271_ vssd1 vssd1 vccd1 vccd1 _10272_ sky130_fd_sc_hd__nor2_1
X_10715_ net6880 net2085 _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _07586_ _07633_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11695_ net4033 net2905 vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nand2_1
X_19010_ net3885 _02976_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16222_ net7406 vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__buf_1
XFILLER_0_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _06541_ _06573_ _06561_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__o21a_1
X_10646_ net7008 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16153_ _08618_ _08665_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer5 _06966_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_1
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13365_ _04635_ _06497_ _06499_ _06503_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a2111o_1
X_15104_ _08218_ net3048 net6282 _08215_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__o211a_1
X_12316_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _05483_ vssd1 vssd1 vccd1 vccd1 _05484_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16084_ _09138_ _08874_ _09158_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13296_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19912_ _08333_ _03480_ _03529_ net2836 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__o211a_1
X_15035_ net7757 _08092_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__nand2_1
X_12247_ rbzero.debug_overlay.facingX\[-9\] _05382_ _05413_ _05415_ vssd1 vssd1 vccd1
+ vccd1 _05416_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19843_ net4335 _03475_ net734 _03454_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _05341_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__nor2_1
X_11129_ net7016 net6980 _04437_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19774_ net2070 _03429_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or2_1
X_16986_ _09988_ _09997_ vssd1 vssd1 vccd1 vccd1 _09998_ sky130_fd_sc_hd__xnor2_1
X_18725_ net6304 _02727_ _02714_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
X_20795__220 clknet_1_1__leaf__03993_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__inv_2
X_15937_ _09008_ _09007_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15868_ _08940_ _08942_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__nor2_4
X_18656_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _02637_
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_204_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17607_ _01657_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__and2b_1
X_14819_ _07691_ _07969_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15799_ _08514_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__clkbuf_4
X_21000__26 clknet_1_1__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
X_18587_ rbzero.wall_tracer.rayAddendX\[0\] _02599_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17538_ _10531_ _10536_ vssd1 vssd1 vccd1 vccd1 _10537_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17469_ _10353_ _10354_ _10351_ vssd1 vssd1 vccd1 vccd1 _10468_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19208_ _03088_ net3129 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20480_ _03858_ net3666 vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__and2_1
Xhold6005 net1516 vssd1 vssd1 vccd1 vccd1 net6529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6016 _04504_ vssd1 vssd1 vccd1 vccd1 net6540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6027 net1512 vssd1 vssd1 vccd1 vccd1 net6551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19139_ net5065 _03053_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__or2_1
Xhold6038 net1625 vssd1 vssd1 vccd1 vccd1 net6562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6049 rbzero.tex_g0\[47\] vssd1 vssd1 vccd1 vccd1 net6573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5304 net2472 vssd1 vssd1 vccd1 vccd1 net5828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5315 _00935_ vssd1 vssd1 vccd1 vccd1 net5839 sky130_fd_sc_hd__dlygate4sd3_1
X_22150_ net282 net2745 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
Xhold5326 net1833 vssd1 vssd1 vccd1 vccd1 net5850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5337 net2155 vssd1 vssd1 vccd1 vccd1 net5861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5348 net2464 vssd1 vssd1 vccd1 vccd1 net5872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4603 rbzero.spi_registers.texadd0\[6\] vssd1 vssd1 vccd1 vccd1 net5127 sky130_fd_sc_hd__dlygate4sd3_1
X_21101_ _04018_ _04091_ net4938 _04017_ net1886 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a32o_1
Xhold5359 net2467 vssd1 vssd1 vccd1 vccd1 net5883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4614 net926 vssd1 vssd1 vccd1 vccd1 net5138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4625 net897 vssd1 vssd1 vccd1 vccd1 net5149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22081_ clknet_leaf_79_i_clk _01250_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4636 rbzero.spi_registers.buf_texadd0\[19\] vssd1 vssd1 vccd1 vccd1 net5160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3902 _01636_ vssd1 vssd1 vccd1 vccd1 net4426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4647 rbzero.spi_registers.texadd0\[10\] vssd1 vssd1 vccd1 vccd1 net5171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4658 net958 vssd1 vssd1 vccd1 vccd1 net5182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3913 net3179 vssd1 vssd1 vccd1 vccd1 net4437 sky130_fd_sc_hd__buf_1
Xhold3924 _01009_ vssd1 vssd1 vccd1 vccd1 net4448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4669 net1290 vssd1 vssd1 vccd1 vccd1 net5193 sky130_fd_sc_hd__dlygate4sd3_1
X_21032_ net5379 net5168 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nor2_1
Xhold3935 rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 net4459 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3946 _01604_ vssd1 vssd1 vccd1 vccd1 net4470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3957 net1077 vssd1 vssd1 vccd1 vccd1 net4481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20290__27 clknet_1_1__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
Xhold3968 rbzero.debug_overlay.vplaneX\[-6\] vssd1 vssd1 vccd1 vccd1 net4492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3979 net1166 vssd1 vssd1 vccd1 vccd1 net4503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21934_ clknet_leaf_9_i_clk net1200 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ clknet_leaf_94_i_clk net3564 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21796_ clknet_leaf_12_i_clk net2815 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11480_ rbzero.texu_hot\[4\] _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7240 _08487_ vssd1 vssd1 vccd1 vccd1 net7764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22417_ net145 net2688 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7251 _08406_ vssd1 vssd1 vccd1 vccd1 net7775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7273 rbzero.wall_tracer.stepDistX\[6\] vssd1 vssd1 vccd1 vccd1 net7797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6550 rbzero.tex_g1\[49\] vssd1 vssd1 vccd1 vccd1 net7074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7295 rbzero.wall_tracer.stepDistY\[-5\] vssd1 vssd1 vccd1 vccd1 net7819 sky130_fd_sc_hd__dlygate4sd3_1
X_13150_ net3472 _06301_ net3321 _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__a2bb2o_1
X_22348_ net480 net1474 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
Xhold6561 net2458 vssd1 vssd1 vccd1 vccd1 net7085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6572 rbzero.tex_b1\[38\] vssd1 vssd1 vccd1 vccd1 net7096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6583 net2587 vssd1 vssd1 vccd1 vccd1 net7107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6594 rbzero.tex_b1\[58\] vssd1 vssd1 vccd1 vccd1 net7118 sky130_fd_sc_hd__dlygate4sd3_1
X_12101_ _05261_ _05269_ _05034_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__o21a_1
Xhold5860 _04399_ vssd1 vssd1 vccd1 vccd1 net6384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5871 net1148 vssd1 vssd1 vccd1 vccd1 net6395 sky130_fd_sc_hd__dlygate4sd3_1
X_13081_ _06231_ _06234_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__or3_1
X_22279_ net411 net2336 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
X_20656__95 clknet_1_1__leaf__03781_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__inv_2
Xhold5882 rbzero.tex_r0\[34\] vssd1 vssd1 vccd1 vccd1 net6406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5893 net1202 vssd1 vssd1 vccd1 vccd1 net6417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ _04816_ _05198_ net4043 _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a211oi_1
Xhold190 net4516 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _09297_ net4106 vssd1 vssd1 vccd1 vccd1 _09910_ sky130_fd_sc_hd__xor2_1
X_16771_ _08872_ _08582_ vssd1 vssd1 vccd1 vccd1 _09841_ sky130_fd_sc_hd__nor2_1
X_13983_ _07127_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15722_ _08699_ _08700_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18510_ _09932_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__clkbuf_4
X_12934_ net4078 _06057_ _06065_ _06060_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__or4bb_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ net6275 _03266_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _08725_ _08726_ _08727_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _02467_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__clkbuf_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ net30 _06003_ _06022_ net32 vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__a22o_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14604_ _07474_ _07304_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ net3026 _04970_ _04985_ _04952_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__o211ai_4
X_18372_ net4538 net4405 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _08642_ _08602_ _08658_ _08645_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__a22o_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ net23 vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _10213_ _10214_ _10323_ vssd1 vssd1 vccd1 vccd1 _10324_ sky130_fd_sc_hd__a21oi_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _07649_ _07667_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__or2b_1
X_11747_ net2931 _04915_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a21boi_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17254_ _10154_ _10159_ vssd1 vssd1 vccd1 vccd1 _10255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03992_ _03992_ vssd1 vssd1 vccd1 vccd1 clknet_0__03992_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14466_ _07604_ _07610_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__xor2_4
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11678_ net3008 net4049 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16205_ _09278_ _09279_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13417_ net7440 _06431_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nor2_1
X_17185_ _09885_ _09887_ vssd1 vssd1 vccd1 vccd1 _10187_ sky130_fd_sc_hd__and2_2
X_10629_ net2751 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__clkbuf_1
X_14397_ _07517_ _07547_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__nand2_1
X_16136_ _09209_ _09210_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13348_ _06430_ _06171_ _06498_ _04635_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_45_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20827__249 clknet_1_0__leaf__03996_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__inv_2
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _09140_ _09141_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__clkbuf_4
Xhold3209 _03922_ vssd1 vssd1 vccd1 vccd1 net3733 sky130_fd_sc_hd__dlygate4sd3_1
X_15018_ net4423 _08155_ _08138_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2508 _03491_ vssd1 vssd1 vccd1 vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2519 rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 net3043 sky130_fd_sc_hd__dlymetal6s2s_1
X_19826_ net55 _03026_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__and2_1
Xhold1807 net6837 vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1818 _01279_ vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1829 net5863 vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
X_19757_ _03426_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16969_ net2787 _09968_ _09982_ vssd1 vssd1 vccd1 vccd1 _09983_ sky130_fd_sc_hd__a21oi_1
X_18708_ _02705_ _02706_ _02711_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19688_ net6104 _03374_ net1769 _03384_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _02647_ rbzero.wall_tracer.rayAddendX\[3\] _02643_ vssd1 vssd1 vccd1 vccd1
+ _02648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21650_ clknet_leaf_33_i_clk net5786 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20601_ _03945_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__clkbuf_1
X_21581_ clknet_leaf_2_i_clk net893 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20532_ net3802 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20463_ net3764 net1278 _03845_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22202_ net334 net1767 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
Xhold5101 rbzero.pov.spi_buffer\[37\] vssd1 vssd1 vccd1 vccd1 net5625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5112 rbzero.pov.spi_buffer\[52\] vssd1 vssd1 vccd1 vccd1 net5636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20394_ _03791_ net3318 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and2_1
Xhold5123 _01074_ vssd1 vssd1 vccd1 vccd1 net5647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5134 net1327 vssd1 vssd1 vccd1 vccd1 net5658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5145 net1350 vssd1 vssd1 vccd1 vccd1 net5669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4400 net1250 vssd1 vssd1 vccd1 vccd1 net4924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4411 rbzero.traced_texa\[3\] vssd1 vssd1 vccd1 vccd1 net4935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22133_ net265 net1236 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
Xhold5156 rbzero.spi_registers.texadd0\[19\] vssd1 vssd1 vccd1 vccd1 net5680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5167 _00786_ vssd1 vssd1 vccd1 vccd1 net5691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4422 _01587_ vssd1 vssd1 vccd1 vccd1 net4946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5178 net1402 vssd1 vssd1 vccd1 vccd1 net5702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4433 _01644_ vssd1 vssd1 vccd1 vccd1 net4957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4444 net690 vssd1 vssd1 vccd1 vccd1 net4968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5189 rbzero.spi_registers.texadd1\[22\] vssd1 vssd1 vccd1 vccd1 net5713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3710 net840 vssd1 vssd1 vccd1 vccd1 net4234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4455 net775 vssd1 vssd1 vccd1 vccd1 net4979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4466 rbzero.spi_registers.buf_texadd0\[17\] vssd1 vssd1 vccd1 vccd1 net4990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3721 _00765_ vssd1 vssd1 vccd1 vccd1 net4245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3732 net1496 vssd1 vssd1 vccd1 vccd1 net4256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22064_ clknet_leaf_7_i_clk net3486 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4477 net804 vssd1 vssd1 vccd1 vccd1 net5001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4488 _00868_ vssd1 vssd1 vccd1 vccd1 net5012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3743 rbzero.spi_registers.texadd2\[10\] vssd1 vssd1 vccd1 vccd1 net4267 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03981_ clknet_0__03981_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03981_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3754 net1673 vssd1 vssd1 vccd1 vccd1 net4278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4499 _00737_ vssd1 vssd1 vccd1 vccd1 net5023 sky130_fd_sc_hd__dlygate4sd3_1
X_21015_ net839 net4975 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__nand2_1
Xhold3765 _00978_ vssd1 vssd1 vccd1 vccd1 net4289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3776 net7427 vssd1 vssd1 vccd1 vccd1 net4300 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3787 _08049_ vssd1 vssd1 vccd1 vccd1 net4311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3798 net4318 vssd1 vssd1 vccd1 vccd1 net4322 sky130_fd_sc_hd__clkbuf_2
X_10980_ net1771 net6415 _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
X_21917_ clknet_leaf_92_i_clk net1344 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ net41 _05795_ _05799_ _05207_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20932__344 clknet_1_1__leaf__04006_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__inv_2
X_21848_ clknet_leaf_83_i_clk net1441 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ rbzero.spi_registers.texadd1\[1\] _04644_ _04709_ vssd1 vssd1 vccd1 vccd1
+ _04773_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12581_ _05744_ _05745_ _05261_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21779_ clknet_leaf_20_i_clk net6035 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _07366_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11532_ rbzero.spi_registers.texadd0\[22\] _04680_ _04703_ vssd1 vssd1 vccd1 vccd1
+ _04704_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14251_ _07356_ _07354_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7070 rbzero.wall_tracer.stepDistX\[-5\] vssd1 vssd1 vccd1 vccd1 net7594 sky130_fd_sc_hd__dlygate4sd3_1
X_13202_ _06349_ _06351_ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14182_ _07326_ _07327_ _07331_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nor3_1
Xhold7092 rbzero.wall_tracer.rayAddendY\[-8\] vssd1 vssd1 vccd1 vccd1 net7616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11394_ net7139 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
Xhold6380 net2334 vssd1 vssd1 vccd1 vccd1 net6904 sky130_fd_sc_hd__dlygate4sd3_1
X_13133_ net3500 _06277_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and2_1
Xhold6391 rbzero.tex_g1\[62\] vssd1 vssd1 vccd1 vccd1 net6915 sky130_fd_sc_hd__dlygate4sd3_1
X_18990_ net6141 net3265 net4902 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5690 _00982_ vssd1 vssd1 vccd1 vccd1 net6214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17941_ _10379_ _09418_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__nor2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _04895_ _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12015_ net1326 _05022_ _05027_ net1402 _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17872_ _10520_ _10407_ _10416_ _01684_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_206_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19611_ net3022 _03340_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or2_1
X_16823_ _09850_ _09891_ _09892_ vssd1 vssd1 vccd1 vccd1 _09893_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19542_ net3866 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__clkbuf_1
X_16754_ _09822_ _09823_ vssd1 vssd1 vccd1 vccd1 _09824_ sky130_fd_sc_hd__nor2_1
X_13966_ _07114_ _07115_ _07116_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15705_ _08773_ _08769_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__or2b_1
X_12917_ net46 _06066_ _06073_ _06057_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a211o_1
X_16685_ _09754_ _09755_ vssd1 vssd1 vccd1 vccd1 _09756_ sky130_fd_sc_hd__and2b_1
X_19473_ net3123 net2951 net3077 vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__mux2_1
X_13897_ _06861_ net79 _06923_ _06844_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ net4573 net4386 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__nor2_1
X_15636_ _08410_ _08470_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ net33 _06005_ net29 net30 vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and4b_1
XFILLER_0_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15567_ _08641_ _08541_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18355_ net4453 net3505 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__nand2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _05933_ _05934_ _05936_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a211o_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17306_ _10292_ _10306_ vssd1 vssd1 vccd1 vccd1 _10307_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14518_ _07617_ _07628_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__xnor2_4
X_15498_ _08533_ _08572_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18286_ _02266_ _02267_ _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17237_ _09813_ _10236_ _10237_ vssd1 vssd1 vccd1 vccd1 _10238_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14449_ _07529_ _07530_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold904 net6513 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ net4954 _08664_ _09870_ _10169_ vssd1 vssd1 vccd1 vccd1 _10170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold915 _01064_ vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _01538_ vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold937 net6505 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ _08529_ _08470_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__nor2_1
Xhold948 net2100 vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17099_ _09795_ _09796_ _09798_ vssd1 vssd1 vccd1 vccd1 _10101_ sky130_fd_sc_hd__o21a_1
Xhold959 net3811 vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3006 net1413 vssd1 vssd1 vccd1 vccd1 net3530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3017 _00414_ vssd1 vssd1 vccd1 vccd1 net3541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3028 _02672_ vssd1 vssd1 vccd1 vccd1 net3552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3039 net7331 vssd1 vssd1 vccd1 vccd1 net3563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2305 _01541_ vssd1 vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2316 net5974 vssd1 vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2327 net7261 vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 net7305 vssd1 vssd1 vccd1 vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1604 net7082 vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2349 net7666 vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 _01573_ vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1626 net6765 vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
X_19809_ net6051 _03428_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__or2_1
Xhold1637 net7039 vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 rbzero.tex_b1\[39\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1659 net5963 vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21702_ clknet_leaf_101_i_clk net862 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21633_ clknet_leaf_28_i_clk net3257 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21564_ clknet_leaf_26_i_clk net5479 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20515_ _03880_ net3612 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__and2_1
X_21495_ clknet_leaf_15_i_clk net2824 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20446_ net3845 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20377_ _03791_ net3738 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4230 _02644_ vssd1 vssd1 vccd1 vccd1 net4754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22116_ net248 net1840 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold4241 net980 vssd1 vssd1 vccd1 vccd1 net4765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4252 net2833 vssd1 vssd1 vccd1 vccd1 net4776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4263 net3006 vssd1 vssd1 vccd1 vccd1 net4787 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold4274 _01030_ vssd1 vssd1 vccd1 vccd1 net4798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3540 _04845_ vssd1 vssd1 vccd1 vccd1 net4064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3551 _09923_ vssd1 vssd1 vccd1 vccd1 net4075 sky130_fd_sc_hd__dlygate4sd3_1
X_22047_ clknet_leaf_91_i_clk net3308 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold4296 net3092 vssd1 vssd1 vccd1 vccd1 net4820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3562 net3480 vssd1 vssd1 vccd1 vccd1 net4086 sky130_fd_sc_hd__buf_2
Xhold3573 _00457_ vssd1 vssd1 vccd1 vccd1 net4097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3584 rbzero.row_render.size\[10\] vssd1 vssd1 vccd1 vccd1 net4108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2850 net3968 vssd1 vssd1 vccd1 vccd1 net3374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3595 _00789_ vssd1 vssd1 vccd1 vccd1 net4119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2861 _03938_ vssd1 vssd1 vccd1 vccd1 net3385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2872 _02408_ vssd1 vssd1 vccd1 vccd1 net3396 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2883 net4693 vssd1 vssd1 vccd1 vccd1 net3407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13820_ _06970_ net529 vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__or2_1
Xhold2894 net7475 vssd1 vssd1 vccd1 vccd1 net3418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ _06892_ net576 vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963_ net6836 net6982 _04355_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12702_ net43 _05844_ _05852_ net46 vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a22o_1
X_16470_ _09539_ _09541_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13682_ _06567_ _06565_ _06688_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__mux2_1
X_10894_ _04169_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _06210_ _08381_ _08479_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__or3_1
X_12633_ net4 net5 vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18140_ _02184_ _02185_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__or2_1
X_15352_ _06163_ _06510_ _08300_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__mux2_1
X_12564_ rbzero.tex_b1\[47\] rbzero.tex_b1\[46\] _04988_ vssd1 vssd1 vccd1 vccd1 _05729_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ _07447_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18071_ _10379_ _09536_ _02117_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__o21ai_1
X_11515_ _04645_ _04683_ _04684_ _04685_ _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15283_ _08356_ _08357_ _06177_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__mux2_1
X_12495_ _05279_ _05658_ _05660_ _05461_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17022_ _10030_ net4597 _09966_ vssd1 vssd1 vccd1 vccd1 _10031_ sky130_fd_sc_hd__mux2_1
X_14234_ _07373_ _07384_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__xnor2_1
X_11446_ net4104 net89 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__nand2_2
XFILLER_0_22_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14165_ _06737_ net545 _06973_ _06931_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__o22a_1
X_11377_ net7048 net6351 _04573_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13116_ net3851 vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__inv_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _07198_ _07226_ _07246_ _07239_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__a2bb2o_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _09952_ _09953_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _01973_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__clkbuf_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ net3507 net4910 vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__or2_1
X_17855_ _01889_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16806_ _09871_ _09872_ _09874_ vssd1 vssd1 vccd1 vccd1 _09876_ sky130_fd_sc_hd__a21o_1
X_17786_ _01832_ _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nand2_1
X_14998_ net4405 _08137_ _08138_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19525_ net1572 _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__or2_1
X_16737_ _09804_ _09806_ vssd1 vssd1 vccd1 vccd1 _09807_ sky130_fd_sc_hd__xor2_1
X_13949_ _07079_ _07073_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19456_ net3182 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__clkbuf_1
X_16668_ net3722 _09304_ _09486_ _09738_ vssd1 vssd1 vccd1 vccd1 _09739_ sky130_fd_sc_hd__or4_4
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18407_ _02437_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15619_ _08687_ _08693_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__xor2_1
XFILLER_0_186_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19387_ net5629 _03198_ _03205_ _03194_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__o211a_1
X_16599_ _09541_ _09668_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18338_ net4491 net4473 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18269_ _02295_ _02314_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20300_ clknet_1_1__leaf__03773_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21280_ clknet_leaf_59_i_clk _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold701 net5531 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 _01302_ vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 net3487 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
X_20231_ net3275 _03730_ _03741_ _03735_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__o211a_1
Xhold734 net6436 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _01322_ vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold756 net5590 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold767 net5194 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20961__370 clknet_1_1__leaf__04009_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__inv_2
X_20162_ net5540 _03691_ _03702_ _03696_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__o211a_1
Xhold778 net4880 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold789 net5679 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2102 _04320_ vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2113 _01553_ vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
X_20093_ net2629 net4796 vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__nor2_1
Xhold2124 _04172_ vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2135 net7098 vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1401 _01307_ vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2146 _01489_ vssd1 vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2157 _01516_ vssd1 vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 net6967 vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 net6731 vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 net7218 vssd1 vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 _04222_ vssd1 vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _01364_ vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1445 _01167_ vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1456 _04382_ vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1467 _00937_ vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 net5855 vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1489 rbzero.spi_registers.buf_texadd3\[11\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21616_ clknet_leaf_25_i_clk net5607 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21547_ clknet_leaf_17_i_clk net848 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11300_ net5819 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
X_12280_ net4532 _05111_ _05095_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21478_ clknet_leaf_102_i_clk net2972 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ net2198 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
X_20429_ _03814_ net3353 vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11162_ net5816 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4060 net3168 vssd1 vssd1 vccd1 vccd1 net4584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4071 net3047 vssd1 vssd1 vccd1 vccd1 net4595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4082 rbzero.spi_registers.buf_texadd0\[20\] vssd1 vssd1 vccd1 vccd1 net4606 sky130_fd_sc_hd__dlygate4sd3_1
X_15970_ _08962_ _08755_ _09020_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__a21bo_1
X_11093_ _04403_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__clkbuf_4
Xhold4093 net1588 vssd1 vssd1 vccd1 vccd1 net4617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3370 _02741_ vssd1 vssd1 vccd1 vccd1 net3894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3381 _02977_ vssd1 vssd1 vccd1 vccd1 net3905 sky130_fd_sc_hd__dlygate4sd3_1
X_14921_ net7771 vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__buf_4
Xhold3392 _00623_ vssd1 vssd1 vccd1 vccd1 net3916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2680 net6079 vssd1 vssd1 vccd1 vccd1 net3204 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _01682_ _01691_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nand2_1
Xhold72 net4292 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2691 _00574_ vssd1 vssd1 vccd1 vccd1 net3215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 _03131_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net7438 _08002_ _06707_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 net3010 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1990 net6957 vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _06880_ _06953_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__nand2_1
X_17571_ _06204_ _10569_ vssd1 vssd1 vccd1 vccd1 _10570_ sky130_fd_sc_hd__nand2_1
X_14783_ _07922_ _07932_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11995_ _05122_ net3987 net2986 _05163_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a221o_1
X_19310_ net5182 _03159_ _03162_ _03155_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__o211a_1
X_16522_ _09593_ _09477_ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__nor2_1
X_13734_ _06806_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10946_ net5897 net6890 _04344_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19241_ net5201 _03120_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__or2_1
X_16453_ _09524_ _09525_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__nor2_1
X_13665_ _06669_ _06687_ _06757_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__o21a_1
X_10877_ net2164 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _05780_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_15404_ net4105 net3028 _08439_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__or3_4
X_16384_ _08394_ _08717_ _09336_ _09334_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__o31a_1
X_19172_ net2590 _03079_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13596_ _06697_ _06698_ _06591_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a21o_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15335_ net3216 _06210_ _08409_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18123_ _02166_ _02169_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__o21a_1
X_12547_ _05710_ _05711_ _05177_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18054_ _01812_ _10416_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__nor2_1
X_15266_ _06535_ _08336_ net7403 _08340_ _06570_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__a41o_2
X_12478_ _05261_ _05641_ _05643_ _05461_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_3 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17005_ net4528 net4727 vssd1 vssd1 vccd1 vccd1 _10015_ sky130_fd_sc_hd__nor2_1
X_14217_ _06737_ _07366_ _07367_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11429_ _04604_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ net4046 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _07297_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14079_ _07191_ _07227_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__and3b_1
X_18956_ _02924_ _02928_ _02937_ _04624_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__a211o_1
X_17907_ _01955_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__and2b_1
XFILLER_0_207_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18887_ _02872_ _02873_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__or2_1
XFILLER_0_206_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17838_ _09562_ net7378 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer15 net538 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 _07109_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_1
XFILLER_0_179_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer37 _06781_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_1
X_17769_ _01706_ _01800_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a21o_1
Xrebuffer48 _06893_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_1
Xrebuffer59 _07106_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19508_ _03141_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__clkbuf_4
X_20780_ clknet_1_0__leaf__03989_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__buf_1
XFILLER_0_147_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19439_ net2230 _03225_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22450_ clknet_leaf_66_i_clk _01619_ vssd1 vssd1 vccd1 vccd1 reg_gpout\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21401_ clknet_leaf_65_i_clk _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22381_ net513 net2558 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6913 _08130_ vssd1 vssd1 vccd1 vccd1 net7437 sky130_fd_sc_hd__buf_1
Xhold6924 rbzero.traced_texVinit\[8\] vssd1 vssd1 vccd1 vccd1 net7448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6935 rbzero.wall_tracer.trackDistY\[-11\] vssd1 vssd1 vccd1 vccd1 net7459 sky130_fd_sc_hd__dlygate4sd3_1
X_21332_ clknet_leaf_55_i_clk net4299 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6957 rbzero.wall_tracer.trackDistY\[5\] vssd1 vssd1 vccd1 vccd1 net7481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6968 net4139 vssd1 vssd1 vccd1 vccd1 net7492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold520 net5436 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
X_21263_ clknet_leaf_71_i_clk net3635 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold531 net5443 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 net5394 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold553 net4480 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
X_20214_ net5439 _03730_ _03732_ _03722_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold564 net6374 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21194_ _02529_ net4439 _04149_ _02528_ net723 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a32o_1
Xhold575 net4414 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold586 net6382 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold597 net6412 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20145_ net3684 _03691_ _03693_ _03683_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ net3428 _03577_ net4460 _03636_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__o211a_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 net6262 vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 _01154_ vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 net6679 vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 net6631 vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1264 _03398_ vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _01385_ vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _04491_ vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 net6835 vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ net6578 net2307 _04266_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__mux2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _04948_ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ net7089 net2382 _04225_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13450_ net4947 _06505_ _06508_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__o21ai_4
X_10662_ net5798 net1762 _04192_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _05550_ _05567_ _05028_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ _06473_ _06435_ _06474_ _06475_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _08218_ _08231_ net3223 _08215_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__o211a_1
X_12332_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _05070_ vssd1 vssd1 vccd1 vccd1 _05500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20296__33 clknet_1_0__leaf__03774_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
X_15051_ _08164_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__inv_2
X_12263_ net3028 _05374_ _05372_ net3821 vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _07108_ net550 _07152_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__a21oi_2
X_11214_ net2228 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12194_ _05357_ _05360_ _05346_ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__and4b_1
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 o_gpout[4] sky130_fd_sc_hd__buf_1
X_18810_ net4626 _02798_ _02797_ _02792_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a211o_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__clkbuf_4
X_11145_ net2350 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
X_19790_ net6650 _03443_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18741_ _06193_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__xnor2_1
X_11076_ net6612 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
X_15953_ _09015_ _09016_ _09026_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__and3_1
XFILLER_0_208_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14904_ _08008_ _08010_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__nor2_1
X_18672_ _02646_ net3242 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__nand2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ net3539 _08311_ _08379_ _08391_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__or4_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _08596_ _08597_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__nand2_2
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14835_ _07584_ _07978_ _07984_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__o31ai_4
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04011_ _04011_ vssd1 vssd1 vccd1 vccd1 clknet_0__04011_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _10529_ _10552_ vssd1 vssd1 vccd1 vccd1 _10553_ sky130_fd_sc_hd__xnor2_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14766_ _07877_ _07884_ _07916_ _07880_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__and4_1
X_11978_ _05141_ _05147_ _05138_ _04604_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16505_ _09574_ _09575_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10929_ net2830 net6752 _04333_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
X_13717_ _06862_ _06865_ _06858_ _06867_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__or4_4
X_17485_ _09051_ _09784_ vssd1 vssd1 vccd1 vccd1 _10484_ sky130_fd_sc_hd__nor2_1
X_14697_ _07444_ _07590_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19224_ net5087 _03107_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__or2_1
X_16436_ _09442_ _09508_ vssd1 vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13648_ _06752_ _06741_ _06797_ _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19155_ net5283 _03066_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__or2_1
X_16367_ _09438_ _09439_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__or2b_1
X_13579_ _06697_ _06698_ _06616_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__a21o_1
Xhold6209 _04582_ vssd1 vssd1 vccd1 vccd1 net6733 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_53_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18106_ _02152_ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15318_ net3149 _06210_ _08391_ _08392_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_48_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16298_ _09369_ _09370_ _09227_ _09371_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__o2bb2a_1
X_19086_ net6324 _03026_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5508 rbzero.spi_registers.spi_buffer\[23\] vssd1 vssd1 vccd1 vccd1 net6032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5519 net1548 vssd1 vssd1 vccd1 vccd1 net6043 sky130_fd_sc_hd__dlygate4sd3_1
X_18037_ _01836_ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ net4315 _08299_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__nor2_1
Xhold4807 _00694_ vssd1 vssd1 vccd1 vccd1 net5331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4818 net966 vssd1 vssd1 vccd1 vccd1 net5342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4829 net1004 vssd1 vssd1 vccd1 vccd1 net5353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_160_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19988_ _03261_ net3140 vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18939_ _02903_ _02909_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21950_ net175 net730 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21881_ clknet_leaf_99_i_clk net1169 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7400 rbzero.wall_tracer.stepDistX\[5\] vssd1 vssd1 vccd1 vccd1 net7924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22433_ clknet_leaf_40_i_clk net4703 vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6710 rbzero.tex_r0\[7\] vssd1 vssd1 vccd1 vccd1 net7234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22364_ net496 net2701 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold6721 net2662 vssd1 vssd1 vccd1 vccd1 net7245 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__04000_ clknet_0__04000_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04000_
+ sky130_fd_sc_hd__clkbuf_16
Xhold6732 rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1 net7256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6743 rbzero.tex_b1\[10\] vssd1 vssd1 vccd1 vccd1 net7267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6754 net2753 vssd1 vssd1 vccd1 vccd1 net7278 sky130_fd_sc_hd__dlygate4sd3_1
X_21315_ clknet_leaf_73_i_clk _00484_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6765 rbzero.tex_r0\[35\] vssd1 vssd1 vccd1 vccd1 net7289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6776 net2714 vssd1 vssd1 vccd1 vccd1 net7300 sky130_fd_sc_hd__dlygate4sd3_1
X_22295_ net427 net2684 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6787 rbzero.spi_registers.spi_cmd\[1\] vssd1 vssd1 vccd1 vccd1 net7311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6798 net7363 vssd1 vssd1 vccd1 vccd1 net7322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21246_ clknet_leaf_55_i_clk net3792 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold350 net5127 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 net5311 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 net5146 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 net5248 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 net5166 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
X_21177_ net4185 _04140_ _04141_ _10205_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__a22o_1
X_20128_ net3590 _03679_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__or2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ net5696 _03613_ _03635_ _03636_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__o211a_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 net6054 vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__buf_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 net5713 vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 net6246 vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 net3948 vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ net6341 _05997_ _06037_ net56 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__a22o_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 net5749 vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11832_ _04992_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__clkbuf_8
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _07749_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14551_ _07697_ _07700_ _07701_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11763_ _04928_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__xnor2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _04169_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__clkbuf_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _06544_ _06645_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17270_ _10141_ _10142_ _10270_ vssd1 vssd1 vccd1 vccd1 _10271_ sky130_fd_sc_hd__a21boi_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _07615_ _07631_ _07632_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11694_ net4033 net2905 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13433_ _06582_ _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__xor2_2
X_16221_ _09295_ _06396_ net4088 vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__mux2_1
X_10645_ net7006 net2405 _04181_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ net3722 _08328_ _08628_ _09226_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__or4_4
X_13364_ _04635_ _06505_ _06508_ _06514_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__o211ai_4
Xrebuffer6 net529 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_1
XFILLER_0_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12315_ _04987_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__buf_4
X_15103_ net6281 _08201_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__or2_1
X_16083_ _09152_ _09153_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19911_ net2835 _03480_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nand2_1
X_15034_ net5686 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
X_12246_ rbzero.debug_overlay.facingX\[-3\] _05373_ _05379_ rbzero.debug_overlay.facingX\[-7\]
+ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19842_ net733 _03477_ _03479_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a211o_1
X_12177_ _05343_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ net6393 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
X_19773_ net3112 _03427_ net1965 _03424_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__o211a_1
X_16985_ _09995_ _09996_ vssd1 vssd1 vccd1 vccd1 _09997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ _04624_ _02725_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a21o_1
X_11059_ net2539 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
X_15936_ _08987_ _08981_ _08986_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__06092_ _06092_ vssd1 vssd1 vccd1 vccd1 clknet_0__06092_ sky130_fd_sc_hd__clkbuf_16
X_18655_ _02643_ _02645_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__and2_1
X_15867_ _08886_ _08889_ _08941_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__o21a_1
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _10509_ _10510_ _10512_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14818_ _07740_ _07741_ _07690_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _02593_ _02598_ _04623_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_130 vssd1 vssd1 vccd1 vccd1 ones[6] top_ew_algofoogle_130/LO sky130_fd_sc_hd__conb_1
X_15798_ _08516_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__buf_4
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _10534_ _10535_ vssd1 vssd1 vccd1 vccd1 _10536_ sky130_fd_sc_hd__xor2_1
X_14749_ _07892_ _07898_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _10374_ _10343_ vssd1 vssd1 vccd1 vccd1 _10467_ sky130_fd_sc_hd__or2b_1
XFILLER_0_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19207_ net3116 net3128 _03038_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__mux2_1
X_16419_ _09485_ _09491_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__xor2_2
XFILLER_0_156_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17399_ _10377_ _10290_ _10398_ vssd1 vssd1 vccd1 vccd1 _10399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6006 rbzero.tex_r0\[10\] vssd1 vssd1 vccd1 vccd1 net6530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6017 net1436 vssd1 vssd1 vccd1 vccd1 net6541 sky130_fd_sc_hd__dlygate4sd3_1
X_19138_ net5559 _03052_ _03060_ _03061_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__o211a_1
Xhold6028 _04348_ vssd1 vssd1 vccd1 vccd1 net6552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6039 rbzero.tex_r1\[45\] vssd1 vssd1 vccd1 vccd1 net6563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5305 _04177_ vssd1 vssd1 vccd1 vccd1 net5829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5316 net649 vssd1 vssd1 vccd1 vccd1 net5840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5327 rbzero.spi_registers.vshift\[3\] vssd1 vssd1 vccd1 vccd1 net5851 sky130_fd_sc_hd__dlygate4sd3_1
X_19069_ net6029 net2843 _03018_ _03011_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5338 _03227_ vssd1 vssd1 vccd1 vccd1 net5862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5349 _04496_ vssd1 vssd1 vccd1 vccd1 net5873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4604 net874 vssd1 vssd1 vccd1 vccd1 net5128 sky130_fd_sc_hd__dlygate4sd3_1
X_21100_ _04087_ net4937 _04089_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4615 rbzero.spi_registers.buf_texadd0\[18\] vssd1 vssd1 vccd1 vccd1 net5139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4626 rbzero.color_floor\[4\] vssd1 vssd1 vccd1 vccd1 net5150 sky130_fd_sc_hd__dlygate4sd3_1
X_22080_ clknet_leaf_6_i_clk net6178 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4637 net835 vssd1 vssd1 vccd1 vccd1 net5161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3903 net702 vssd1 vssd1 vccd1 vccd1 net4427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4648 net847 vssd1 vssd1 vccd1 vccd1 net5172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3914 rbzero.debug_overlay.vplaneY\[-9\] vssd1 vssd1 vccd1 vccd1 net4438 sky130_fd_sc_hd__buf_2
Xhold4659 _00742_ vssd1 vssd1 vccd1 vccd1 net5183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21031_ _04028_ _04029_ _04030_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold3925 net1299 vssd1 vssd1 vccd1 vccd1 net4449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_201_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20804__228 clknet_1_1__leaf__03994_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__inv_2
Xhold3936 _03646_ vssd1 vssd1 vccd1 vccd1 net4460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3947 net1584 vssd1 vssd1 vccd1 vccd1 net4471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3958 net7481 vssd1 vssd1 vccd1 vccd1 net4482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3969 net4476 vssd1 vssd1 vccd1 vccd1 net4493 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21933_ clknet_leaf_8_i_clk net1242 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ clknet_leaf_94_i_clk net3828 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21795_ clknet_leaf_12_i_clk net6157 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20746_ clknet_1_0__leaf__03780_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7230 net4518 vssd1 vssd1 vccd1 vccd1 net7754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22416_ net144 net2649 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7263 rbzero.wall_tracer.stepDistY\[6\] vssd1 vssd1 vccd1 vccd1 net7787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7274 _01977_ vssd1 vssd1 vccd1 vccd1 net7798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6540 net2439 vssd1 vssd1 vccd1 vccd1 net7064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold7285 _08368_ vssd1 vssd1 vccd1 vccd1 net7809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6551 net2246 vssd1 vssd1 vccd1 vccd1 net7075 sky130_fd_sc_hd__dlygate4sd3_1
X_22347_ net479 net2681 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
Xhold7296 net4472 vssd1 vssd1 vccd1 vccd1 net7820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6562 rbzero.tex_b0\[62\] vssd1 vssd1 vccd1 vccd1 net7086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6573 net2596 vssd1 vssd1 vccd1 vccd1 net7097 sky130_fd_sc_hd__dlygate4sd3_1
X_12100_ rbzero.tex_r1\[3\] rbzero.tex_r1\[2\] _05263_ vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6584 rbzero.tex_g1\[21\] vssd1 vssd1 vccd1 vccd1 net7108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5850 rbzero.tex_b1\[16\] vssd1 vssd1 vccd1 vccd1 net6374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6595 net2212 vssd1 vssd1 vccd1 vccd1 net7119 sky130_fd_sc_hd__dlygate4sd3_1
X_13080_ net3996 _06216_ net4821 _04827_ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22278_ net410 net1556 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
Xhold5861 net1111 vssd1 vssd1 vccd1 vccd1 net6385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5872 _04256_ vssd1 vssd1 vccd1 vccd1 net6396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5883 net1153 vssd1 vssd1 vccd1 vccd1 net6407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5894 rbzero.tex_r1\[30\] vssd1 vssd1 vccd1 vccd1 net6418 sky130_fd_sc_hd__dlygate4sd3_1
X_12031_ net6041 _05200_ net6220 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a21o_4
Xhold180 net5031 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
X_21229_ clknet_leaf_51_i_clk _00398_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold191 net7614 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
X_20744__175 clknet_1_0__leaf__03987_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__inv_2
X_16770_ _08684_ _09216_ vssd1 vssd1 vccd1 vccd1 _09840_ sky130_fd_sc_hd__nor2_1
X_13982_ _07127_ _07128_ _07132_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__nand3_1
X_15721_ _08325_ _08795_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__or2_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _06076_ _06078_ _06088_ _06089_ net39 vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__o221a_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18440_ _02466_ net4513 _02411_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _08310_ _08707_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__nor2_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ net29 net30 net31 vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a21oi_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14603_ _07367_ _07523_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__or2_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _04950_ _04951_ _04947_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__o21ai_2
X_18371_ net4538 net4405 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__and2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _08596_ _08597_ _08613_ _08644_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__nand4_1
XFILLER_0_29_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ net27 _05953_ net23 net24 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__and4b_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _10090_ _10322_ vssd1 vssd1 vccd1 vccd1 _10323_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ net1060 net1915 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nand2_1
X_14534_ _07643_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17253_ _10136_ _10146_ _10144_ vssd1 vssd1 vccd1 vccd1 _10254_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0__03991_ _03991_ vssd1 vssd1 vccd1 vccd1 clknet_0__03991_ sky130_fd_sc_hd__clkbuf_16
X_14465_ _07551_ _07552_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__xnor2_1
X_11677_ net3028 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16204_ _09276_ net2943 vssd1 vssd1 vccd1 vccd1 _09279_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10628_ net7161 net7272 _04170_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__mux2_1
X_13416_ _06561_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__xor2_1
X_17184_ _10184_ _10185_ vssd1 vssd1 vccd1 vccd1 _10186_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14396_ _07515_ _07516_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16135_ _08449_ _08588_ _08565_ _09064_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13347_ net645 _06430_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16066_ _09138_ _08517_ _08874_ _09139_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__o22ai_1
X_13278_ _06414_ _06415_ _06419_ _06424_ _06428_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12229_ rbzero.debug_overlay.vplaneY\[-3\] _05373_ _05395_ _05397_ vssd1 vssd1 vccd1
+ vccd1 _05398_ sky130_fd_sc_hd__a211o_1
X_15017_ _08150_ _08095_ _08154_ _08068_ net6162 vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__a221o_4
Xhold2509 net4339 vssd1 vssd1 vccd1 vccd1 net3033 sky130_fd_sc_hd__dlygate4sd3_1
X_19825_ net3927 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1808 net6839 vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1819 net7055 vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19756_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__buf_2
X_16968_ net2787 _09968_ _09980_ vssd1 vssd1 vccd1 vccd1 _09982_ sky130_fd_sc_hd__o21a_1
XFILLER_0_194_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18707_ _02696_ _02700_ _02710_ _04623_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15919_ _08947_ _08993_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__06044_ clknet_0__06044_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__06044_
+ sky130_fd_sc_hd__clkbuf_16
X_19687_ net1768 _03375_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__or2_1
X_16899_ net1011 _09937_ _09938_ rbzero.wall_tracer.visualWallDist\[-9\] vssd1 vssd1
+ vccd1 vccd1 _00501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18638_ _02646_ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ _02574_ _02580_ net7585 net4691 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20600_ net56 _03026_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__and2_1
X_21580_ clknet_leaf_2_i_clk net5277 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20531_ _03880_ net3801 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20884__300 clknet_1_1__leaf__04002_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__inv_2
XFILLER_0_144_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20462_ net3784 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22201_ net333 net2426 vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5102 net1341 vssd1 vssd1 vccd1 vccd1 net5626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5113 _01088_ vssd1 vssd1 vccd1 vccd1 net5637 sky130_fd_sc_hd__dlygate4sd3_1
X_20393_ net3317 net1245 _03801_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__mux2_1
Xhold5124 rbzero.spi_registers.texadd0\[9\] vssd1 vssd1 vccd1 vccd1 net5648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5135 rbzero.spi_registers.texadd1\[21\] vssd1 vssd1 vccd1 vccd1 net5659 sky130_fd_sc_hd__dlygate4sd3_1
X_22132_ net264 net2229 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4401 rbzero.wall_tracer.trackDistX\[-4\] vssd1 vssd1 vccd1 vccd1 net4925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5146 _00708_ vssd1 vssd1 vccd1 vccd1 net5670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4412 net1144 vssd1 vssd1 vccd1 vccd1 net4936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5157 net1379 vssd1 vssd1 vccd1 vccd1 net5681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4423 _04636_ vssd1 vssd1 vccd1 vccd1 net4947 sky130_fd_sc_hd__buf_4
Xhold5168 net1416 vssd1 vssd1 vccd1 vccd1 net5692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4434 gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 net4958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5179 _00686_ vssd1 vssd1 vccd1 vccd1 net5703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3700 _03382_ vssd1 vssd1 vccd1 vccd1 net4224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4445 _01035_ vssd1 vssd1 vccd1 vccd1 net4969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22063_ clknet_leaf_7_i_clk net3571 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3711 net4242 vssd1 vssd1 vccd1 vccd1 net4235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4456 _00799_ vssd1 vssd1 vccd1 vccd1 net4980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4467 net736 vssd1 vssd1 vccd1 vccd1 net4991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3722 net1960 vssd1 vssd1 vccd1 vccd1 net4246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4478 rbzero.spi_registers.texadd3\[17\] vssd1 vssd1 vccd1 vccd1 net5002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3733 net7669 vssd1 vssd1 vccd1 vccd1 net4257 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0__f__03980_ clknet_0__03980_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03980_
+ sky130_fd_sc_hd__clkbuf_16
Xhold3744 net2280 vssd1 vssd1 vccd1 vccd1 net4268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4489 rbzero.spi_registers.buf_mapdy\[3\] vssd1 vssd1 vccd1 vccd1 net5013 sky130_fd_sc_hd__dlygate4sd3_1
X_21014_ net839 net4975 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__or2_1
Xhold3755 _00485_ vssd1 vssd1 vccd1 vccd1 net4279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3766 net1020 vssd1 vssd1 vccd1 vccd1 net4290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3777 _00960_ vssd1 vssd1 vccd1 vccd1 net4301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3788 net7739 vssd1 vssd1 vccd1 vccd1 net4312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3799 _00945_ vssd1 vssd1 vccd1 vccd1 net4323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21916_ clknet_leaf_92_i_clk net1494 vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21847_ clknet_leaf_82_i_clk net1227 vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11600_ rbzero.spi_registers.texadd3\[1\] _04640_ _04642_ rbzero.spi_registers.texadd2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _05476_ vssd1 vssd1 vccd1 vccd1 _05745_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21778_ clknet_leaf_20_i_clk net2284 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd3\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ rbzero.spi_registers.texadd2\[22\] _04693_ _04644_ rbzero.spi_registers.texadd1\[22\]
+ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250_ _06859_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__or2_1
X_11462_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__buf_4
XFILLER_0_191_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13201_ _06353_ _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nor2_1
Xhold7071 net4398 vssd1 vssd1 vccd1 vccd1 net7595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _07326_ _07327_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7082 rbzero.wall_tracer.stepDistX\[-4\] vssd1 vssd1 vccd1 vccd1 net7606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11393_ net7137 net2809 _04573_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold7093 rbzero.spi_registers.texadd1\[16\] vssd1 vssd1 vccd1 vccd1 net7617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6370 net2524 vssd1 vssd1 vccd1 vccd1 net6894 sky130_fd_sc_hd__dlygate4sd3_1
X_13132_ _06287_ net3426 vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__nor2_1
Xhold6381 rbzero.tex_r1\[48\] vssd1 vssd1 vccd1 vccd1 net6905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6392 net2110 vssd1 vssd1 vccd1 vccd1 net6916 sky130_fd_sc_hd__dlygate4sd3_1
X_17940_ _08546_ _09538_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ net6251 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__inv_2
Xhold5680 _08212_ vssd1 vssd1 vccd1 vccd1 net6204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold5691 net749 vssd1 vssd1 vccd1 vccd1 net6215 sky130_fd_sc_hd__dlygate4sd3_1
X_12014_ net1524 _04999_ _05022_ net1326 _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__o221a_1
X_17871_ _01684_ _10520_ _10407_ _10416_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__or4_1
Xhold4990 _00682_ vssd1 vssd1 vccd1 vccd1 net5514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19610_ net5030 net799 _03341_ _03330_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__o211a_1
X_16822_ _09887_ _09888_ _09890_ vssd1 vssd1 vccd1 vccd1 _09892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19541_ _08279_ net3865 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__and2_1
X_16753_ _09820_ _09821_ vssd1 vssd1 vccd1 vccd1 _09823_ sky130_fd_sc_hd__and2_1
X_13965_ _06862_ net564 vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15704_ _08772_ _08770_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__or2b_1
X_19472_ _02996_ net3077 net1616 _03233_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__o211a_1
X_12916_ net35 _06046_ net4043 _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a31o_1
X_16684_ _09751_ _09753_ vssd1 vssd1 vccd1 vccd1 _09755_ sky130_fd_sc_hd__nand2_1
X_13896_ _06837_ _06922_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__nor2_1
X_18423_ _02451_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__clkbuf_1
X_15635_ _08704_ _08709_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ net32 _06001_ _06003_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18354_ net4453 net3505 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__nor2_1
X_15566_ _06211_ _08540_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12778_ _05904_ _05937_ _05896_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__a21o_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17305_ _10304_ _10305_ vssd1 vssd1 vccd1 vccd1 _10306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ _07649_ _07667_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_154_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11729_ net4345 net2825 net2895 net2774 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__or4_1
X_18285_ _02270_ _02327_ _02328_ _02330_ _09999_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a311o_1
X_15497_ _08570_ _08571_ vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17236_ _09251_ _09562_ _08849_ _09306_ vssd1 vssd1 vccd1 vccd1 _10237_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _07444_ _07598_ _07439_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _08632_ _08664_ vssd1 vssd1 vccd1 vccd1 _10169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold905 _01418_ vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ _07471_ _07400_ _07439_ _07367_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__o22a_1
Xhold916 net5695 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold927 net4102 vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ _08394_ _08484_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__or2_1
Xhold938 _04532_ vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17098_ _10098_ _10099_ vssd1 vssd1 vccd1 vccd1 _10100_ sky130_fd_sc_hd__xnor2_1
Xhold949 _04250_ vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3007 _03870_ vssd1 vssd1 vccd1 vccd1 net3531 sky130_fd_sc_hd__dlygate4sd3_1
X_16049_ _09102_ _09110_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__or2_1
Xhold3018 net4590 vssd1 vssd1 vccd1 vccd1 net3542 sky130_fd_sc_hd__buf_1
Xhold3029 net4769 vssd1 vssd1 vccd1 vccd1 net3553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2306 net7287 vssd1 vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2317 net3944 vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2328 _04286_ vssd1 vssd1 vccd1 vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2339 _01451_ vssd1 vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 _04430_ vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1616 net6883 vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_19808_ net4401 _03426_ net2231 _03454_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__o211a_1
Xhold1627 _01320_ vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1638 _01165_ vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 net1756 vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19739_ net6058 _03407_ net1785 _03413_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20916__329 clknet_1_1__leaf__04005_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__inv_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21701_ clknet_leaf_101_i_clk net4993 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.buf_texadd0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21632_ clknet_leaf_19_i_clk net5093 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21563_ clknet_leaf_17_i_clk net5269 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20514_ net3611 net1324 _03867_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21494_ clknet_leaf_15_i_clk net2537 vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20445_ _03836_ net3844 vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20376_ net3615 net3737 _03782_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
Xhold4220 net2909 vssd1 vssd1 vccd1 vccd1 net4744 sky130_fd_sc_hd__dlygate4sd3_1
X_22115_ net247 net1882 vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold4231 _00585_ vssd1 vssd1 vccd1 vccd1 net4755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4253 _01008_ vssd1 vssd1 vccd1 vccd1 net4777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_140_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4264 _00591_ vssd1 vssd1 vccd1 vccd1 net4788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4275 rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 net4799 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3530 _09924_ vssd1 vssd1 vccd1 vccd1 net4054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4286 _02689_ vssd1 vssd1 vccd1 vccd1 net4810 sky130_fd_sc_hd__dlygate4sd3_1
X_22046_ clknet_leaf_91_i_clk net3340 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold3541 _04859_ vssd1 vssd1 vccd1 vccd1 net4065 sky130_fd_sc_hd__buf_1
Xhold3552 net5995 vssd1 vssd1 vccd1 vccd1 net4076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4297 net6112 vssd1 vssd1 vccd1 vccd1 net4821 sky130_fd_sc_hd__buf_2
Xhold3563 _04646_ vssd1 vssd1 vccd1 vccd1 net4087 sky130_fd_sc_hd__clkbuf_2
Xhold3574 gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 net4098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3585 net694 vssd1 vssd1 vccd1 vccd1 net4109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2840 rbzero.pov.ready_buffer\[44\] vssd1 vssd1 vccd1 vccd1 net3364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2851 _02983_ vssd1 vssd1 vccd1 vccd1 net3375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3596 net599 vssd1 vssd1 vccd1 vccd1 net4120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2862 _01245_ vssd1 vssd1 vccd1 vccd1 net3386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2873 net3418 vssd1 vssd1 vccd1 vccd1 net3397 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2895 net3397 vssd1 vssd1 vccd1 vccd1 net3419 sky130_fd_sc_hd__buf_1
X_10962_ net2491 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
X_13750_ _06894_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20856__276 clknet_1_0__leaf__03998_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__inv_2
XFILLER_0_211_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12701_ net44 _05854_ _05843_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ net2626 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13681_ _06659_ _06791_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__or3b_2
XFILLER_0_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ _06178_ _08314_ _08473_ _08494_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ net9 _05793_ net5 net6 vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__and4b_1
XFILLER_0_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _05726_ _05727_ _05019_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__mux2_1
X_15351_ _08423_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14302_ _07448_ _07452_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__xor2_1
X_11514_ rbzero.spi_registers.texadd3\[14\] _04640_ _04642_ rbzero.spi_registers.texadd2\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a22oi_2
X_18070_ _10379_ _09536_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12494_ _05229_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15282_ net2940 vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17021_ net7796 _10028_ _10029_ vssd1 vssd1 vccd1 vccd1 _10030_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14233_ _07374_ _07383_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__xor2_1
X_11445_ net4103 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__inv_2
XFILLER_0_180_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _06931_ _06973_ _07268_ _06866_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__and4bb_1
X_11376_ net2712 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13115_ net3494 vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__inv_2
X_14095_ _07159_ _06970_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__nand2_1
X_18972_ net3999 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__clkbuf_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _06180_ net4823 vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__nand2_1
X_17923_ _01972_ net4558 _01749_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17854_ _01902_ _01903_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16805_ _09871_ _09872_ _09874_ vssd1 vssd1 vccd1 vccd1 _09875_ sky130_fd_sc_hd__nand3_1
X_17785_ _01835_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__buf_2
X_14997_ _08026_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__buf_4
XFILLER_0_205_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19524_ _02492_ _02497_ _02498_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__nand3_2
X_16736_ _08310_ _09805_ vssd1 vssd1 vccd1 vccd1 _09806_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13948_ _07086_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19455_ _03088_ net3181 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or2_1
X_16667_ _08633_ _09736_ _09737_ _08610_ vssd1 vssd1 vccd1 vccd1 _09738_ sky130_fd_sc_hd__a31o_4
X_13879_ _07026_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18406_ _02436_ net4613 _02411_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
X_15618_ _08691_ _08692_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19386_ net2354 _03199_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__or2_1
X_16598_ _09541_ _09668_ vssd1 vssd1 vccd1 vccd1 _09669_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18337_ net4491 net4473 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15549_ _08622_ _08612_ net7444 _08596_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__or4b_4
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18268_ _02312_ _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17219_ _10106_ _10120_ _10118_ vssd1 vssd1 vccd1 vccd1 _10220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18199_ _02244_ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__nand2_1
Xhold702 net3351 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 net3640 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
X_20230_ net5219 _03731_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold724 net5771 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 net6438 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 net5239 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold757 net5592 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 net5543 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
X_20161_ net1276 _03692_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold779 net4882 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2103 _01453_ vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 net7108 vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
X_20092_ net2628 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__inv_2
Xhold2125 _01585_ vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2136 _04395_ vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2147 net7259 vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1402 net7070 vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2158 net7246 vssd1 vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _01346_ vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1424 net6733 vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold2169 _04586_ vssd1 vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 net7663 vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 net5952 vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1457 _01398_ vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1468 net5810 vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1479 _01426_ vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21615_ clknet_leaf_25_i_clk net5538 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21546_ clknet_leaf_27_i_clk net1321 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.texadd0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21477_ clknet_leaf_102_i_clk net3110 vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11230_ net6504 net2197 _04492_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__mux2_1
X_20428_ net3352 net1280 _03823_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ net2140 net5814 _04459_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
Xhold4050 net7914 vssd1 vssd1 vccd1 vccd1 net4574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4061 net7899 vssd1 vssd1 vccd1 vccd1 net4585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold4072 net7560 vssd1 vssd1 vccd1 vccd1 net4596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11092_ net2049 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
Xhold4083 net767 vssd1 vssd1 vccd1 vccd1 net4607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4094 rbzero.wall_tracer.stepDistX\[8\] vssd1 vssd1 vccd1 vccd1 net4618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3360 _00594_ vssd1 vssd1 vccd1 vccd1 net3884 sky130_fd_sc_hd__dlygate4sd3_1
X_22029_ clknet_leaf_96_i_clk net3299 vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14920_ net7436 vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__clkbuf_4
Xhold3371 _02742_ vssd1 vssd1 vccd1 vccd1 net3895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold3382 _02978_ vssd1 vssd1 vccd1 vccd1 net3906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3393 net6206 vssd1 vssd1 vccd1 vccd1 net3917 sky130_fd_sc_hd__clkbuf_4
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2670 rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 net3194 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2681 _00579_ vssd1 vssd1 vccd1 vccd1 net3205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 net2013 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net7434 _07986_ _07988_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__and3_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2692 net4718 vssd1 vssd1 vccd1 vccd1 net3216 sky130_fd_sc_hd__clkbuf_2
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 net4128 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 _03158_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _06929_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__inv_2
Xhold1980 _01157_ vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_17570_ _10462_ _10464_ _10568_ vssd1 vssd1 vccd1 vccd1 _10569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1991 net6959 vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_14782_ _07922_ _07932_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__or2_1
X_11994_ net3016 _04713_ _04719_ net1603 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a211oi_1
X_16521_ _08587_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__clkbuf_4
X_13733_ net578 _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__nand2_1
X_10945_ net6553 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19240_ net5128 _03119_ _03122_ _03115_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16452_ _09405_ _09408_ _09523_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__nor3_1
X_13664_ _06657_ _06814_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10876_ net6922 net5911 _04310_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ net7939 _08298_ _08327_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__a21oi_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ net5656 _03078_ _03080_ _03074_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12615_ reg_rgb\[23\] _05779_ _05204_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__mux2_2
X_16383_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__xnor2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _06744_ _06745_ _06692_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__a21oi_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18122_ _02166_ _02169_ net3508 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a21oi_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _08298_ _08407_ _08408_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__a21oi_4
X_12546_ rbzero.tex_b1\[59\] rbzero.tex_b1\[58\] _05541_ vssd1 vssd1 vccd1 vccd1 _05711_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18053_ _02099_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15265_ _06470_ _06489_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__nor2_1
X_12477_ _05248_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__or2_1
X_17004_ _10005_ _10006_ _10007_ vssd1 vssd1 vccd1 vccd1 _10014_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ net544 vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__buf_2
X_11428_ net3760 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__clkbuf_4
X_15196_ _08276_ net4045 vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ net6479 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
X_14147_ _07071_ _07255_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14078_ _07163_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__xnor2_1
X_18955_ net4634 _05391_ _02928_ _02864_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _01953_ _01954_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__nand2_1
X_13029_ net4896 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__buf_2
X_18886_ _02844_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__and3_1
X_17837_ _01885_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer16 net3132 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_6
Xrebuffer27 _07137_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_1
X_17768_ _01808_ _01818_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__xnor2_1
Xrebuffer38 _06819_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_6
X_20839__260 clknet_1_1__leaf__03997_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__inv_2
Xrebuffer49 _06858_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_1
XFILLER_0_117_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16719_ _09669_ _09786_ vssd1 vssd1 vccd1 vccd1 _09789_ sky130_fd_sc_hd__nand2_1
X_19507_ net3096 _03275_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17699_ _01750_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__clkbuf_1
X_19438_ net5106 _03224_ _03234_ _03233_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ net4291 _03185_ net595 _03194_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21400_ clknet_leaf_64_i_clk _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22380_ net512 net2780 vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold6903 rbzero.debug_overlay.playerX\[-4\] vssd1 vssd1 vccd1 vccd1 net7427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ clknet_leaf_57_i_clk net4234 vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6914 _07311_ vssd1 vssd1 vccd1 vccd1 net7438 sky130_fd_sc_hd__buf_2
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6925 net4184 vssd1 vssd1 vccd1 vccd1 net7449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6936 rbzero.wall_tracer.trackDistX\[-11\] vssd1 vssd1 vccd1 vccd1 net7460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold6947 rbzero.traced_texVinit\[7\] vssd1 vssd1 vccd1 vccd1 net7471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6958 rbzero.traced_texVinit\[0\] vssd1 vssd1 vccd1 vccd1 net7482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6969 rbzero.wall_tracer.stepDistX\[1\] vssd1 vssd1 vccd1 vccd1 net7493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold510 net3309 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
X_21262_ clknet_leaf_71_i_clk net3774 vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold521 net5390 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold532 net5397 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20213_ net3530 _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__or2_1
Xhold543 net5396 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 net5476 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 net6376 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21193_ net4438 net723 vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold576 net7569 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold587 net6384 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 _01452_ vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
X_20144_ net5209 _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__or2_1
X_20981__8 clknet_1_0__leaf__04011_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ net4459 _03581_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__or2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _01503_ vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _03439_ vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 net2172 vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1243 _01371_ vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1254 net6633 vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1265 _00903_ vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1276 net6695 vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 _01299_ vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _04359_ vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ net6900 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10661_ net5823 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _04979_ _05554_ _05558_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__o31a_1
X_13380_ _06519_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__or2b_4
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12331_ _05495_ _05498_ net80 vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21529_ clknet_leaf_34_i_clk net5153 vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20667__105 clknet_1_1__leaf__03980_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__inv_2
XFILLER_0_181_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ _08182_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ _05390_ _05411_ _05419_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a31o_1
XFILLER_0_161_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ net6790 net6912 _04481_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14001_ _07085_ net75 vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12193_ _05343_ _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__nand2_1
X_11144_ net6756 net6570 _04448_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__mux2_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__buf_1
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18740_ _06183_ _06396_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__xnor2_1
X_15952_ _09015_ _09016_ _09026_ vssd1 vssd1 vccd1 vccd1 _09027_ sky130_fd_sc_hd__a21o_1
X_11075_ net6610 net2237 _04415_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__mux2_1
Xhold3190 _03885_ vssd1 vssd1 vccd1 vccd1 net3714 sky130_fd_sc_hd__dlygate4sd3_1
X_14903_ net7566 _08051_ vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__nand2_1
X_18671_ _02646_ net3242 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__or2_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08410_ _08625_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _10537_ _10530_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__or2b_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14834_ _07578_ _07581_ _07983_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__04010_ _04010_ vssd1 vssd1 vccd1 vccd1 clknet_0__04010_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17553_ _10550_ _10551_ vssd1 vssd1 vccd1 vccd1 _10552_ sky130_fd_sc_hd__nor2_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _07913_ _07915_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11977_ net1673 _04726_ _04776_ _05140_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _09574_ _09575_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__nor2_1
X_13716_ _06866_ _06857_ _06668_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__a21o_2
X_10928_ net2210 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
X_17484_ _10481_ _10482_ vssd1 vssd1 vccd1 vccd1 _10483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14696_ _07846_ _07844_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ net5802 _03106_ _03112_ _03096_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__o211a_1
X_16435_ _09506_ _09507_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ _06662_ _06746_ _06749_ _06762_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__o31a_1
X_10859_ net6992 net6531 _04299_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ net5497 _03065_ _03070_ _03061_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__o211a_1
X_16366_ _09345_ _09417_ _09437_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__nand3_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13578_ _06720_ _06726_ _06728_ _06725_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o22a_1
X_18105_ _02019_ _02057_ _02055_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15317_ net3315 _08305_ _08311_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19085_ _03027_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
X_12529_ _05189_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__nand2_1
X_16297_ net3539 _08313_ _08628_ _09368_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__or4_2
XFILLER_0_140_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5509 net1613 vssd1 vssd1 vccd1 vccd1 net6033 sky130_fd_sc_hd__buf_1
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _02023_ _02083_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15248_ _06625_ _08024_ _08320_ net7590 vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4808 net916 vssd1 vssd1 vccd1 vccd1 net5332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4819 _00734_ vssd1 vssd1 vccd1 vccd1 net5343 sky130_fd_sc_hd__dlygate4sd3_1
X_15179_ _08268_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19987_ rbzero.debug_overlay.facingX\[-3\] net3139 _03581_ vssd1 vssd1 vccd1 vccd1
+ _03591_ sky130_fd_sc_hd__mux2_1
X_20995__21 clknet_1_1__leaf__04012_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
X_18938_ _02919_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__nand2_1
.ends

