VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 587.945 BY 598.665 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 594.665 575.830 598.665 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 355.680 587.945 356.280 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 255.720 587.945 256.320 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 84.360 587.945 84.960 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 98.640 587.945 99.240 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 112.920 587.945 113.520 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 127.200 587.945 127.800 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 141.480 587.945 142.080 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 155.760 587.945 156.360 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 170.040 587.945 170.640 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 184.320 587.945 184.920 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 198.600 587.945 199.200 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 212.880 587.945 213.480 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 227.160 587.945 227.760 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 241.440 587.945 242.040 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 270.000 587.945 270.600 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 284.280 587.945 284.880 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 298.560 587.945 299.160 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 312.840 587.945 313.440 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 327.120 587.945 327.720 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 341.400 587.945 342.000 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 369.960 587.945 370.560 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 384.240 587.945 384.840 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 398.520 587.945 399.120 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 412.800 587.945 413.400 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 427.080 587.945 427.680 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 441.360 587.945 441.960 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 455.640 587.945 456.240 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 469.920 587.945 470.520 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 484.200 587.945 484.800 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 498.480 587.945 499.080 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 512.760 587.945 513.360 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 527.040 587.945 527.640 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 541.320 587.945 541.920 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 555.600 587.945 556.200 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 569.880 587.945 570.480 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 27.240 587.945 27.840 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 41.520 587.945 42.120 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 55.800 587.945 56.400 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 70.080 587.945 70.680 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 584.160 587.945 584.760 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 594.665 12.330 598.665 ;
    END
  END i_spare_1
  PIN i_test_uc2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 583.945 12.960 587.945 13.560 ;
    END
  END i_test_uc2
  PIN i_test_wci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END i_test_wci
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 594.665 58.330 598.665 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 594.665 46.830 598.665 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 594.665 35.330 598.665 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 594.665 23.830 598.665 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 594.665 127.330 598.665 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 594.665 115.830 598.665 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 594.665 104.330 598.665 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 594.665 92.830 598.665 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 594.665 81.330 598.665 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 594.665 69.830 598.665 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 594.665 196.330 598.665 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 594.665 173.330 598.665 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 594.665 161.830 598.665 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 594.665 150.330 598.665 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 594.665 138.830 598.665 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 594.665 184.830 598.665 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 594.665 564.330 598.665 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 594.665 449.330 598.665 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 594.665 437.830 598.665 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 594.665 426.330 598.665 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 594.665 414.830 598.665 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 594.665 403.330 598.665 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 594.665 391.830 598.665 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 594.665 552.830 598.665 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 594.665 541.330 598.665 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 594.665 529.830 598.665 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 594.665 518.330 598.665 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 594.665 506.830 598.665 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 594.665 495.330 598.665 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 594.665 483.830 598.665 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 594.665 472.330 598.665 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 594.665 460.830 598.665 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 594.665 380.330 598.665 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 594.665 265.330 598.665 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 594.665 253.830 598.665 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 594.665 242.330 598.665 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 594.665 230.830 598.665 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 594.665 219.330 598.665 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 594.665 207.830 598.665 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 594.665 368.830 598.665 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 594.665 357.330 598.665 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 594.665 345.830 598.665 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 594.665 334.330 598.665 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 594.665 322.830 598.665 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 594.665 311.330 598.665 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 594.665 299.830 598.665 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 594.665 288.330 598.665 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 594.665 276.830 598.665 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 582.550 586.215 ;
        RECT 5.330 577.945 582.550 580.775 ;
        RECT 5.330 572.505 582.550 575.335 ;
        RECT 5.330 567.065 582.550 569.895 ;
        RECT 5.330 561.625 582.550 564.455 ;
        RECT 5.330 556.185 582.550 559.015 ;
        RECT 5.330 550.745 582.550 553.575 ;
        RECT 5.330 545.305 582.550 548.135 ;
        RECT 5.330 539.865 582.550 542.695 ;
        RECT 5.330 534.425 582.550 537.255 ;
        RECT 5.330 528.985 582.550 531.815 ;
        RECT 5.330 523.545 582.550 526.375 ;
        RECT 5.330 518.105 582.550 520.935 ;
        RECT 5.330 512.665 582.550 515.495 ;
        RECT 5.330 507.225 582.550 510.055 ;
        RECT 5.330 501.785 582.550 504.615 ;
        RECT 5.330 496.345 582.550 499.175 ;
        RECT 5.330 490.905 582.550 493.735 ;
        RECT 5.330 485.465 582.550 488.295 ;
        RECT 5.330 480.025 582.550 482.855 ;
        RECT 5.330 474.585 582.550 477.415 ;
        RECT 5.330 469.145 582.550 471.975 ;
        RECT 5.330 463.705 582.550 466.535 ;
        RECT 5.330 458.265 582.550 461.095 ;
        RECT 5.330 452.825 582.550 455.655 ;
        RECT 5.330 447.385 582.550 450.215 ;
        RECT 5.330 441.945 582.550 444.775 ;
        RECT 5.330 436.505 582.550 439.335 ;
        RECT 5.330 431.065 582.550 433.895 ;
        RECT 5.330 425.625 582.550 428.455 ;
        RECT 5.330 420.185 582.550 423.015 ;
        RECT 5.330 414.745 582.550 417.575 ;
        RECT 5.330 409.305 582.550 412.135 ;
        RECT 5.330 403.865 582.550 406.695 ;
        RECT 5.330 398.425 582.550 401.255 ;
        RECT 5.330 392.985 582.550 395.815 ;
        RECT 5.330 387.545 582.550 390.375 ;
        RECT 5.330 382.105 582.550 384.935 ;
        RECT 5.330 376.665 582.550 379.495 ;
        RECT 5.330 371.225 582.550 374.055 ;
        RECT 5.330 365.785 582.550 368.615 ;
        RECT 5.330 360.345 582.550 363.175 ;
        RECT 5.330 354.905 582.550 357.735 ;
        RECT 5.330 349.465 582.550 352.295 ;
        RECT 5.330 344.025 582.550 346.855 ;
        RECT 5.330 338.585 582.550 341.415 ;
        RECT 5.330 333.145 582.550 335.975 ;
        RECT 5.330 327.705 582.550 330.535 ;
        RECT 5.330 322.265 582.550 325.095 ;
        RECT 5.330 316.825 582.550 319.655 ;
        RECT 5.330 311.385 582.550 314.215 ;
        RECT 5.330 305.945 582.550 308.775 ;
        RECT 5.330 300.505 582.550 303.335 ;
        RECT 5.330 295.065 582.550 297.895 ;
        RECT 5.330 289.625 582.550 292.455 ;
        RECT 5.330 284.185 582.550 287.015 ;
        RECT 5.330 278.745 582.550 281.575 ;
        RECT 5.330 273.305 582.550 276.135 ;
        RECT 5.330 267.865 582.550 270.695 ;
        RECT 5.330 262.425 582.550 265.255 ;
        RECT 5.330 256.985 582.550 259.815 ;
        RECT 5.330 251.545 582.550 254.375 ;
        RECT 5.330 246.105 582.550 248.935 ;
        RECT 5.330 240.665 582.550 243.495 ;
        RECT 5.330 235.225 582.550 238.055 ;
        RECT 5.330 229.785 582.550 232.615 ;
        RECT 5.330 224.345 582.550 227.175 ;
        RECT 5.330 218.905 582.550 221.735 ;
        RECT 5.330 213.465 582.550 216.295 ;
        RECT 5.330 208.025 582.550 210.855 ;
        RECT 5.330 202.585 582.550 205.415 ;
        RECT 5.330 197.145 582.550 199.975 ;
        RECT 5.330 191.705 582.550 194.535 ;
        RECT 5.330 186.265 582.550 189.095 ;
        RECT 5.330 180.825 582.550 183.655 ;
        RECT 5.330 175.385 582.550 178.215 ;
        RECT 5.330 169.945 582.550 172.775 ;
        RECT 5.330 164.505 582.550 167.335 ;
        RECT 5.330 159.065 582.550 161.895 ;
        RECT 5.330 153.625 582.550 156.455 ;
        RECT 5.330 148.185 582.550 151.015 ;
        RECT 5.330 142.745 582.550 145.575 ;
        RECT 5.330 137.305 582.550 140.135 ;
        RECT 5.330 131.865 582.550 134.695 ;
        RECT 5.330 126.425 582.550 129.255 ;
        RECT 5.330 120.985 582.550 123.815 ;
        RECT 5.330 115.545 582.550 118.375 ;
        RECT 5.330 110.105 582.550 112.935 ;
        RECT 5.330 104.665 582.550 107.495 ;
        RECT 5.330 99.225 582.550 102.055 ;
        RECT 5.330 93.785 582.550 96.615 ;
        RECT 5.330 88.345 582.550 91.175 ;
        RECT 5.330 82.905 582.550 85.735 ;
        RECT 5.330 77.465 582.550 80.295 ;
        RECT 5.330 72.025 582.550 74.855 ;
        RECT 5.330 66.585 582.550 69.415 ;
        RECT 5.330 61.145 582.550 63.975 ;
        RECT 5.330 55.705 582.550 58.535 ;
        RECT 5.330 50.265 582.550 53.095 ;
        RECT 5.330 44.825 582.550 47.655 ;
        RECT 5.330 39.385 582.550 42.215 ;
        RECT 5.330 33.945 582.550 36.775 ;
        RECT 5.330 28.505 582.550 31.335 ;
        RECT 5.330 23.065 582.550 25.895 ;
        RECT 5.330 17.625 582.550 20.455 ;
        RECT 5.330 12.185 582.550 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 582.360 587.605 ;
      LAYER met1 ;
        RECT 5.520 9.900 582.360 587.760 ;
      LAYER met2 ;
        RECT 7.920 594.385 11.770 595.410 ;
        RECT 12.610 594.385 23.270 595.410 ;
        RECT 24.110 594.385 34.770 595.410 ;
        RECT 35.610 594.385 46.270 595.410 ;
        RECT 47.110 594.385 57.770 595.410 ;
        RECT 58.610 594.385 69.270 595.410 ;
        RECT 70.110 594.385 80.770 595.410 ;
        RECT 81.610 594.385 92.270 595.410 ;
        RECT 93.110 594.385 103.770 595.410 ;
        RECT 104.610 594.385 115.270 595.410 ;
        RECT 116.110 594.385 126.770 595.410 ;
        RECT 127.610 594.385 138.270 595.410 ;
        RECT 139.110 594.385 149.770 595.410 ;
        RECT 150.610 594.385 161.270 595.410 ;
        RECT 162.110 594.385 172.770 595.410 ;
        RECT 173.610 594.385 184.270 595.410 ;
        RECT 185.110 594.385 195.770 595.410 ;
        RECT 196.610 594.385 207.270 595.410 ;
        RECT 208.110 594.385 218.770 595.410 ;
        RECT 219.610 594.385 230.270 595.410 ;
        RECT 231.110 594.385 241.770 595.410 ;
        RECT 242.610 594.385 253.270 595.410 ;
        RECT 254.110 594.385 264.770 595.410 ;
        RECT 265.610 594.385 276.270 595.410 ;
        RECT 277.110 594.385 287.770 595.410 ;
        RECT 288.610 594.385 299.270 595.410 ;
        RECT 300.110 594.385 310.770 595.410 ;
        RECT 311.610 594.385 322.270 595.410 ;
        RECT 323.110 594.385 333.770 595.410 ;
        RECT 334.610 594.385 345.270 595.410 ;
        RECT 346.110 594.385 356.770 595.410 ;
        RECT 357.610 594.385 368.270 595.410 ;
        RECT 369.110 594.385 379.770 595.410 ;
        RECT 380.610 594.385 391.270 595.410 ;
        RECT 392.110 594.385 402.770 595.410 ;
        RECT 403.610 594.385 414.270 595.410 ;
        RECT 415.110 594.385 425.770 595.410 ;
        RECT 426.610 594.385 437.270 595.410 ;
        RECT 438.110 594.385 448.770 595.410 ;
        RECT 449.610 594.385 460.270 595.410 ;
        RECT 461.110 594.385 471.770 595.410 ;
        RECT 472.610 594.385 483.270 595.410 ;
        RECT 484.110 594.385 494.770 595.410 ;
        RECT 495.610 594.385 506.270 595.410 ;
        RECT 507.110 594.385 517.770 595.410 ;
        RECT 518.610 594.385 529.270 595.410 ;
        RECT 530.110 594.385 540.770 595.410 ;
        RECT 541.610 594.385 552.270 595.410 ;
        RECT 553.110 594.385 563.770 595.410 ;
        RECT 564.610 594.385 575.270 595.410 ;
        RECT 576.110 594.385 579.960 595.410 ;
        RECT 7.920 4.280 579.960 594.385 ;
        RECT 7.920 4.000 13.610 4.280 ;
        RECT 14.450 4.000 28.330 4.280 ;
        RECT 29.170 4.000 43.050 4.280 ;
        RECT 43.890 4.000 57.770 4.280 ;
        RECT 58.610 4.000 72.490 4.280 ;
        RECT 73.330 4.000 87.210 4.280 ;
        RECT 88.050 4.000 101.930 4.280 ;
        RECT 102.770 4.000 116.650 4.280 ;
        RECT 117.490 4.000 131.370 4.280 ;
        RECT 132.210 4.000 146.090 4.280 ;
        RECT 146.930 4.000 160.810 4.280 ;
        RECT 161.650 4.000 175.530 4.280 ;
        RECT 176.370 4.000 190.250 4.280 ;
        RECT 191.090 4.000 204.970 4.280 ;
        RECT 205.810 4.000 219.690 4.280 ;
        RECT 220.530 4.000 234.410 4.280 ;
        RECT 235.250 4.000 249.130 4.280 ;
        RECT 249.970 4.000 263.850 4.280 ;
        RECT 264.690 4.000 278.570 4.280 ;
        RECT 279.410 4.000 293.290 4.280 ;
        RECT 294.130 4.000 308.010 4.280 ;
        RECT 308.850 4.000 322.730 4.280 ;
        RECT 323.570 4.000 337.450 4.280 ;
        RECT 338.290 4.000 352.170 4.280 ;
        RECT 353.010 4.000 366.890 4.280 ;
        RECT 367.730 4.000 381.610 4.280 ;
        RECT 382.450 4.000 396.330 4.280 ;
        RECT 397.170 4.000 411.050 4.280 ;
        RECT 411.890 4.000 425.770 4.280 ;
        RECT 426.610 4.000 440.490 4.280 ;
        RECT 441.330 4.000 455.210 4.280 ;
        RECT 456.050 4.000 469.930 4.280 ;
        RECT 470.770 4.000 484.650 4.280 ;
        RECT 485.490 4.000 499.370 4.280 ;
        RECT 500.210 4.000 514.090 4.280 ;
        RECT 514.930 4.000 528.810 4.280 ;
        RECT 529.650 4.000 543.530 4.280 ;
        RECT 544.370 4.000 558.250 4.280 ;
        RECT 559.090 4.000 572.970 4.280 ;
        RECT 573.810 4.000 579.960 4.280 ;
      LAYER met3 ;
        RECT 13.405 585.160 583.945 587.685 ;
        RECT 13.405 583.760 583.545 585.160 ;
        RECT 13.405 570.880 583.945 583.760 ;
        RECT 13.405 569.480 583.545 570.880 ;
        RECT 13.405 556.600 583.945 569.480 ;
        RECT 13.405 555.200 583.545 556.600 ;
        RECT 13.405 542.320 583.945 555.200 ;
        RECT 13.405 540.920 583.545 542.320 ;
        RECT 13.405 528.040 583.945 540.920 ;
        RECT 13.405 526.640 583.545 528.040 ;
        RECT 13.405 513.760 583.945 526.640 ;
        RECT 13.405 512.360 583.545 513.760 ;
        RECT 13.405 499.480 583.945 512.360 ;
        RECT 13.405 498.080 583.545 499.480 ;
        RECT 13.405 485.200 583.945 498.080 ;
        RECT 13.405 483.800 583.545 485.200 ;
        RECT 13.405 470.920 583.945 483.800 ;
        RECT 13.405 469.520 583.545 470.920 ;
        RECT 13.405 456.640 583.945 469.520 ;
        RECT 13.405 455.240 583.545 456.640 ;
        RECT 13.405 442.360 583.945 455.240 ;
        RECT 13.405 440.960 583.545 442.360 ;
        RECT 13.405 428.080 583.945 440.960 ;
        RECT 13.405 426.680 583.545 428.080 ;
        RECT 13.405 413.800 583.945 426.680 ;
        RECT 13.405 412.400 583.545 413.800 ;
        RECT 13.405 399.520 583.945 412.400 ;
        RECT 13.405 398.120 583.545 399.520 ;
        RECT 13.405 385.240 583.945 398.120 ;
        RECT 13.405 383.840 583.545 385.240 ;
        RECT 13.405 370.960 583.945 383.840 ;
        RECT 13.405 369.560 583.545 370.960 ;
        RECT 13.405 356.680 583.945 369.560 ;
        RECT 13.405 355.280 583.545 356.680 ;
        RECT 13.405 342.400 583.945 355.280 ;
        RECT 13.405 341.000 583.545 342.400 ;
        RECT 13.405 328.120 583.945 341.000 ;
        RECT 13.405 326.720 583.545 328.120 ;
        RECT 13.405 313.840 583.945 326.720 ;
        RECT 13.405 312.440 583.545 313.840 ;
        RECT 13.405 299.560 583.945 312.440 ;
        RECT 13.405 298.160 583.545 299.560 ;
        RECT 13.405 285.280 583.945 298.160 ;
        RECT 13.405 283.880 583.545 285.280 ;
        RECT 13.405 271.000 583.945 283.880 ;
        RECT 13.405 269.600 583.545 271.000 ;
        RECT 13.405 256.720 583.945 269.600 ;
        RECT 13.405 255.320 583.545 256.720 ;
        RECT 13.405 242.440 583.945 255.320 ;
        RECT 13.405 241.040 583.545 242.440 ;
        RECT 13.405 228.160 583.945 241.040 ;
        RECT 13.405 226.760 583.545 228.160 ;
        RECT 13.405 213.880 583.945 226.760 ;
        RECT 13.405 212.480 583.545 213.880 ;
        RECT 13.405 199.600 583.945 212.480 ;
        RECT 13.405 198.200 583.545 199.600 ;
        RECT 13.405 185.320 583.945 198.200 ;
        RECT 13.405 183.920 583.545 185.320 ;
        RECT 13.405 171.040 583.945 183.920 ;
        RECT 13.405 169.640 583.545 171.040 ;
        RECT 13.405 156.760 583.945 169.640 ;
        RECT 13.405 155.360 583.545 156.760 ;
        RECT 13.405 142.480 583.945 155.360 ;
        RECT 13.405 141.080 583.545 142.480 ;
        RECT 13.405 128.200 583.945 141.080 ;
        RECT 13.405 126.800 583.545 128.200 ;
        RECT 13.405 113.920 583.945 126.800 ;
        RECT 13.405 112.520 583.545 113.920 ;
        RECT 13.405 99.640 583.945 112.520 ;
        RECT 13.405 98.240 583.545 99.640 ;
        RECT 13.405 85.360 583.945 98.240 ;
        RECT 13.405 83.960 583.545 85.360 ;
        RECT 13.405 71.080 583.945 83.960 ;
        RECT 13.405 69.680 583.545 71.080 ;
        RECT 13.405 56.800 583.945 69.680 ;
        RECT 13.405 55.400 583.545 56.800 ;
        RECT 13.405 42.520 583.945 55.400 ;
        RECT 13.405 41.120 583.545 42.520 ;
        RECT 13.405 28.240 583.945 41.120 ;
        RECT 13.405 26.840 583.545 28.240 ;
        RECT 13.405 13.960 583.945 26.840 ;
        RECT 13.405 12.560 583.545 13.960 ;
        RECT 13.405 10.715 583.945 12.560 ;
      LAYER met4 ;
        RECT 49.975 11.735 97.440 585.305 ;
        RECT 99.840 11.735 174.240 585.305 ;
        RECT 176.640 11.735 251.040 585.305 ;
        RECT 253.440 11.735 327.840 585.305 ;
        RECT 330.240 11.735 404.640 585.305 ;
        RECT 407.040 11.735 481.440 585.305 ;
        RECT 483.840 11.735 558.240 585.305 ;
        RECT 560.640 11.735 570.105 585.305 ;
  END
END top_ew_algofoogle
END LIBRARY

